//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n773_, new_n774_, new_n775_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n785_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n902_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n927_, new_n928_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n941_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n951_, new_n953_, new_n954_, new_n955_, new_n956_, new_n958_,
    new_n959_, new_n960_;
  INV_X1    g000(.A(G183gat), .ZN(new_n202_));
  INV_X1    g001(.A(G190gat), .ZN(new_n203_));
  NOR3_X1   g002(.A1(new_n202_), .A2(new_n203_), .A3(KEYINPUT23), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT23), .B1(new_n202_), .B2(new_n203_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(KEYINPUT81), .B(G190gat), .Z(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(new_n202_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(G169gat), .ZN(new_n212_));
  AND2_X1   g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n206_), .A2(KEYINPUT84), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT84), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n215_), .B(KEYINPUT23), .C1(new_n202_), .C2(new_n203_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n204_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT26), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(G190gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT82), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n208_), .A2(KEYINPUT26), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT25), .B(G183gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n218_), .A2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(G169gat), .ZN(new_n228_));
  INV_X1    g027(.A(G176gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n227_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT83), .ZN(new_n231_));
  OR3_X1    g030(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT83), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n227_), .B(new_n233_), .C1(new_n228_), .C2(new_n229_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n231_), .A2(new_n232_), .A3(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n213_), .B1(new_n225_), .B2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G211gat), .B(G218gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT94), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G197gat), .B(G204gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT21), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n241_), .A2(new_n242_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n240_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT95), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n238_), .B(KEYINPUT94), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(new_n243_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n246_), .A2(new_n247_), .A3(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n247_), .B1(new_n246_), .B2(new_n249_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n237_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n246_), .A2(new_n249_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT26), .B(G190gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(new_n223_), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n207_), .A2(new_n232_), .A3(new_n230_), .A4(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(G183gat), .A2(G190gat), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n212_), .B1(new_n217_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT98), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT98), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n261_), .A2(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n259_), .B1(new_n263_), .B2(new_n265_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n253_), .B(KEYINPUT20), .C1(new_n255_), .C2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G226gat), .A2(G233gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT19), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT20), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n251_), .A2(new_n252_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n210_), .A2(new_n212_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n218_), .A2(new_n224_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n274_), .B1(new_n275_), .B2(new_n235_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n272_), .B1(new_n273_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n265_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n261_), .A2(new_n264_), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n255_), .B(new_n258_), .C1(new_n278_), .C2(new_n279_), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n267_), .A2(new_n269_), .B1(new_n277_), .B2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G8gat), .B(G36gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT18), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G64gat), .B(G92gat), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n283_), .B(new_n284_), .Z(new_n285_));
  NAND2_X1  g084(.A1(new_n281_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n285_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n269_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n252_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(new_n250_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n270_), .B1(new_n290_), .B2(new_n237_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n258_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(new_n254_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n288_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n289_), .A2(new_n276_), .A3(new_n250_), .ZN(new_n295_));
  AND3_X1   g094(.A1(new_n295_), .A2(new_n280_), .A3(new_n271_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n287_), .B1(new_n294_), .B2(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(KEYINPUT27), .B1(new_n286_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT27), .ZN(new_n299_));
  XOR2_X1   g098(.A(KEYINPUT100), .B(KEYINPUT20), .Z(new_n300_));
  NAND3_X1  g099(.A1(new_n246_), .A2(new_n249_), .A3(new_n258_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n300_), .B1(new_n301_), .B2(new_n262_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n302_), .B1(new_n273_), .B2(new_n276_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT101), .B1(new_n303_), .B2(new_n288_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n291_), .A2(new_n288_), .A3(new_n293_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT101), .ZN(new_n306_));
  INV_X1    g105(.A(new_n295_), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n306_), .B(new_n269_), .C1(new_n307_), .C2(new_n302_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n304_), .A2(new_n305_), .A3(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n299_), .B1(new_n309_), .B2(new_n287_), .ZN(new_n310_));
  AOI21_X1  g109(.A(KEYINPUT102), .B1(new_n281_), .B2(new_n285_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT102), .ZN(new_n312_));
  NOR4_X1   g111(.A1(new_n294_), .A2(new_n296_), .A3(new_n312_), .A4(new_n287_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n310_), .B1(new_n311_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT103), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT103), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n310_), .B(new_n316_), .C1(new_n311_), .C2(new_n313_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n298_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G78gat), .B(G106gat), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT96), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT1), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT87), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  OR2_X1    g124(.A1(new_n322_), .A2(KEYINPUT1), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT86), .ZN(new_n327_));
  INV_X1    g126(.A(G155gat), .ZN(new_n328_));
  INV_X1    g127(.A(G162gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT86), .B1(G155gat), .B2(G162gat), .ZN(new_n331_));
  AND3_X1   g130(.A1(new_n326_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n325_), .A2(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(G141gat), .A2(G148gat), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G141gat), .A2(G148gat), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n333_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n330_), .A2(new_n331_), .A3(new_n322_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT89), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n334_), .A2(KEYINPUT88), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n341_), .A2(KEYINPUT3), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(KEYINPUT3), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n336_), .B(KEYINPUT2), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n340_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT90), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT90), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n340_), .A2(new_n348_), .A3(new_n345_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n338_), .B1(new_n347_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT29), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n321_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n349_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n348_), .B1(new_n340_), .B2(new_n345_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n337_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n355_), .A2(KEYINPUT96), .A3(KEYINPUT29), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n352_), .A2(new_n254_), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(G233gat), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT93), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n359_), .A2(G228gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(G228gat), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n358_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n357_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT92), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n364_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n355_), .A2(KEYINPUT92), .A3(KEYINPUT29), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n290_), .A2(new_n362_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n320_), .B1(new_n363_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G22gat), .B(G50gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n350_), .A2(new_n351_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n373_), .A2(KEYINPUT28), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(KEYINPUT28), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n372_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n376_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n372_), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n378_), .A2(new_n374_), .A3(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n377_), .A2(new_n380_), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n357_), .A2(new_n362_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(new_n320_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n371_), .A2(new_n381_), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n371_), .A2(KEYINPUT97), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT97), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n370_), .A2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n386_), .A2(new_n388_), .A3(new_n383_), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT91), .B1(new_n377_), .B2(new_n380_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n379_), .B1(new_n378_), .B2(new_n374_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n375_), .A2(new_n376_), .A3(new_n372_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT91), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n391_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n390_), .A2(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n385_), .B1(new_n389_), .B2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G1gat), .B(G29gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(G85gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT0), .B(G57gat), .ZN(new_n399_));
  XOR2_X1   g198(.A(new_n398_), .B(new_n399_), .Z(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G127gat), .B(G134gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G113gat), .B(G120gat), .ZN(new_n403_));
  XOR2_X1   g202(.A(new_n402_), .B(new_n403_), .Z(new_n404_));
  NAND2_X1  g203(.A1(new_n355_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n404_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n350_), .A2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n405_), .A2(new_n407_), .A3(KEYINPUT4), .ZN(new_n408_));
  OR3_X1    g207(.A1(new_n350_), .A2(KEYINPUT4), .A3(new_n406_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G225gat), .A2(G233gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n408_), .A2(new_n409_), .A3(KEYINPUT99), .A4(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n405_), .A2(new_n407_), .A3(new_n410_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n411_), .B1(new_n405_), .B2(KEYINPUT4), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(KEYINPUT99), .B1(new_n416_), .B2(new_n408_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n401_), .B1(new_n414_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT99), .ZN(new_n419_));
  INV_X1    g218(.A(new_n408_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n419_), .B1(new_n420_), .B2(new_n415_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n421_), .A2(new_n413_), .A3(new_n400_), .A4(new_n412_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n418_), .A2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G71gat), .B(G99gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(G43gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n276_), .B(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G227gat), .A2(G233gat), .ZN(new_n427_));
  XOR2_X1   g226(.A(new_n427_), .B(G15gat), .Z(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(KEYINPUT30), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT31), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n426_), .A2(new_n430_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n426_), .A2(new_n430_), .ZN(new_n432_));
  OR3_X1    g231(.A1(new_n431_), .A2(new_n432_), .A3(KEYINPUT85), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT85), .B1(new_n431_), .B2(new_n432_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(new_n404_), .A3(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n434_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n406_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n423_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n318_), .A2(new_n396_), .A3(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n383_), .B1(new_n370_), .B2(new_n387_), .ZN(new_n440_));
  NOR3_X1   g239(.A1(new_n382_), .A2(KEYINPUT97), .A3(new_n320_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n395_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n423_), .B1(new_n442_), .B2(new_n384_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT33), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n422_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n414_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n446_), .A2(KEYINPUT33), .A3(new_n400_), .A4(new_n421_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n408_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n405_), .A2(new_n407_), .A3(new_n411_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n448_), .A2(new_n401_), .A3(new_n449_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n450_), .A2(new_n286_), .A3(new_n297_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n445_), .A2(new_n447_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n423_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n285_), .A2(KEYINPUT32), .ZN(new_n454_));
  MUX2_X1   g253(.A(new_n309_), .B(new_n281_), .S(new_n454_), .Z(new_n455_));
  OAI21_X1  g254(.A(new_n452_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n318_), .A2(new_n443_), .B1(new_n456_), .B2(new_n396_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n437_), .A2(new_n435_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n439_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT67), .ZN(new_n460_));
  XOR2_X1   g259(.A(G120gat), .B(G148gat), .Z(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT5), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G176gat), .B(G204gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(G64gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(G57gat), .ZN(new_n467_));
  INV_X1    g266(.A(G57gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(G64gat), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT66), .ZN(new_n470_));
  AND3_X1   g269(.A1(new_n467_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n470_), .B1(new_n467_), .B2(new_n469_), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT11), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n468_), .A2(G64gat), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n466_), .A2(G57gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT66), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT11), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n467_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G71gat), .B(G78gat), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n473_), .A2(new_n479_), .A3(new_n481_), .ZN(new_n482_));
  OAI211_X1 g281(.A(KEYINPUT11), .B(new_n480_), .C1(new_n471_), .C2(new_n472_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(G85gat), .ZN(new_n485_));
  INV_X1    g284(.A(G92gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G85gat), .A2(G92gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT64), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT7), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n491_), .B(new_n492_), .C1(G99gat), .C2(G106gat), .ZN(new_n493_));
  INV_X1    g292(.A(G99gat), .ZN(new_n494_));
  INV_X1    g293(.A(G106gat), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n494_), .B(new_n495_), .C1(KEYINPUT64), .C2(KEYINPUT7), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT65), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n493_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT6), .B1(new_n494_), .B2(new_n495_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT6), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(G99gat), .A3(G106gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n498_), .A2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n497_), .B1(new_n493_), .B2(new_n496_), .ZN(new_n504_));
  OAI211_X1 g303(.A(KEYINPUT8), .B(new_n490_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT8), .ZN(new_n506_));
  AOI22_X1  g305(.A1(new_n493_), .A2(new_n496_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n506_), .B1(new_n507_), .B2(new_n489_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n487_), .A2(KEYINPUT9), .A3(new_n488_), .ZN(new_n509_));
  OR2_X1    g308(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(new_n495_), .A3(new_n511_), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n488_), .A2(KEYINPUT9), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n502_), .A2(new_n509_), .A3(new_n512_), .A4(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n505_), .A2(new_n508_), .A3(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(KEYINPUT12), .B1(new_n484_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n482_), .A2(new_n483_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n493_), .A2(new_n496_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(new_n502_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(new_n490_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n502_), .A2(new_n513_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n512_), .A2(new_n509_), .ZN(new_n522_));
  AOI22_X1  g321(.A1(new_n520_), .A2(new_n506_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n517_), .A2(new_n523_), .A3(new_n505_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n490_), .A2(KEYINPUT8), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n498_), .A2(new_n502_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n504_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n525_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n489_), .B1(new_n518_), .B2(new_n502_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n514_), .B1(new_n529_), .B2(KEYINPUT8), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n483_), .B(new_n482_), .C1(new_n528_), .C2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n524_), .A2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n516_), .B1(new_n532_), .B2(KEYINPUT12), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G230gat), .A2(G233gat), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n534_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n532_), .A2(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n465_), .B1(new_n535_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT12), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n539_), .B1(new_n524_), .B2(new_n531_), .ZN(new_n540_));
  NOR3_X1   g339(.A1(new_n540_), .A2(new_n536_), .A3(new_n516_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n537_), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n541_), .A2(new_n542_), .A3(new_n464_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n460_), .B1(new_n538_), .B2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n535_), .A2(new_n537_), .A3(new_n465_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n464_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n545_), .A2(new_n546_), .A3(KEYINPUT67), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n544_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT13), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n544_), .A2(KEYINPUT13), .A3(new_n547_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G29gat), .B(G36gat), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT68), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n554_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G43gat), .B(G50gat), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n557_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G1gat), .B(G8gat), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT73), .ZN(new_n563_));
  INV_X1    g362(.A(G8gat), .ZN(new_n564_));
  INV_X1    g363(.A(G1gat), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(KEYINPUT72), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT72), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(G1gat), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n564_), .B1(new_n566_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT14), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n563_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(KEYINPUT72), .B(G1gat), .ZN(new_n572_));
  OAI211_X1 g371(.A(KEYINPUT73), .B(KEYINPUT14), .C1(new_n572_), .C2(new_n564_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  XOR2_X1   g373(.A(G15gat), .B(G22gat), .Z(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT74), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT74), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n574_), .A2(new_n579_), .A3(new_n576_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n562_), .B1(new_n578_), .B2(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n579_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n582_));
  AOI211_X1 g381(.A(KEYINPUT74), .B(new_n575_), .C1(new_n571_), .C2(new_n573_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n562_), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n582_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n561_), .B1(new_n581_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT78), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n578_), .A2(new_n580_), .A3(new_n562_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n584_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n561_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n588_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n586_), .A2(new_n587_), .A3(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n581_), .A2(new_n585_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n593_), .A2(KEYINPUT78), .A3(new_n590_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G229gat), .A2(G233gat), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT15), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n599_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n553_), .B(new_n554_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n557_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(KEYINPUT15), .A3(new_n558_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n600_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT79), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n588_), .A2(new_n605_), .A3(new_n589_), .A4(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n588_), .A2(new_n605_), .A3(new_n589_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT79), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n590_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n596_), .B(new_n607_), .C1(new_n609_), .C2(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(G113gat), .B(G141gat), .Z(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT80), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G169gat), .B(G197gat), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n613_), .B(new_n614_), .Z(new_n615_));
  NAND3_X1  g414(.A1(new_n598_), .A2(new_n611_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n615_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n611_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n596_), .B1(new_n592_), .B2(new_n594_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n617_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n552_), .B1(new_n616_), .B2(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n459_), .A2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G190gat), .B(G218gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G134gat), .B(G162gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT36), .Z(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n605_), .A2(new_n515_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n561_), .A2(new_n505_), .A3(new_n523_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G232gat), .A2(G233gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT34), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT35), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n628_), .A2(new_n629_), .A3(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n635_), .A2(KEYINPUT35), .A3(new_n631_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n631_), .A2(KEYINPUT35), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n628_), .A2(new_n637_), .A3(new_n629_), .A4(new_n634_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n627_), .B1(new_n636_), .B2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n625_), .A2(KEYINPUT36), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n636_), .A2(new_n640_), .A3(new_n638_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT69), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n636_), .A2(KEYINPUT69), .A3(new_n640_), .A4(new_n638_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n639_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT37), .ZN(new_n646_));
  OR3_X1    g445(.A1(new_n645_), .A2(KEYINPUT70), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT71), .ZN(new_n648_));
  INV_X1    g447(.A(new_n636_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n638_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n648_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n636_), .A2(KEYINPUT71), .A3(new_n638_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n651_), .A2(new_n652_), .A3(new_n626_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n643_), .A2(new_n644_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n653_), .A2(new_n654_), .A3(new_n646_), .ZN(new_n655_));
  OAI21_X1  g454(.A(KEYINPUT70), .B1(new_n645_), .B2(new_n646_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n647_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  XOR2_X1   g456(.A(G127gat), .B(G155gat), .Z(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n658_), .B(new_n659_), .ZN(new_n660_));
  XOR2_X1   g459(.A(G183gat), .B(G211gat), .Z(new_n661_));
  XNOR2_X1  g460(.A(new_n660_), .B(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT17), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(G231gat), .A2(G233gat), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT75), .Z(new_n666_));
  XNOR2_X1  g465(.A(new_n517_), .B(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n593_), .B(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n668_), .A2(KEYINPUT17), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n664_), .B1(new_n669_), .B2(new_n662_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n668_), .A2(KEYINPUT77), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n671_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n657_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n622_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n677_), .A2(new_n572_), .A3(new_n423_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT38), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT104), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n653_), .A2(new_n654_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n674_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n622_), .A2(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G1gat), .B1(new_n684_), .B2(new_n453_), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n681_), .B(new_n685_), .C1(new_n679_), .C2(new_n678_), .ZN(G1324gat));
  OAI21_X1  g485(.A(G8gat), .B1(new_n684_), .B2(new_n318_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT39), .ZN(new_n688_));
  INV_X1    g487(.A(new_n318_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n677_), .A2(new_n564_), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g491(.A(new_n458_), .ZN(new_n693_));
  OAI21_X1  g492(.A(G15gat), .B1(new_n684_), .B2(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT41), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n676_), .A2(G15gat), .A3(new_n693_), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1326gat));
  OAI21_X1  g496(.A(G22gat), .B1(new_n684_), .B2(new_n396_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT42), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n396_), .A2(G22gat), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n699_), .B1(new_n676_), .B2(new_n700_), .ZN(G1327gat));
  INV_X1    g500(.A(new_n674_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n682_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n622_), .A2(new_n704_), .ZN(new_n705_));
  OR3_X1    g504(.A1(new_n705_), .A2(G29gat), .A3(new_n453_), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n318_), .A2(new_n396_), .A3(new_n438_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n443_), .A2(new_n318_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n456_), .A2(new_n396_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n707_), .B1(new_n710_), .B2(new_n693_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n657_), .ZN(new_n712_));
  OAI21_X1  g511(.A(KEYINPUT43), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT43), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n459_), .A2(new_n714_), .A3(new_n657_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n713_), .A2(KEYINPUT105), .A3(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n621_), .A2(new_n674_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT105), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n716_), .A2(new_n717_), .A3(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n717_), .B1(new_n716_), .B2(new_n719_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n423_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n722_), .A2(KEYINPUT106), .A3(G29gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(KEYINPUT106), .B1(new_n722_), .B2(G29gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n706_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT107), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n727_), .B(new_n706_), .C1(new_n723_), .C2(new_n724_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1328gat));
  NOR3_X1   g528(.A1(new_n705_), .A2(G36gat), .A3(new_n318_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT45), .ZN(new_n731_));
  INV_X1    g530(.A(new_n721_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n716_), .A2(new_n717_), .A3(new_n719_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(new_n689_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n731_), .B1(new_n735_), .B2(G36gat), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT46), .ZN(G1329gat));
  INV_X1    g536(.A(new_n705_), .ZN(new_n738_));
  AOI21_X1  g537(.A(G43gat), .B1(new_n738_), .B2(new_n458_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n458_), .A2(G43gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n734_), .B2(new_n740_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT47), .Z(G1330gat));
  OR3_X1    g541(.A1(new_n705_), .A2(G50gat), .A3(new_n396_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n396_), .ZN(new_n744_));
  AOI21_X1  g543(.A(KEYINPUT108), .B1(new_n734_), .B2(new_n744_), .ZN(new_n745_));
  OAI211_X1 g544(.A(KEYINPUT108), .B(new_n744_), .C1(new_n720_), .C2(new_n721_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(G50gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n743_), .B1(new_n745_), .B2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT109), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT109), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n750_), .B(new_n743_), .C1(new_n745_), .C2(new_n747_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(G1331gat));
  INV_X1    g551(.A(new_n552_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n616_), .A2(new_n620_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n459_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n683_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n757_), .A2(new_n468_), .A3(new_n453_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT110), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n756_), .A2(new_n675_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(G57gat), .B1(new_n761_), .B2(new_n423_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n759_), .A2(new_n762_), .ZN(G1332gat));
  OAI21_X1  g562(.A(G64gat), .B1(new_n757_), .B2(new_n318_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT48), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n761_), .A2(new_n466_), .A3(new_n689_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n767_), .B(KEYINPUT111), .Z(G1333gat));
  OAI21_X1  g567(.A(G71gat), .B1(new_n757_), .B2(new_n693_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT49), .ZN(new_n770_));
  OR2_X1    g569(.A1(new_n693_), .A2(G71gat), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n760_), .B2(new_n771_), .ZN(G1334gat));
  OAI21_X1  g571(.A(G78gat), .B1(new_n757_), .B2(new_n396_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT50), .ZN(new_n774_));
  OR2_X1    g573(.A1(new_n396_), .A2(G78gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n760_), .B2(new_n775_), .ZN(G1335gat));
  NAND2_X1  g575(.A1(new_n755_), .A2(new_n674_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n777_), .B1(new_n713_), .B2(new_n715_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n485_), .B1(new_n778_), .B2(new_n423_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n756_), .A2(new_n704_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n780_), .A2(G85gat), .A3(new_n453_), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1336gat));
  AOI21_X1  g581(.A(new_n486_), .B1(new_n778_), .B2(new_n689_), .ZN(new_n783_));
  NOR3_X1   g582(.A1(new_n780_), .A2(G92gat), .A3(new_n318_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  XOR2_X1   g584(.A(new_n785_), .B(KEYINPUT112), .Z(G1337gat));
  AOI21_X1  g585(.A(new_n494_), .B1(new_n778_), .B2(new_n458_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n780_), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n458_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n787_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  XOR2_X1   g589(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n791_));
  XNOR2_X1  g590(.A(new_n790_), .B(new_n791_), .ZN(G1338gat));
  NAND2_X1  g591(.A1(new_n778_), .A2(new_n744_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT114), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(new_n794_), .A3(G106gat), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT52), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n794_), .B1(new_n793_), .B2(G106gat), .ZN(new_n797_));
  OR2_X1    g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n797_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n788_), .A2(new_n495_), .A3(new_n744_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n798_), .A2(new_n799_), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT53), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n798_), .A2(new_n803_), .A3(new_n799_), .A4(new_n800_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(G1339gat));
  AOI21_X1  g604(.A(new_n615_), .B1(new_n598_), .B2(new_n611_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n607_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT118), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  OAI211_X1 g608(.A(KEYINPUT118), .B(new_n607_), .C1(new_n609_), .C2(new_n610_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(new_n597_), .A3(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n592_), .A2(new_n596_), .A3(new_n594_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n812_), .A2(new_n615_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n806_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n535_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n541_), .A2(KEYINPUT55), .ZN(new_n818_));
  OAI21_X1  g617(.A(KEYINPUT115), .B1(new_n533_), .B2(new_n534_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n820_), .B(new_n536_), .C1(new_n540_), .C2(new_n516_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n817_), .A2(new_n818_), .A3(new_n819_), .A4(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n815_), .B1(new_n822_), .B2(new_n464_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n823_), .A2(new_n543_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n819_), .A2(new_n821_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT55), .B1(new_n533_), .B2(new_n534_), .ZN(new_n826_));
  NOR4_X1   g625(.A1(new_n540_), .A2(new_n516_), .A3(new_n816_), .A4(new_n536_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n465_), .B1(new_n825_), .B2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n815_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n814_), .A2(new_n824_), .A3(KEYINPUT58), .A4(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n822_), .A2(new_n815_), .A3(new_n464_), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n834_), .A2(new_n823_), .A3(new_n543_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n835_), .A2(KEYINPUT119), .A3(KEYINPUT58), .A4(new_n814_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT58), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n822_), .A2(new_n464_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT56), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n830_), .A2(new_n839_), .A3(new_n545_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n811_), .A2(new_n813_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n620_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n837_), .B1(new_n840_), .B2(new_n842_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n833_), .A2(new_n657_), .A3(new_n836_), .A4(new_n843_), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n548_), .A2(new_n841_), .A3(new_n620_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n815_), .B1(new_n829_), .B2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n543_), .B1(new_n616_), .B2(new_n620_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n838_), .A2(KEYINPUT116), .A3(KEYINPUT56), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n847_), .A2(new_n848_), .A3(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n845_), .B1(new_n850_), .B2(KEYINPUT117), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n847_), .A2(new_n848_), .A3(new_n849_), .A4(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n682_), .B1(new_n851_), .B2(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n844_), .B1(new_n854_), .B2(KEYINPUT57), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n856_));
  AOI211_X1 g655(.A(new_n856_), .B(new_n682_), .C1(new_n851_), .C2(new_n853_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n674_), .B1(new_n855_), .B2(new_n857_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n550_), .A2(new_n616_), .A3(new_n620_), .A4(new_n551_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n657_), .A2(new_n859_), .A3(new_n674_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n860_), .B(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n693_), .B1(new_n858_), .B2(new_n862_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n863_), .A2(new_n423_), .A3(new_n396_), .A4(new_n318_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT59), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n864_), .A2(new_n867_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n866_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n754_), .A2(G113gat), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(G113gat), .B1(new_n865_), .B2(new_n754_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n872_), .A2(new_n873_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n871_), .A2(new_n874_), .A3(new_n875_), .ZN(G1340gat));
  NOR2_X1   g675(.A1(new_n753_), .A2(KEYINPUT60), .ZN(new_n877_));
  MUX2_X1   g676(.A(new_n877_), .B(KEYINPUT60), .S(G120gat), .Z(new_n878_));
  NAND2_X1  g677(.A1(new_n865_), .A2(new_n878_), .ZN(new_n879_));
  XOR2_X1   g678(.A(new_n879_), .B(KEYINPUT121), .Z(new_n880_));
  AOI21_X1  g679(.A(new_n753_), .B1(new_n866_), .B2(new_n868_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT122), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(G120gat), .B1(new_n881_), .B2(new_n882_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n880_), .B1(new_n883_), .B2(new_n884_), .ZN(G1341gat));
  OAI21_X1  g684(.A(G127gat), .B1(new_n869_), .B2(new_n674_), .ZN(new_n886_));
  OR3_X1    g685(.A1(new_n864_), .A2(G127gat), .A3(new_n674_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1342gat));
  INV_X1    g687(.A(G134gat), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n869_), .A2(new_n889_), .A3(new_n712_), .ZN(new_n890_));
  AOI211_X1 g689(.A(KEYINPUT123), .B(G134gat), .C1(new_n865_), .C2(new_n682_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n865_), .A2(new_n682_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n889_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n890_), .A2(new_n891_), .A3(new_n894_), .ZN(G1343gat));
  AOI21_X1  g694(.A(new_n458_), .B1(new_n858_), .B2(new_n862_), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n689_), .A2(new_n453_), .A3(new_n396_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n754_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n552_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g702(.A1(new_n898_), .A2(new_n674_), .ZN(new_n904_));
  XOR2_X1   g703(.A(KEYINPUT61), .B(G155gat), .Z(new_n905_));
  XNOR2_X1  g704(.A(new_n904_), .B(new_n905_), .ZN(G1346gat));
  OAI21_X1  g705(.A(G162gat), .B1(new_n898_), .B2(new_n712_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n682_), .A2(new_n329_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n898_), .B2(new_n908_), .ZN(G1347gat));
  NAND2_X1  g708(.A1(new_n858_), .A2(new_n862_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n318_), .A2(new_n744_), .A3(new_n423_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n910_), .A2(new_n458_), .A3(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n228_), .B1(new_n913_), .B2(new_n754_), .ZN(new_n914_));
  XOR2_X1   g713(.A(new_n914_), .B(KEYINPUT62), .Z(new_n915_));
  NAND2_X1  g714(.A1(new_n912_), .A2(KEYINPUT124), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n863_), .A2(new_n917_), .A3(new_n911_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n916_), .A2(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n920_));
  AND2_X1   g719(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n921_));
  OAI211_X1 g720(.A(new_n919_), .B(new_n754_), .C1(new_n920_), .C2(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n915_), .A2(new_n922_), .ZN(G1348gat));
  NAND3_X1  g722(.A1(new_n919_), .A2(new_n229_), .A3(new_n552_), .ZN(new_n924_));
  OAI21_X1  g723(.A(G176gat), .B1(new_n912_), .B2(new_n753_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(G1349gat));
  AOI21_X1  g725(.A(G183gat), .B1(new_n913_), .B2(new_n702_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n674_), .A2(new_n223_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n927_), .B1(new_n919_), .B2(new_n928_), .ZN(G1350gat));
  NAND3_X1  g728(.A1(new_n919_), .A2(new_n682_), .A3(new_n256_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n712_), .B1(new_n916_), .B2(new_n918_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n931_), .A2(KEYINPUT125), .A3(new_n203_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT125), .ZN(new_n933_));
  AND4_X1   g732(.A1(new_n917_), .A2(new_n910_), .A3(new_n458_), .A4(new_n911_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n917_), .B1(new_n863_), .B2(new_n911_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n657_), .B1(new_n934_), .B2(new_n935_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n933_), .B1(new_n936_), .B2(G190gat), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n930_), .B1(new_n932_), .B2(new_n937_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  OAI211_X1 g739(.A(KEYINPUT126), .B(new_n930_), .C1(new_n932_), .C2(new_n937_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(G1351gat));
  NOR3_X1   g741(.A1(new_n318_), .A2(new_n396_), .A3(new_n423_), .ZN(new_n943_));
  AND2_X1   g742(.A1(new_n896_), .A2(new_n943_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(new_n754_), .ZN(new_n945_));
  INV_X1    g744(.A(G197gat), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n945_), .A2(KEYINPUT127), .A3(new_n946_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n944_), .A2(G197gat), .A3(new_n754_), .ZN(new_n948_));
  AND2_X1   g747(.A1(new_n948_), .A2(KEYINPUT127), .ZN(new_n949_));
  AOI211_X1 g748(.A(new_n947_), .B(new_n949_), .C1(new_n946_), .C2(new_n945_), .ZN(G1352gat));
  NAND2_X1  g749(.A1(new_n944_), .A2(new_n552_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n951_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g751(.A1(new_n944_), .A2(new_n702_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n954_));
  AND2_X1   g753(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n955_));
  NOR3_X1   g754(.A1(new_n953_), .A2(new_n954_), .A3(new_n955_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n956_), .B1(new_n953_), .B2(new_n954_), .ZN(G1354gat));
  INV_X1    g756(.A(new_n944_), .ZN(new_n958_));
  OAI21_X1  g757(.A(G218gat), .B1(new_n958_), .B2(new_n712_), .ZN(new_n959_));
  OR2_X1    g758(.A1(new_n703_), .A2(G218gat), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n959_), .B1(new_n958_), .B2(new_n960_), .ZN(G1355gat));
endmodule


