//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n867_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n906_,
    new_n907_, new_n908_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G64gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(KEYINPUT11), .ZN(new_n205_));
  XOR2_X1   g004(.A(G71gat), .B(G78gat), .Z(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n205_), .A2(new_n206_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT12), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G85gat), .A2(G92gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G85gat), .A2(G92gat), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT8), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT7), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n219_), .B(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G99gat), .A2(G106gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT6), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT67), .B1(new_n221_), .B2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n219_), .B(KEYINPUT7), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT67), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n222_), .B(KEYINPUT6), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n218_), .B1(new_n225_), .B2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT69), .ZN(new_n232_));
  OR2_X1    g031(.A1(KEYINPUT68), .A2(KEYINPUT6), .ZN(new_n233_));
  NAND2_X1  g032(.A1(KEYINPUT68), .A2(KEYINPUT6), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(new_n222_), .A3(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n222_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n232_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n237_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n239_), .A2(KEYINPUT69), .A3(new_n235_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n238_), .A2(new_n240_), .A3(new_n226_), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n241_), .A2(new_n216_), .ZN(new_n242_));
  OAI211_X1 g041(.A(KEYINPUT71), .B(new_n231_), .C1(new_n242_), .C2(new_n217_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT71), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n217_), .B1(new_n241_), .B2(new_n216_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n244_), .B1(new_n245_), .B2(new_n230_), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT10), .B(G99gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT65), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n249_), .A2(G106gat), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT9), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n215_), .A2(KEYINPUT66), .A3(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(KEYINPUT66), .B1(new_n215_), .B2(new_n251_), .ZN(new_n253_));
  OAI221_X1 g052(.A(new_n214_), .B1(new_n251_), .B2(new_n215_), .C1(new_n252_), .C2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n250_), .A2(new_n254_), .A3(new_n228_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n202_), .B(new_n212_), .C1(new_n247_), .C2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n231_), .B1(new_n242_), .B2(new_n217_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(new_n209_), .A3(new_n255_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G230gat), .A2(G233gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT64), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n256_), .B1(new_n243_), .B2(new_n246_), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT72), .B1(new_n264_), .B2(new_n211_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n258_), .A2(new_n255_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(new_n210_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT12), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n257_), .A2(new_n263_), .A3(new_n265_), .A4(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n267_), .A2(new_n271_), .A3(new_n259_), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n272_), .B(new_n262_), .C1(new_n271_), .C2(new_n267_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(G120gat), .B(G148gat), .Z(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G176gat), .B(G204gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n274_), .A2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n270_), .A2(new_n273_), .A3(new_n279_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(KEYINPUT74), .B(KEYINPUT13), .Z(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT13), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n281_), .B(new_n282_), .C1(KEYINPUT74), .C2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT75), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT75), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n285_), .A2(new_n290_), .A3(new_n287_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(KEYINPUT80), .B(G1gat), .Z(new_n293_));
  INV_X1    g092(.A(G8gat), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT14), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G15gat), .B(G22gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G1gat), .B(G8gat), .ZN(new_n298_));
  XOR2_X1   g097(.A(new_n297_), .B(new_n298_), .Z(new_n299_));
  XNOR2_X1  g098(.A(G29gat), .B(G36gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G43gat), .B(G50gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(new_n302_), .B(KEYINPUT84), .Z(new_n303_));
  XNOR2_X1  g102(.A(new_n299_), .B(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G229gat), .A2(G233gat), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n302_), .B(KEYINPUT15), .Z(new_n307_));
  OR2_X1    g106(.A1(new_n299_), .A2(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n306_), .B1(new_n299_), .B2(new_n303_), .ZN(new_n309_));
  AOI22_X1  g108(.A1(new_n304_), .A2(new_n306_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(G113gat), .B(G141gat), .Z(new_n311_));
  XNOR2_X1  g110(.A(G169gat), .B(G197gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n310_), .B(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n292_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT85), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT85), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(G169gat), .A3(G176gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT86), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n321_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT86), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n323_), .A2(new_n324_), .A3(new_n317_), .A4(new_n319_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT25), .B(G183gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT26), .B(G190gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NOR3_X1   g127(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G183gat), .A2(G190gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT23), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT23), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(G183gat), .A3(G190gat), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n329_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n322_), .A2(new_n325_), .A3(new_n328_), .A4(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(G176gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT22), .B(G169gat), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n320_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(G183gat), .A2(G190gat), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n339_), .B1(new_n332_), .B2(new_n330_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n340_), .B1(new_n332_), .B2(new_n330_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n335_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT87), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n335_), .A2(KEYINPUT87), .A3(new_n342_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G71gat), .B(G99gat), .ZN(new_n348_));
  INV_X1    g147(.A(G43gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n347_), .B(new_n350_), .Z(new_n351_));
  XOR2_X1   g150(.A(G127gat), .B(G134gat), .Z(new_n352_));
  XOR2_X1   g151(.A(G113gat), .B(G120gat), .Z(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n351_), .B(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G227gat), .A2(G233gat), .ZN(new_n357_));
  INV_X1    g156(.A(G15gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT30), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT31), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n356_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n351_), .B(new_n354_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n361_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n362_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(G155gat), .A2(G162gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT88), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G155gat), .A2(G162gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(G141gat), .ZN(new_n372_));
  INV_X1    g171(.A(G148gat), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(new_n373_), .A3(KEYINPUT3), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT3), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n375_), .B1(G141gat), .B2(G148gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G141gat), .A2(G148gat), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT89), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT2), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT2), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n378_), .A2(new_n379_), .A3(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n377_), .A2(new_n381_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT90), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT90), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n377_), .A2(new_n381_), .A3(new_n386_), .A4(new_n383_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n371_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n372_), .A2(new_n373_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n378_), .ZN(new_n390_));
  XOR2_X1   g189(.A(new_n370_), .B(KEYINPUT1), .Z(new_n391_));
  AOI21_X1  g190(.A(new_n390_), .B1(new_n391_), .B2(new_n369_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n355_), .B1(new_n388_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n371_), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n378_), .A2(new_n379_), .A3(new_n382_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n382_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n386_), .B1(new_n397_), .B2(new_n377_), .ZN(new_n398_));
  AND4_X1   g197(.A1(new_n386_), .A2(new_n377_), .A3(new_n381_), .A4(new_n383_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n394_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n392_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n400_), .A2(new_n354_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G225gat), .A2(G233gat), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n393_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G1gat), .B(G29gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(G85gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT0), .B(G57gat), .ZN(new_n407_));
  XOR2_X1   g206(.A(new_n406_), .B(new_n407_), .Z(new_n408_));
  INV_X1    g207(.A(KEYINPUT4), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n409_), .B(new_n355_), .C1(new_n388_), .C2(new_n392_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT97), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n393_), .A2(new_n402_), .A3(KEYINPUT4), .ZN(new_n412_));
  INV_X1    g211(.A(new_n403_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n404_), .B(new_n408_), .C1(new_n411_), .C2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT97), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n410_), .A2(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n410_), .A2(new_n417_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n413_), .B(new_n412_), .C1(new_n418_), .C2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n408_), .B1(new_n420_), .B2(new_n404_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n416_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n367_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT27), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G226gat), .A2(G233gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT19), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  AOI22_X1  g226(.A1(new_n326_), .A2(new_n327_), .B1(new_n323_), .B2(new_n316_), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n428_), .A2(KEYINPUT95), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n334_), .B1(new_n428_), .B2(KEYINPUT95), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n342_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(G197gat), .A2(G204gat), .ZN(new_n432_));
  INV_X1    g231(.A(G197gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT91), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT91), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(G197gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n432_), .B1(new_n437_), .B2(G204gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G211gat), .B(G218gat), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT21), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n438_), .A2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n438_), .A2(KEYINPUT21), .ZN(new_n443_));
  INV_X1    g242(.A(G204gat), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n434_), .A2(new_n436_), .A3(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n440_), .B1(G197gat), .B2(G204gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n439_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n442_), .B1(new_n443_), .B2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT20), .B1(new_n431_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(KEYINPUT96), .B1(new_n347_), .B2(new_n449_), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n335_), .A2(KEYINPUT87), .A3(new_n342_), .ZN(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT87), .B1(new_n335_), .B2(new_n342_), .ZN(new_n454_));
  OAI211_X1 g253(.A(KEYINPUT96), .B(new_n449_), .C1(new_n453_), .C2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n427_), .B(new_n451_), .C1(new_n452_), .C2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G8gat), .B(G36gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT18), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G64gat), .B(G92gat), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n459_), .B(new_n460_), .Z(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT91), .B(G197gat), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n462_), .A2(new_n444_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n440_), .B1(new_n463_), .B2(new_n432_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n439_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n465_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n466_));
  AOI22_X1  g265(.A1(new_n464_), .A2(new_n466_), .B1(new_n438_), .B2(new_n441_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n345_), .A2(new_n346_), .A3(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT20), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n469_), .B1(new_n431_), .B2(new_n449_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n427_), .B1(new_n468_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n457_), .A2(new_n461_), .A3(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n461_), .B1(new_n457_), .B2(new_n472_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n424_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n457_), .A2(new_n461_), .A3(new_n472_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n468_), .A2(new_n470_), .A3(new_n427_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n451_), .B1(new_n452_), .B2(new_n456_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n478_), .B1(new_n479_), .B2(new_n426_), .ZN(new_n480_));
  OAI211_X1 g279(.A(KEYINPUT27), .B(new_n476_), .C1(new_n480_), .C2(new_n461_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n475_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G78gat), .B(G106gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G228gat), .A2(G233gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n485_), .B1(new_n388_), .B2(new_n392_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n484_), .B1(new_n486_), .B2(new_n449_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n449_), .A2(new_n484_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n400_), .A2(new_n401_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n488_), .B1(KEYINPUT29), .B2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n483_), .B1(new_n487_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n484_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n467_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n385_), .A2(new_n387_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n392_), .B1(new_n494_), .B2(new_n394_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT29), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n493_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n483_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n467_), .B1(new_n489_), .B2(new_n485_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n497_), .B(new_n498_), .C1(new_n499_), .C2(new_n484_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n491_), .A2(new_n500_), .A3(KEYINPUT93), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n487_), .A2(new_n490_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT93), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(new_n503_), .A3(new_n498_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G22gat), .B(G50gat), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT28), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n507_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n508_));
  NOR4_X1   g307(.A1(new_n388_), .A2(KEYINPUT28), .A3(KEYINPUT29), .A4(new_n392_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n506_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n400_), .A2(new_n496_), .A3(new_n401_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT28), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n495_), .A2(new_n507_), .A3(new_n496_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(new_n513_), .A3(new_n505_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n510_), .A2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n501_), .A2(new_n504_), .A3(new_n515_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n491_), .A2(new_n500_), .A3(new_n514_), .A4(new_n510_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT94), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NOR3_X1   g318(.A1(new_n508_), .A2(new_n509_), .A3(new_n506_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n505_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n522_), .A2(KEYINPUT94), .A3(new_n500_), .A4(new_n491_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n516_), .A2(new_n519_), .A3(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n482_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT101), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT101), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n527_), .B1(new_n482_), .B2(new_n524_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n423_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n524_), .A2(new_n422_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n461_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n449_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT96), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  AOI211_X1 g333(.A(new_n426_), .B(new_n450_), .C1(new_n534_), .C2(new_n455_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n531_), .B1(new_n535_), .B2(new_n471_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(new_n476_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n450_), .B1(new_n534_), .B2(new_n455_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n471_), .B1(new_n538_), .B2(new_n427_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n424_), .B1(new_n539_), .B2(new_n461_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n477_), .B1(new_n538_), .B2(new_n427_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n531_), .ZN(new_n542_));
  AOI22_X1  g341(.A1(new_n537_), .A2(new_n424_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT100), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n530_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n475_), .A2(new_n524_), .A3(new_n481_), .A4(new_n422_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT100), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n461_), .A2(KEYINPUT32), .ZN(new_n549_));
  OAI21_X1  g348(.A(KEYINPUT98), .B1(new_n480_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n420_), .A2(new_n404_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n408_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(new_n415_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT98), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n541_), .A2(new_n555_), .A3(KEYINPUT32), .A4(new_n461_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n539_), .A2(new_n549_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n550_), .A2(new_n554_), .A3(new_n556_), .A4(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n415_), .A2(KEYINPUT33), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT33), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n420_), .A2(new_n560_), .A3(new_n404_), .A4(new_n408_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n393_), .A2(new_n402_), .A3(new_n413_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n412_), .A2(new_n403_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n552_), .B(new_n563_), .C1(new_n411_), .C2(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n562_), .A2(new_n476_), .A3(new_n536_), .A4(new_n565_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n558_), .A2(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT99), .B1(new_n567_), .B2(new_n524_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n524_), .B1(new_n558_), .B2(new_n566_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT99), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n548_), .A2(new_n568_), .A3(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n529_), .B1(new_n572_), .B2(new_n366_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n315_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G231gat), .A2(G233gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n209_), .B(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n576_), .B(new_n299_), .Z(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT82), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n578_), .B(KEYINPUT83), .Z(new_n579_));
  INV_X1    g378(.A(KEYINPUT17), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n577_), .A2(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(G127gat), .B(G155gat), .Z(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G183gat), .B(G211gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n581_), .A2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n587_), .B1(KEYINPUT17), .B2(new_n586_), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n579_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n579_), .A2(new_n588_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n264_), .A2(new_n307_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G232gat), .A2(G233gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT34), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT35), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n595_), .A2(new_n596_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n302_), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n598_), .B(new_n599_), .C1(new_n266_), .C2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT77), .ZN(new_n602_));
  OR3_X1    g401(.A1(new_n592_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n602_), .B1(new_n592_), .B2(new_n601_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G190gat), .B(G218gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G134gat), .B(G162gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n608_), .A2(KEYINPUT36), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n599_), .B1(new_n266_), .B2(new_n600_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT76), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT76), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n612_), .B(new_n599_), .C1(new_n266_), .C2(new_n600_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n597_), .B1(new_n614_), .B2(new_n592_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n605_), .A2(new_n609_), .A3(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n608_), .B(KEYINPUT36), .Z(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT78), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT79), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n619_), .B1(new_n605_), .B2(new_n615_), .ZN(new_n620_));
  OAI21_X1  g419(.A(KEYINPUT37), .B1(new_n616_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT37), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n605_), .A2(new_n609_), .A3(new_n615_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n605_), .A2(new_n615_), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n622_), .B(new_n623_), .C1(new_n624_), .C2(new_n618_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n591_), .B1(new_n621_), .B2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n574_), .A2(new_n626_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n627_), .A2(KEYINPUT102), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(KEYINPUT102), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n628_), .A2(new_n293_), .A3(new_n554_), .A4(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT38), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n545_), .B(new_n547_), .C1(new_n569_), .C2(new_n570_), .ZN(new_n633_));
  AOI211_X1 g432(.A(KEYINPUT99), .B(new_n524_), .C1(new_n558_), .C2(new_n566_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n366_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n529_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n623_), .B1(new_n624_), .B2(new_n618_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n639_), .A2(new_n591_), .A3(new_n315_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(new_n554_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(G1gat), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n630_), .A2(new_n631_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n632_), .A2(new_n642_), .A3(new_n643_), .ZN(G1324gat));
  NAND4_X1  g443(.A1(new_n628_), .A2(new_n294_), .A3(new_n482_), .A4(new_n629_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n640_), .A2(new_n482_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n646_), .B1(new_n647_), .B2(G8gat), .ZN(new_n648_));
  AOI211_X1 g447(.A(KEYINPUT39), .B(new_n294_), .C1(new_n640_), .C2(new_n482_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n645_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT40), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(G1325gat));
  INV_X1    g451(.A(new_n627_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n653_), .A2(new_n358_), .A3(new_n367_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n640_), .A2(new_n367_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n655_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n656_));
  AOI21_X1  g455(.A(KEYINPUT41), .B1(new_n655_), .B2(G15gat), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n654_), .B1(new_n656_), .B2(new_n657_), .ZN(G1326gat));
  INV_X1    g457(.A(G22gat), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n653_), .A2(new_n659_), .A3(new_n524_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n640_), .A2(new_n524_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(G22gat), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n662_), .A2(KEYINPUT42), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(KEYINPUT42), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n660_), .B1(new_n663_), .B2(new_n664_), .ZN(G1327gat));
  INV_X1    g464(.A(new_n638_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(new_n591_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT104), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n574_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(G29gat), .B1(new_n670_), .B2(new_n554_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n292_), .A2(new_n591_), .A3(new_n314_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n625_), .A2(new_n621_), .ZN(new_n673_));
  OAI21_X1  g472(.A(KEYINPUT43), .B1(new_n573_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n675_));
  INV_X1    g474(.A(new_n673_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n637_), .A2(new_n675_), .A3(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n672_), .B1(new_n674_), .B2(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n672_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n675_), .B1(new_n637_), .B2(new_n676_), .ZN(new_n682_));
  AOI211_X1 g481(.A(KEYINPUT43), .B(new_n673_), .C1(new_n635_), .C2(new_n636_), .ZN(new_n683_));
  OAI211_X1 g482(.A(KEYINPUT44), .B(new_n681_), .C1(new_n682_), .C2(new_n683_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n680_), .A2(new_n684_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n554_), .A2(G29gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n671_), .B1(new_n685_), .B2(new_n686_), .ZN(G1328gat));
  XNOR2_X1  g486(.A(new_n482_), .B(KEYINPUT106), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n669_), .A2(G36gat), .A3(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT45), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n689_), .B(new_n690_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n684_), .B(new_n482_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n692_), .A2(KEYINPUT105), .A3(G36gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(KEYINPUT105), .B1(new_n692_), .B2(G36gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n691_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT46), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  OAI211_X1 g496(.A(new_n691_), .B(KEYINPUT46), .C1(new_n693_), .C2(new_n694_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(G1329gat));
  NAND4_X1  g498(.A1(new_n680_), .A2(G43gat), .A3(new_n367_), .A4(new_n684_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n349_), .B1(new_n669_), .B2(new_n366_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g502(.A(G50gat), .B1(new_n670_), .B2(new_n524_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n524_), .A2(G50gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n685_), .B2(new_n705_), .ZN(G1331gat));
  INV_X1    g505(.A(new_n291_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n290_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n314_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n639_), .A2(new_n711_), .A3(new_n591_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n554_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n292_), .A2(new_n314_), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n714_), .A2(new_n626_), .A3(new_n637_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n422_), .A2(G57gat), .ZN(new_n716_));
  AOI22_X1  g515(.A1(new_n713_), .A2(G57gat), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT107), .Z(G1332gat));
  INV_X1    g517(.A(G64gat), .ZN(new_n719_));
  INV_X1    g518(.A(new_n688_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n715_), .A2(new_n719_), .A3(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n712_), .A2(new_n720_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(KEYINPUT108), .B(KEYINPUT48), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n722_), .A2(G64gat), .A3(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n723_), .B1(new_n722_), .B2(G64gat), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n721_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT109), .ZN(G1333gat));
  INV_X1    g526(.A(G71gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n712_), .B2(new_n367_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT49), .Z(new_n730_));
  NAND3_X1  g529(.A1(new_n715_), .A2(new_n728_), .A3(new_n367_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1334gat));
  INV_X1    g531(.A(G78gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n712_), .B2(new_n524_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT50), .Z(new_n735_));
  NAND3_X1  g534(.A1(new_n715_), .A2(new_n733_), .A3(new_n524_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1335gat));
  NAND2_X1  g536(.A1(new_n674_), .A2(new_n677_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n591_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n711_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G85gat), .B1(new_n741_), .B2(new_n422_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n668_), .A2(new_n637_), .A3(new_n714_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT110), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n668_), .A2(new_n745_), .A3(new_n637_), .A4(new_n714_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n422_), .A2(G85gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n742_), .B1(new_n748_), .B2(new_n749_), .ZN(G1336gat));
  OAI21_X1  g549(.A(G92gat), .B1(new_n741_), .B2(new_n688_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n543_), .A2(G92gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n748_), .B2(new_n752_), .ZN(G1337gat));
  NAND3_X1  g552(.A1(new_n738_), .A2(new_n367_), .A3(new_n740_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(G99gat), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT111), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n366_), .A2(new_n249_), .ZN(new_n758_));
  AOI22_X1  g557(.A1(new_n747_), .A2(new_n758_), .B1(KEYINPUT112), .B2(KEYINPUT51), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n754_), .A2(KEYINPUT111), .A3(G99gat), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n757_), .A2(new_n759_), .A3(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT113), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n761_), .B(new_n763_), .ZN(G1338gat));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n740_), .B(new_n524_), .C1(new_n682_), .C2(new_n683_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(G106gat), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n766_), .A2(G106gat), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(KEYINPUT114), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n767_), .A2(new_n768_), .ZN(new_n773_));
  INV_X1    g572(.A(G106gat), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n747_), .A2(new_n774_), .A3(new_n524_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n771_), .A2(new_n772_), .A3(new_n773_), .A4(new_n775_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n770_), .A2(KEYINPUT114), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n777_), .A2(new_n768_), .A3(new_n767_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n773_), .A2(new_n775_), .ZN(new_n779_));
  OAI21_X1  g578(.A(KEYINPUT53), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n776_), .A2(new_n780_), .ZN(G1339gat));
  AOI21_X1  g580(.A(new_n314_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n626_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n783_), .B(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n313_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n305_), .B1(new_n299_), .B2(new_n303_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n308_), .A2(new_n787_), .ZN(new_n788_));
  AOI22_X1  g587(.A1(new_n310_), .A2(new_n313_), .B1(new_n786_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n283_), .A2(new_n789_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n264_), .A2(new_n211_), .ZN(new_n791_));
  AOI22_X1  g590(.A1(new_n791_), .A2(new_n202_), .B1(new_n268_), .B2(new_n267_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n792_), .A2(KEYINPUT55), .A3(new_n265_), .A4(new_n263_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n270_), .A2(new_n794_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n257_), .A2(new_n265_), .A3(new_n269_), .A4(new_n259_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n262_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n793_), .A2(new_n795_), .A3(new_n797_), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n798_), .A2(KEYINPUT56), .A3(new_n280_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT56), .B1(new_n798_), .B2(new_n280_), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n799_), .A2(new_n800_), .A3(KEYINPUT116), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n798_), .A2(new_n280_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT56), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(KEYINPUT116), .A3(new_n803_), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n282_), .A2(new_n314_), .A3(KEYINPUT115), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT115), .B1(new_n282_), .B2(new_n314_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n804_), .A2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n790_), .B1(new_n801_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT57), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n666_), .A2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n282_), .B(new_n789_), .C1(new_n799_), .C2(new_n800_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT58), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n673_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n802_), .A2(new_n803_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n798_), .A2(KEYINPUT56), .A3(new_n280_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n818_), .A2(KEYINPUT58), .A3(new_n282_), .A4(new_n789_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n815_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n816_), .A2(new_n821_), .A3(new_n817_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n822_), .A2(new_n804_), .A3(new_n807_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n666_), .B1(new_n823_), .B2(new_n790_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n812_), .B(new_n820_), .C1(new_n824_), .C2(KEYINPUT57), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n785_), .B1(new_n825_), .B2(new_n591_), .ZN(new_n826_));
  AOI211_X1 g625(.A(new_n366_), .B(new_n422_), .C1(new_n526_), .C2(new_n528_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(G113gat), .B1(new_n829_), .B2(new_n314_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT118), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n828_), .A2(KEYINPUT117), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT59), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n833_), .B1(new_n828_), .B2(KEYINPUT117), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n832_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n831_), .B1(new_n826_), .B2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT59), .B1(new_n826_), .B2(new_n828_), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n819_), .A2(new_n815_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n809_), .A2(new_n638_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n810_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n739_), .B1(new_n839_), .B2(new_n841_), .ZN(new_n842_));
  OAI211_X1 g641(.A(KEYINPUT118), .B(new_n835_), .C1(new_n842_), .C2(new_n785_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n837_), .A2(new_n838_), .A3(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n710_), .A2(KEYINPUT119), .ZN(new_n846_));
  MUX2_X1   g645(.A(KEYINPUT119), .B(new_n846_), .S(G113gat), .Z(new_n847_));
  AOI21_X1  g646(.A(new_n830_), .B1(new_n845_), .B2(new_n847_), .ZN(G1340gat));
  OAI21_X1  g647(.A(G120gat), .B1(new_n844_), .B2(new_n292_), .ZN(new_n849_));
  INV_X1    g648(.A(G120gat), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n850_), .B1(new_n292_), .B2(KEYINPUT60), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n829_), .B(new_n851_), .C1(KEYINPUT60), .C2(new_n850_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n849_), .A2(new_n852_), .ZN(G1341gat));
  INV_X1    g652(.A(G127gat), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n591_), .A2(new_n854_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n837_), .A2(new_n838_), .A3(new_n843_), .A4(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n826_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n857_), .A2(new_n739_), .A3(new_n827_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n854_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n856_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT120), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT120), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n856_), .A2(new_n859_), .A3(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n863_), .ZN(G1342gat));
  OAI21_X1  g663(.A(G134gat), .B1(new_n844_), .B2(new_n673_), .ZN(new_n865_));
  INV_X1    g664(.A(G134gat), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n829_), .A2(new_n866_), .A3(new_n666_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n867_), .ZN(G1343gat));
  AND3_X1   g667(.A1(new_n688_), .A2(new_n524_), .A3(new_n554_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n366_), .B(new_n869_), .C1(new_n842_), .C2(new_n785_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n870_), .A2(new_n710_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(new_n372_), .ZN(G1344gat));
  NOR2_X1   g671(.A1(new_n870_), .A2(new_n292_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(new_n373_), .ZN(G1345gat));
  NOR2_X1   g673(.A1(new_n870_), .A2(new_n591_), .ZN(new_n875_));
  XOR2_X1   g674(.A(KEYINPUT61), .B(G155gat), .Z(new_n876_));
  XNOR2_X1  g675(.A(new_n875_), .B(new_n876_), .ZN(G1346gat));
  INV_X1    g676(.A(G162gat), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n870_), .A2(new_n878_), .A3(new_n673_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n870_), .B2(new_n638_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT121), .ZN(new_n881_));
  OR2_X1    g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n881_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n879_), .B1(new_n882_), .B2(new_n883_), .ZN(G1347gat));
  NOR3_X1   g683(.A1(new_n688_), .A2(new_n524_), .A3(new_n423_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  OR3_X1    g685(.A1(new_n826_), .A2(KEYINPUT122), .A3(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT122), .B1(new_n826_), .B2(new_n886_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n889_), .A2(new_n337_), .A3(new_n314_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT62), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n857_), .A2(new_n314_), .A3(new_n885_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(G169gat), .ZN(new_n893_));
  AND3_X1   g692(.A1(new_n892_), .A2(new_n891_), .A3(G169gat), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n890_), .B1(new_n893_), .B2(new_n894_), .ZN(G1348gat));
  NAND3_X1  g694(.A1(new_n889_), .A2(new_n336_), .A3(new_n709_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n857_), .A2(new_n709_), .A3(new_n885_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(G176gat), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n896_), .A2(new_n898_), .ZN(G1349gat));
  NOR3_X1   g698(.A1(new_n826_), .A2(new_n591_), .A3(new_n886_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT123), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(G183gat), .B1(new_n900_), .B2(new_n901_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n591_), .A2(new_n326_), .ZN(new_n904_));
  AOI22_X1  g703(.A1(new_n902_), .A2(new_n903_), .B1(new_n889_), .B2(new_n904_), .ZN(G1350gat));
  NAND3_X1  g704(.A1(new_n889_), .A2(new_n666_), .A3(new_n327_), .ZN(new_n906_));
  INV_X1    g705(.A(G190gat), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n673_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n906_), .B1(new_n907_), .B2(new_n908_), .ZN(G1351gat));
  AND2_X1   g708(.A1(new_n720_), .A2(new_n530_), .ZN(new_n910_));
  OAI211_X1 g709(.A(new_n366_), .B(new_n910_), .C1(new_n842_), .C2(new_n785_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(new_n710_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(new_n433_), .ZN(G1352gat));
  INV_X1    g712(.A(KEYINPUT124), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n709_), .B1(new_n914_), .B2(new_n444_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n911_), .A2(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n444_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(KEYINPUT125), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n916_), .B(new_n918_), .ZN(G1353gat));
  NOR2_X1   g718(.A1(new_n826_), .A2(new_n367_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT127), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT63), .ZN(new_n922_));
  INV_X1    g721(.A(G211gat), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n739_), .B1(new_n922_), .B2(new_n923_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(KEYINPUT126), .ZN(new_n925_));
  NAND4_X1  g724(.A1(new_n920_), .A2(new_n921_), .A3(new_n910_), .A4(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n925_), .ZN(new_n927_));
  OAI21_X1  g726(.A(KEYINPUT127), .B1(new_n911_), .B2(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n926_), .A2(new_n928_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n929_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n930_));
  NAND4_X1  g729(.A1(new_n926_), .A2(new_n928_), .A3(new_n922_), .A4(new_n923_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1354gat));
  OAI21_X1  g731(.A(G218gat), .B1(new_n911_), .B2(new_n673_), .ZN(new_n933_));
  OR2_X1    g732(.A1(new_n638_), .A2(G218gat), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n933_), .B1(new_n911_), .B2(new_n934_), .ZN(G1355gat));
endmodule


