//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 1 0 0 1 1 0 0 0 0 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n850_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n892_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_;
  INV_X1    g000(.A(KEYINPUT20), .ZN(new_n202_));
  NOR2_X1   g001(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G169gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G183gat), .A2(G190gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n204_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G169gat), .ZN(new_n210_));
  INV_X1    g009(.A(G176gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n210_), .A2(new_n211_), .A3(KEYINPUT81), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT81), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n213_), .B1(G169gat), .B2(G176gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT82), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT24), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n218_), .B1(G169gat), .B2(G176gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n217_), .A2(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n207_), .B1(new_n218_), .B2(new_n215_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT26), .B(G190gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT92), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n223_), .B(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(KEYINPUT25), .B(G183gat), .Z(new_n226_));
  OAI21_X1  g025(.A(new_n222_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n209_), .B1(new_n221_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT89), .ZN(new_n229_));
  INV_X1    g028(.A(G197gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(new_n230_), .A3(G204gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G197gat), .B(G204gat), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  OAI211_X1 g032(.A(KEYINPUT21), .B(new_n231_), .C1(new_n233_), .C2(new_n229_), .ZN(new_n234_));
  XOR2_X1   g033(.A(G211gat), .B(G218gat), .Z(new_n235_));
  XOR2_X1   g034(.A(KEYINPUT90), .B(KEYINPUT21), .Z(new_n236_));
  AOI21_X1  g035(.A(new_n235_), .B1(new_n232_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n234_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n233_), .A2(new_n235_), .A3(KEYINPUT21), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n202_), .B1(new_n228_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n217_), .A2(new_n218_), .ZN(new_n242_));
  INV_X1    g041(.A(G190gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT26), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n226_), .B1(KEYINPUT80), .B2(new_n244_), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n223_), .A2(KEYINPUT80), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n207_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n242_), .B(new_n247_), .C1(new_n217_), .C2(new_n220_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n240_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(new_n249_), .A3(new_n209_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n241_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G226gat), .A2(G233gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT19), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n248_), .A2(new_n209_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(new_n240_), .ZN(new_n256_));
  OR2_X1    g055(.A1(new_n228_), .A2(new_n240_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n253_), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n256_), .A2(new_n257_), .A3(KEYINPUT20), .A4(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(G8gat), .B(G36gat), .Z(new_n260_));
  XNOR2_X1  g059(.A(G64gat), .B(G92gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n263_));
  XOR2_X1   g062(.A(new_n262_), .B(new_n263_), .Z(new_n264_));
  NAND3_X1  g063(.A1(new_n254_), .A2(new_n259_), .A3(new_n264_), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n265_), .A2(KEYINPUT97), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(KEYINPUT97), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT20), .B1(new_n228_), .B2(new_n240_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n249_), .B1(new_n248_), .B2(new_n209_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n253_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n270_), .B1(new_n253_), .B2(new_n251_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n264_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n266_), .A2(KEYINPUT27), .A3(new_n267_), .A4(new_n273_), .ZN(new_n274_));
  NOR3_X1   g073(.A1(new_n268_), .A2(new_n269_), .A3(new_n253_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n258_), .B1(new_n241_), .B2(new_n250_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n272_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n265_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT98), .B(KEYINPUT27), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n274_), .A2(new_n280_), .ZN(new_n281_));
  NOR3_X1   g080(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT86), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G141gat), .A2(G148gat), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n284_), .A2(KEYINPUT2), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(KEYINPUT2), .ZN(new_n286_));
  INV_X1    g085(.A(G141gat), .ZN(new_n287_));
  INV_X1    g086(.A(G148gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  AOI22_X1  g088(.A1(new_n285_), .A2(new_n286_), .B1(KEYINPUT3), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n283_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT87), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT87), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n283_), .A2(new_n293_), .A3(new_n290_), .ZN(new_n294_));
  XOR2_X1   g093(.A(G155gat), .B(G162gat), .Z(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT88), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n292_), .A2(new_n294_), .A3(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G155gat), .A2(G162gat), .ZN(new_n298_));
  NOR2_X1   g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n298_), .B1(new_n299_), .B2(KEYINPUT1), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT84), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT85), .ZN(new_n302_));
  OR3_X1    g101(.A1(new_n298_), .A2(new_n302_), .A3(KEYINPUT1), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n302_), .B1(new_n298_), .B2(KEYINPUT1), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n301_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n300_), .A2(KEYINPUT84), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n289_), .B(new_n284_), .C1(new_n305_), .C2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n297_), .A2(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n249_), .B1(new_n308_), .B2(KEYINPUT29), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G228gat), .A2(G233gat), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n309_), .B(new_n310_), .Z(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G22gat), .B(G50gat), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT28), .B1(new_n308_), .B2(KEYINPUT29), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT28), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT29), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n297_), .A2(new_n316_), .A3(new_n317_), .A4(new_n307_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n314_), .B1(new_n315_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G78gat), .B(G106gat), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n315_), .A2(new_n318_), .A3(new_n314_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n320_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n323_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n325_), .A2(new_n319_), .ZN(new_n326_));
  OR2_X1    g125(.A1(new_n322_), .A2(KEYINPUT91), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n312_), .B(new_n324_), .C1(new_n326_), .C2(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n327_), .B1(new_n320_), .B2(new_n323_), .ZN(new_n329_));
  NOR3_X1   g128(.A1(new_n325_), .A2(new_n321_), .A3(new_n319_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n311_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n281_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G225gat), .A2(G233gat), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT4), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G127gat), .B(G134gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G113gat), .B(G120gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT83), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n308_), .A2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n297_), .A2(new_n340_), .A3(new_n307_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n337_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(KEYINPUT4), .B1(new_n308_), .B2(new_n341_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n336_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT95), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n342_), .A2(new_n343_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n347_), .B1(new_n348_), .B2(new_n336_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n342_), .A2(KEYINPUT95), .A3(new_n335_), .A4(new_n343_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n346_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  XOR2_X1   g150(.A(G1gat), .B(G29gat), .Z(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT94), .B(G85gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT0), .B(G57gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n351_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n356_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n346_), .A2(new_n358_), .A3(new_n349_), .A4(new_n350_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G227gat), .A2(G233gat), .ZN(new_n361_));
  INV_X1    g160(.A(G15gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT30), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n255_), .B(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(new_n341_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G71gat), .B(G99gat), .ZN(new_n367_));
  INV_X1    g166(.A(G43gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT31), .ZN(new_n370_));
  XOR2_X1   g169(.A(new_n366_), .B(new_n370_), .Z(new_n371_));
  NOR3_X1   g170(.A1(new_n334_), .A2(new_n360_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT96), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n358_), .A2(KEYINPUT33), .ZN(new_n374_));
  OR2_X1    g173(.A1(new_n351_), .A2(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n356_), .B1(new_n348_), .B2(new_n335_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n348_), .A2(KEYINPUT4), .ZN(new_n377_));
  INV_X1    g176(.A(new_n345_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n376_), .B1(new_n379_), .B2(new_n335_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n278_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT33), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n359_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n375_), .A2(new_n381_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n264_), .A2(KEYINPUT32), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NOR3_X1   g185(.A1(new_n275_), .A2(new_n276_), .A3(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n387_), .B1(new_n271_), .B2(new_n386_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n360_), .A2(new_n388_), .ZN(new_n389_));
  AND2_X1   g188(.A1(new_n384_), .A2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n373_), .B1(new_n390_), .B2(new_n332_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n332_), .B1(new_n384_), .B2(new_n389_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT96), .ZN(new_n393_));
  INV_X1    g192(.A(new_n360_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n332_), .A2(new_n394_), .A3(new_n274_), .A4(new_n280_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n391_), .A2(new_n393_), .A3(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n372_), .B1(new_n396_), .B2(new_n371_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT74), .B(G1gat), .ZN(new_n398_));
  INV_X1    g197(.A(G8gat), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT14), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G15gat), .B(G22gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G1gat), .B(G8gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G29gat), .B(G36gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT72), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G43gat), .B(G50gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT72), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n405_), .B(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n407_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n408_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n404_), .B(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G229gat), .A2(G233gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n408_), .A2(new_n412_), .A3(KEYINPUT15), .ZN(new_n418_));
  AOI21_X1  g217(.A(KEYINPUT15), .B1(new_n408_), .B2(new_n412_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n404_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n404_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n413_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n420_), .A2(new_n423_), .A3(new_n415_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n417_), .A2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G113gat), .B(G141gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT77), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G169gat), .B(G197gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n427_), .B(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT78), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n425_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n417_), .A2(new_n424_), .A3(new_n429_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(KEYINPUT79), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT79), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n425_), .A2(new_n434_), .A3(new_n430_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n397_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT70), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT69), .ZN(new_n439_));
  INV_X1    g238(.A(G64gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(G57gat), .ZN(new_n441_));
  INV_X1    g240(.A(G57gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(G64gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n441_), .A2(new_n443_), .A3(KEYINPUT11), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT67), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G57gat), .B(G64gat), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT67), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n446_), .A2(new_n447_), .A3(KEYINPUT11), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n441_), .A2(new_n443_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT11), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  XOR2_X1   g250(.A(G71gat), .B(G78gat), .Z(new_n452_));
  AND4_X1   g251(.A1(new_n445_), .A2(new_n448_), .A3(new_n451_), .A4(new_n452_), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n445_), .A2(new_n448_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT68), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n445_), .A2(new_n448_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n451_), .A2(new_n452_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT68), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n445_), .A2(new_n448_), .A3(new_n451_), .A4(new_n452_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n455_), .A2(KEYINPUT12), .A3(new_n461_), .ZN(new_n462_));
  OR2_X1    g261(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n463_));
  INV_X1    g262(.A(G106gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT64), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT64), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(G106gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n463_), .A2(new_n465_), .A3(new_n467_), .A4(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G99gat), .A2(G106gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT6), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT6), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n472_), .A2(G99gat), .A3(G106gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G85gat), .A2(G92gat), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT9), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(G85gat), .ZN(new_n479_));
  INV_X1    g278(.A(G92gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(KEYINPUT9), .A3(new_n475_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n469_), .A2(new_n474_), .A3(new_n478_), .A4(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT65), .ZN(new_n484_));
  AOI22_X1  g283(.A1(new_n471_), .A2(new_n473_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT65), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n485_), .A2(new_n469_), .A3(new_n486_), .A4(new_n482_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n484_), .A2(new_n487_), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n481_), .A2(new_n475_), .ZN(new_n489_));
  OR3_X1    g288(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n474_), .A2(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT66), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT66), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n494_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  OAI211_X1 g295(.A(KEYINPUT8), .B(new_n489_), .C1(new_n491_), .C2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n489_), .B1(new_n491_), .B2(new_n496_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT8), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n488_), .A2(new_n497_), .A3(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n462_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G230gat), .A2(G233gat), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n488_), .A2(new_n497_), .A3(new_n500_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n458_), .A2(new_n460_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n503_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(KEYINPUT12), .B1(new_n504_), .B2(new_n505_), .ZN(new_n507_));
  NOR3_X1   g306(.A1(new_n502_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n453_), .A2(new_n454_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n501_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n504_), .A2(new_n505_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n503_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n439_), .B1(new_n508_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n506_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n507_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n504_), .A2(KEYINPUT12), .A3(new_n455_), .A4(new_n461_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n514_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n503_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n504_), .A2(new_n505_), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n484_), .A2(new_n487_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n509_), .B1(new_n520_), .B2(new_n497_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n518_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n517_), .A2(KEYINPUT69), .A3(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G120gat), .B(G148gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT5), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G176gat), .B(G204gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  AND4_X1   g327(.A1(new_n438_), .A2(new_n513_), .A3(new_n523_), .A4(new_n528_), .ZN(new_n529_));
  OAI22_X1  g328(.A1(new_n521_), .A2(KEYINPUT12), .B1(new_n462_), .B2(new_n501_), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n522_), .B(new_n527_), .C1(new_n530_), .C2(new_n506_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT70), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n522_), .B1(new_n530_), .B2(new_n506_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n527_), .B1(new_n533_), .B2(new_n439_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n532_), .B1(new_n534_), .B2(new_n523_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n529_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT13), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n536_), .A2(KEYINPUT71), .A3(new_n537_), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n537_), .A2(KEYINPUT71), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(KEYINPUT71), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n539_), .B(new_n540_), .C1(new_n529_), .C2(new_n535_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n538_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G127gat), .B(G155gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT16), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G183gat), .B(G211gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT76), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G231gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n509_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(new_n421_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n550_), .B1(new_n553_), .B2(KEYINPUT68), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n554_), .B1(KEYINPUT68), .B2(new_n553_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n553_), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n547_), .B(KEYINPUT17), .Z(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n555_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n501_), .A2(new_n422_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n504_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G232gat), .A2(G233gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT34), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n563_), .A2(KEYINPUT35), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n560_), .A2(new_n561_), .A3(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(KEYINPUT35), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G190gat), .B(G218gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT73), .ZN(new_n569_));
  XOR2_X1   g368(.A(G134gat), .B(G162gat), .Z(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT36), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n567_), .A2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n571_), .B(new_n572_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n574_), .B1(new_n567_), .B2(new_n575_), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n576_), .A2(KEYINPUT37), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(KEYINPUT37), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n559_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  AND3_X1   g378(.A1(new_n437_), .A2(new_n543_), .A3(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n580_), .A2(new_n360_), .A3(new_n398_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT38), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n576_), .A2(KEYINPUT99), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT99), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n574_), .B(new_n584_), .C1(new_n567_), .C2(new_n575_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n397_), .A2(new_n586_), .ZN(new_n587_));
  NOR3_X1   g386(.A1(new_n542_), .A2(new_n559_), .A3(new_n436_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT100), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(new_n360_), .ZN(new_n591_));
  AND3_X1   g390(.A1(new_n591_), .A2(KEYINPUT101), .A3(G1gat), .ZN(new_n592_));
  AOI21_X1  g391(.A(KEYINPUT101), .B1(new_n591_), .B2(G1gat), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n582_), .B1(new_n592_), .B2(new_n593_), .ZN(G1324gat));
  INV_X1    g393(.A(new_n281_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n580_), .A2(new_n399_), .A3(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n587_), .A2(new_n595_), .A3(new_n588_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT39), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n597_), .A2(new_n598_), .A3(G8gat), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n598_), .B1(new_n597_), .B2(G8gat), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n596_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n601_), .B(new_n602_), .Z(G1325gat));
  INV_X1    g402(.A(new_n371_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n362_), .B1(new_n590_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT41), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n606_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n580_), .A2(new_n362_), .A3(new_n604_), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n609_), .B(KEYINPUT103), .Z(new_n610_));
  NAND3_X1  g409(.A1(new_n607_), .A2(new_n608_), .A3(new_n610_), .ZN(G1326gat));
  INV_X1    g410(.A(G22gat), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n580_), .A2(new_n612_), .A3(new_n332_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n590_), .A2(new_n332_), .ZN(new_n614_));
  XOR2_X1   g413(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n615_));
  AND3_X1   g414(.A1(new_n614_), .A2(G22gat), .A3(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n615_), .B1(new_n614_), .B2(G22gat), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n613_), .B1(new_n616_), .B2(new_n617_), .ZN(G1327gat));
  INV_X1    g417(.A(new_n586_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n559_), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n542_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n437_), .A2(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(G29gat), .B1(new_n622_), .B2(new_n360_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n577_), .A2(new_n578_), .ZN(new_n624_));
  OAI21_X1  g423(.A(KEYINPUT43), .B1(new_n397_), .B2(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n395_), .B1(new_n392_), .B2(KEYINPUT96), .ZN(new_n626_));
  AOI211_X1 g425(.A(new_n373_), .B(new_n332_), .C1(new_n384_), .C2(new_n389_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n371_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n372_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT43), .ZN(new_n631_));
  INV_X1    g430(.A(new_n624_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n630_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n625_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n436_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n543_), .A2(new_n559_), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(KEYINPUT44), .B1(new_n634_), .B2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT44), .ZN(new_n639_));
  AOI211_X1 g438(.A(new_n639_), .B(new_n636_), .C1(new_n625_), .C2(new_n633_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n360_), .A2(G29gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n623_), .B1(new_n641_), .B2(new_n642_), .ZN(G1328gat));
  XNOR2_X1  g442(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(G36gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n646_), .B1(new_n641_), .B2(new_n595_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n622_), .A2(new_n646_), .A3(new_n595_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT45), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n645_), .B1(new_n647_), .B2(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n648_), .B(KEYINPUT45), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n638_), .A2(new_n640_), .A3(new_n281_), .ZN(new_n653_));
  OAI211_X1 g452(.A(new_n652_), .B(new_n644_), .C1(new_n646_), .C2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n651_), .A2(new_n654_), .ZN(G1329gat));
  AOI21_X1  g454(.A(new_n631_), .B1(new_n630_), .B2(new_n632_), .ZN(new_n656_));
  AOI211_X1 g455(.A(KEYINPUT43), .B(new_n624_), .C1(new_n628_), .C2(new_n629_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n637_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(new_n639_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n634_), .A2(KEYINPUT44), .A3(new_n637_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n371_), .A2(new_n368_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n659_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(KEYINPUT106), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT106), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n659_), .A2(new_n660_), .A3(new_n664_), .A4(new_n661_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n622_), .A2(new_n604_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(new_n368_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n663_), .A2(new_n665_), .A3(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n663_), .A2(new_n665_), .A3(new_n667_), .A4(new_n669_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1330gat));
  AOI21_X1  g472(.A(G50gat), .B1(new_n622_), .B2(new_n332_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n332_), .A2(G50gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n641_), .B2(new_n675_), .ZN(G1331gat));
  NOR2_X1   g475(.A1(new_n397_), .A2(new_n635_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n677_), .A2(new_n620_), .A3(new_n542_), .A4(new_n624_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT108), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n680_), .A2(new_n442_), .A3(new_n360_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n543_), .A2(new_n559_), .A3(new_n635_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n587_), .A2(new_n682_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n683_), .A2(new_n360_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n681_), .B1(new_n442_), .B2(new_n684_), .ZN(G1332gat));
  AOI211_X1 g484(.A(KEYINPUT48), .B(new_n440_), .C1(new_n683_), .C2(new_n595_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT48), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n683_), .A2(new_n595_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n688_), .B2(G64gat), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n595_), .A2(new_n440_), .ZN(new_n690_));
  OAI22_X1  g489(.A1(new_n686_), .A2(new_n689_), .B1(new_n679_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT109), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  OAI221_X1 g492(.A(KEYINPUT109), .B1(new_n679_), .B2(new_n690_), .C1(new_n686_), .C2(new_n689_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1333gat));
  INV_X1    g494(.A(G71gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n696_), .B1(new_n683_), .B2(new_n604_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT110), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n698_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT49), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n680_), .A2(new_n696_), .A3(new_n604_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n699_), .A2(KEYINPUT49), .A3(new_n700_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n703_), .A2(new_n704_), .A3(new_n705_), .ZN(G1334gat));
  INV_X1    g505(.A(G78gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n707_), .B1(new_n683_), .B2(new_n332_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT50), .Z(new_n709_));
  NAND3_X1  g508(.A1(new_n680_), .A2(new_n707_), .A3(new_n332_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1335gat));
  NOR3_X1   g510(.A1(new_n543_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n677_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(new_n479_), .A3(new_n360_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n543_), .A2(new_n620_), .A3(new_n635_), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n634_), .A2(KEYINPUT111), .A3(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT111), .B1(new_n634_), .B2(new_n715_), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n716_), .A2(new_n717_), .A3(new_n394_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n714_), .B1(new_n718_), .B2(new_n479_), .ZN(G1336gat));
  AOI21_X1  g518(.A(G92gat), .B1(new_n713_), .B2(new_n595_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT112), .Z(new_n721_));
  NOR2_X1   g520(.A1(new_n716_), .A2(new_n717_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n281_), .A2(new_n480_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n721_), .B1(new_n722_), .B2(new_n723_), .ZN(G1337gat));
  AND2_X1   g523(.A1(new_n463_), .A2(new_n468_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n713_), .A2(new_n604_), .A3(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT113), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n634_), .A2(new_n604_), .A3(new_n715_), .ZN(new_n728_));
  INV_X1    g527(.A(G99gat), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  OAI211_X1 g529(.A(KEYINPUT114), .B(KEYINPUT51), .C1(new_n727_), .C2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT113), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n726_), .B(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n733_), .B(new_n734_), .C1(new_n728_), .C2(new_n729_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n731_), .A2(new_n735_), .ZN(G1338gat));
  NAND3_X1  g535(.A1(new_n634_), .A2(new_n332_), .A3(new_n715_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(G106gat), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT52), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n737_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n332_), .A2(new_n465_), .A3(new_n467_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n677_), .A2(new_n712_), .A3(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT115), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n740_), .A2(new_n741_), .A3(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT53), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT53), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n740_), .A2(new_n747_), .A3(new_n741_), .A4(new_n744_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(G1339gat));
  INV_X1    g548(.A(KEYINPUT117), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n433_), .A2(new_n531_), .A3(new_n435_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT55), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n517_), .A2(new_n752_), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n514_), .A2(new_n515_), .A3(KEYINPUT55), .A4(new_n516_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n518_), .B1(new_n530_), .B2(new_n519_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n753_), .A2(new_n754_), .A3(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n528_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT56), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n756_), .A2(KEYINPUT56), .A3(new_n528_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n751_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT116), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n429_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n420_), .A2(new_n423_), .A3(new_n416_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n432_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n763_), .B1(new_n536_), .B2(new_n768_), .ZN(new_n769_));
  NOR4_X1   g568(.A1(new_n529_), .A2(new_n535_), .A3(KEYINPUT116), .A4(new_n767_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n762_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n583_), .A2(KEYINPUT57), .A3(new_n585_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n750_), .B1(new_n771_), .B2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n534_), .A2(new_n438_), .A3(new_n523_), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n513_), .A2(new_n523_), .A3(new_n528_), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n775_), .B(new_n768_), .C1(new_n776_), .C2(new_n532_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT116), .ZN(new_n778_));
  INV_X1    g577(.A(new_n535_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n779_), .A2(new_n763_), .A3(new_n775_), .A4(new_n768_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n761_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n781_), .A2(KEYINPUT117), .A3(new_n772_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n774_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT57), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n784_), .B1(new_n781_), .B2(new_n586_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n759_), .A2(new_n760_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n768_), .A2(new_n531_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT58), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n786_), .A2(KEYINPUT58), .A3(new_n787_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n632_), .A2(new_n790_), .A3(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n785_), .A2(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n559_), .B1(new_n783_), .B2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n543_), .A2(new_n579_), .A3(new_n436_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT54), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n334_), .A2(new_n394_), .A3(new_n371_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n799_), .A2(KEYINPUT59), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n797_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n802_), .B1(new_n783_), .B2(new_n793_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n771_), .A2(new_n750_), .A3(new_n773_), .ZN(new_n804_));
  OAI21_X1  g603(.A(KEYINPUT117), .B1(new_n781_), .B2(new_n772_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n806_), .A2(KEYINPUT118), .A3(new_n785_), .A4(new_n792_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n803_), .A2(new_n559_), .A3(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n799_), .B1(new_n808_), .B2(new_n796_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT59), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n635_), .B(new_n801_), .C1(new_n809_), .C2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(G113gat), .ZN(new_n812_));
  INV_X1    g611(.A(G113gat), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n809_), .A2(new_n813_), .A3(new_n635_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT119), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT119), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n812_), .A2(new_n817_), .A3(new_n814_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(G1340gat));
  OAI211_X1 g618(.A(new_n542_), .B(new_n801_), .C1(new_n809_), .C2(new_n810_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(G120gat), .ZN(new_n821_));
  INV_X1    g620(.A(G120gat), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n822_), .B1(new_n543_), .B2(KEYINPUT60), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n809_), .B(new_n823_), .C1(KEYINPUT60), .C2(new_n822_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n821_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT120), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n821_), .A2(KEYINPUT120), .A3(new_n824_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(G1341gat));
  INV_X1    g628(.A(G127gat), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n809_), .A2(new_n830_), .A3(new_n620_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n809_), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n832_), .A2(KEYINPUT59), .B1(new_n797_), .B2(new_n800_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n620_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n831_), .B1(new_n835_), .B2(new_n830_), .ZN(G1342gat));
  INV_X1    g635(.A(G134gat), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(new_n832_), .B2(new_n619_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT121), .ZN(new_n839_));
  OR2_X1    g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n839_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n624_), .A2(new_n837_), .ZN(new_n842_));
  AOI22_X1  g641(.A1(new_n840_), .A2(new_n841_), .B1(new_n833_), .B2(new_n842_), .ZN(G1343gat));
  NAND2_X1  g642(.A1(new_n808_), .A2(new_n796_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n371_), .A2(new_n332_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n595_), .A2(new_n845_), .A3(new_n394_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n847_), .A2(new_n436_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(new_n287_), .ZN(G1344gat));
  NOR2_X1   g648(.A1(new_n847_), .A2(new_n543_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(new_n288_), .ZN(G1345gat));
  NOR2_X1   g650(.A1(new_n847_), .A2(new_n559_), .ZN(new_n852_));
  XOR2_X1   g651(.A(KEYINPUT61), .B(G155gat), .Z(new_n853_));
  XNOR2_X1  g652(.A(new_n852_), .B(new_n853_), .ZN(G1346gat));
  OAI21_X1  g653(.A(G162gat), .B1(new_n847_), .B2(new_n624_), .ZN(new_n855_));
  OR2_X1    g654(.A1(new_n619_), .A2(G162gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n847_), .B2(new_n856_), .ZN(G1347gat));
  INV_X1    g656(.A(KEYINPUT22), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n595_), .A2(new_n394_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n859_), .A2(new_n332_), .A3(new_n371_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n797_), .A2(new_n858_), .A3(new_n635_), .A4(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(KEYINPUT62), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT62), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n797_), .A2(new_n863_), .A3(new_n635_), .A4(new_n860_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n210_), .B1(new_n862_), .B2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(G169gat), .B1(new_n861_), .B2(KEYINPUT62), .ZN(new_n866_));
  OR3_X1    g665(.A1(new_n865_), .A2(KEYINPUT122), .A3(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(KEYINPUT122), .B1(new_n865_), .B2(new_n866_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1348gat));
  NAND2_X1  g668(.A1(new_n844_), .A2(new_n333_), .ZN(new_n870_));
  OR2_X1    g669(.A1(new_n870_), .A2(KEYINPUT124), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n859_), .A2(new_n371_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n870_), .A2(KEYINPUT124), .ZN(new_n873_));
  AND3_X1   g672(.A1(new_n871_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n543_), .A2(new_n211_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n797_), .A2(new_n860_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n211_), .B1(new_n876_), .B2(new_n543_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT123), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n877_), .A2(new_n878_), .ZN(new_n880_));
  AOI22_X1  g679(.A1(new_n874_), .A2(new_n875_), .B1(new_n879_), .B2(new_n880_), .ZN(G1349gat));
  NAND4_X1  g680(.A1(new_n797_), .A2(new_n226_), .A3(new_n620_), .A4(new_n860_), .ZN(new_n882_));
  XOR2_X1   g681(.A(new_n882_), .B(KEYINPUT125), .Z(new_n883_));
  NAND4_X1  g682(.A1(new_n871_), .A2(new_n620_), .A3(new_n872_), .A4(new_n873_), .ZN(new_n884_));
  INV_X1    g683(.A(G183gat), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n883_), .B1(new_n884_), .B2(new_n885_), .ZN(G1350gat));
  OAI21_X1  g685(.A(G190gat), .B1(new_n876_), .B2(new_n624_), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n619_), .A2(new_n225_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n876_), .B2(new_n888_), .ZN(G1351gat));
  NOR2_X1   g688(.A1(new_n859_), .A2(new_n845_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n844_), .A2(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n436_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(new_n230_), .ZN(G1352gat));
  INV_X1    g692(.A(new_n891_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n542_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g695(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n897_));
  XOR2_X1   g696(.A(new_n897_), .B(KEYINPUT126), .Z(new_n898_));
  INV_X1    g697(.A(KEYINPUT127), .ZN(new_n899_));
  AOI22_X1  g698(.A1(new_n898_), .A2(new_n899_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n894_), .A2(new_n620_), .A3(new_n900_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n898_), .A2(new_n899_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1354gat));
  OR3_X1    g702(.A1(new_n891_), .A2(G218gat), .A3(new_n619_), .ZN(new_n904_));
  OAI21_X1  g703(.A(G218gat), .B1(new_n891_), .B2(new_n624_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1355gat));
endmodule


