//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1 0 1 1 1 0 0 1 0 0 0 0 1 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n614_, new_n615_, new_n616_, new_n617_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n832_, new_n833_, new_n834_, new_n836_, new_n837_, new_n838_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n845_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n879_, new_n880_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NOR3_X1   g004(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(G183gat), .A3(G190gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT85), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G183gat), .ZN(new_n211_));
  INV_X1    g010(.A(G190gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT23), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n206_), .B1(new_n210_), .B2(new_n213_), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n214_), .A2(KEYINPUT86), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(KEYINPUT86), .ZN(new_n216_));
  XOR2_X1   g015(.A(KEYINPUT25), .B(G183gat), .Z(new_n217_));
  NAND2_X1  g016(.A1(new_n212_), .A2(KEYINPUT26), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n217_), .B1(KEYINPUT84), .B2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT26), .B(G190gat), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n220_), .A2(KEYINPUT84), .ZN(new_n221_));
  XOR2_X1   g020(.A(G169gat), .B(G176gat), .Z(new_n222_));
  AOI22_X1  g021(.A1(new_n219_), .A2(new_n221_), .B1(KEYINPUT24), .B2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n215_), .A2(new_n216_), .A3(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(G169gat), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n213_), .A2(new_n208_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n226_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n224_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G71gat), .B(G99gat), .ZN(new_n231_));
  INV_X1    g030(.A(G43gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n230_), .A2(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n230_), .A2(new_n233_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G227gat), .A2(G233gat), .ZN(new_n236_));
  INV_X1    g035(.A(G15gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT30), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT31), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NOR3_X1   g040(.A1(new_n234_), .A2(new_n235_), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT87), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n241_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n244_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n205_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n245_), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT87), .B1(new_n250_), .B2(new_n242_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n251_), .A2(new_n246_), .A3(new_n204_), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n249_), .A2(KEYINPUT88), .A3(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(KEYINPUT88), .B1(new_n249_), .B2(new_n252_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT1), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(G155gat), .A3(G162gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT90), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT89), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G155gat), .A2(G162gat), .ZN(new_n260_));
  NOR2_X1   g059(.A1(G155gat), .A2(G162gat), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n260_), .B1(new_n261_), .B2(KEYINPUT1), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n258_), .B1(new_n259_), .B2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n263_), .B1(new_n259_), .B2(new_n262_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G141gat), .A2(G148gat), .ZN(new_n265_));
  NOR2_X1   g064(.A1(G141gat), .A2(G148gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n264_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n266_), .B(KEYINPUT3), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n265_), .B(KEYINPUT2), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n261_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(new_n260_), .A3(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n268_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT29), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(G22gat), .B(G50gat), .Z(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT28), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n277_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G78gat), .B(G106gat), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(G197gat), .B(G204gat), .Z(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT21), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G211gat), .B(G218gat), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT92), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n283_), .A2(KEYINPUT21), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n288_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(KEYINPUT91), .A2(G233gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(KEYINPUT91), .A2(G233gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(G228gat), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n290_), .B(new_n294_), .C1(new_n275_), .C2(new_n276_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n294_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n264_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n276_), .B1(new_n297_), .B2(new_n273_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n290_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n296_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n282_), .B1(new_n295_), .B2(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n280_), .B1(new_n301_), .B2(KEYINPUT93), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n295_), .A2(new_n300_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n281_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n295_), .A2(new_n300_), .A3(new_n282_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n302_), .A2(new_n306_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n304_), .A2(new_n280_), .A3(KEYINPUT93), .A4(new_n305_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n210_), .A2(new_n213_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n311_), .B1(G183gat), .B2(G190gat), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT96), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n313_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(new_n226_), .A3(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n220_), .B(KEYINPUT94), .ZN(new_n317_));
  INV_X1    g116(.A(new_n217_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(G169gat), .A2(G176gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT95), .B(KEYINPUT24), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n227_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n222_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n319_), .B(new_n322_), .C1(new_n323_), .C2(new_n321_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n316_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(new_n290_), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n326_), .B(KEYINPUT20), .C1(new_n290_), .C2(new_n230_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G226gat), .A2(G233gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT19), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G8gat), .B(G36gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT18), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G64gat), .B(G92gat), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n332_), .B(new_n333_), .Z(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT32), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n316_), .A2(new_n299_), .A3(new_n324_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n230_), .A2(new_n290_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(new_n337_), .A3(KEYINPUT20), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n338_), .A2(new_n329_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n330_), .A2(new_n335_), .A3(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(KEYINPUT97), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT97), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n330_), .A2(new_n342_), .A3(new_n339_), .A4(new_n335_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n204_), .B1(new_n268_), .B2(new_n274_), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n345_), .A2(KEYINPUT4), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n297_), .A2(new_n205_), .A3(new_n273_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n345_), .A2(KEYINPUT4), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G225gat), .A2(G233gat), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n345_), .A2(new_n347_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n353_), .A2(new_n351_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G1gat), .B(G29gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(G85gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT0), .B(G57gat), .ZN(new_n358_));
  XOR2_X1   g157(.A(new_n357_), .B(new_n358_), .Z(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n352_), .A2(new_n355_), .A3(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n350_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n359_), .B1(new_n362_), .B2(new_n354_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n335_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n338_), .A2(new_n329_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n365_), .B1(new_n327_), .B2(new_n329_), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n361_), .A2(new_n363_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n344_), .A2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n359_), .B1(new_n353_), .B2(new_n351_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n346_), .A2(new_n350_), .A3(new_n348_), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT33), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n363_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n330_), .A2(new_n334_), .A3(new_n339_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n330_), .A2(new_n339_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n334_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  OAI211_X1 g176(.A(KEYINPUT33), .B(new_n359_), .C1(new_n362_), .C2(new_n354_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n373_), .A2(new_n374_), .A3(new_n377_), .A4(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n310_), .B1(new_n368_), .B2(new_n379_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n307_), .A2(new_n363_), .A3(new_n361_), .A4(new_n308_), .ZN(new_n381_));
  AOI21_X1  g180(.A(KEYINPUT27), .B1(new_n377_), .B2(new_n374_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n366_), .A2(new_n376_), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n383_), .A2(KEYINPUT27), .A3(new_n374_), .ZN(new_n384_));
  NOR3_X1   g183(.A1(new_n381_), .A2(new_n382_), .A3(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n255_), .B1(new_n380_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n249_), .A2(new_n252_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n361_), .A2(new_n363_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n382_), .A2(new_n384_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n389_), .A2(new_n309_), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n386_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT69), .ZN(new_n393_));
  XOR2_X1   g192(.A(G85gat), .B(G92gat), .Z(new_n394_));
  INV_X1    g193(.A(KEYINPUT6), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n395_), .B1(G99gat), .B2(G106gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G99gat), .A2(G106gat), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n397_), .A2(KEYINPUT6), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT7), .ZN(new_n400_));
  INV_X1    g199(.A(G99gat), .ZN(new_n401_));
  INV_X1    g200(.A(G106gat), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n400_), .A2(new_n401_), .A3(new_n402_), .A4(KEYINPUT68), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT68), .ZN(new_n404_));
  OAI22_X1  g203(.A1(new_n404_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n393_), .B(new_n394_), .C1(new_n399_), .C2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT8), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n405_), .B(new_n403_), .C1(new_n396_), .C2(new_n398_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n393_), .B1(new_n409_), .B2(new_n394_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  AOI211_X1 g210(.A(new_n393_), .B(KEYINPUT8), .C1(new_n409_), .C2(new_n394_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT10), .B(G99gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT64), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n399_), .B1(new_n415_), .B2(new_n402_), .ZN(new_n416_));
  INV_X1    g215(.A(G85gat), .ZN(new_n417_));
  INV_X1    g216(.A(G92gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT9), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT65), .B(G85gat), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n422_), .B1(new_n423_), .B2(new_n418_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT66), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n421_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  OAI211_X1 g225(.A(KEYINPUT66), .B(new_n422_), .C1(new_n423_), .C2(new_n418_), .ZN(new_n427_));
  AOI21_X1  g226(.A(KEYINPUT67), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n417_), .A2(KEYINPUT65), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT65), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(G85gat), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n418_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n425_), .B1(new_n432_), .B2(KEYINPUT9), .ZN(new_n433_));
  INV_X1    g232(.A(new_n421_), .ZN(new_n434_));
  AND4_X1   g233(.A1(KEYINPUT67), .A2(new_n433_), .A3(new_n427_), .A4(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n416_), .B1(new_n428_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n413_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G29gat), .B(G36gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G43gat), .B(G50gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT15), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n437_), .A2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT73), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G232gat), .A2(G233gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT34), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT35), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT75), .B1(new_n445_), .B2(KEYINPUT35), .ZN(new_n447_));
  INV_X1    g246(.A(new_n437_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n447_), .B1(new_n448_), .B2(new_n440_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n443_), .A2(new_n446_), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G190gat), .B(G218gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(KEYINPUT74), .ZN(new_n453_));
  XOR2_X1   g252(.A(G134gat), .B(G162gat), .Z(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  OR2_X1    g255(.A1(new_n456_), .A2(KEYINPUT36), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n446_), .B1(new_n443_), .B2(new_n449_), .ZN(new_n458_));
  OR3_X1    g257(.A1(new_n451_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n456_), .A2(KEYINPUT36), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n457_), .B(new_n460_), .C1(new_n451_), .C2(new_n458_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n392_), .A2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G57gat), .B(G64gat), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n464_), .A2(KEYINPUT11), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(KEYINPUT11), .ZN(new_n466_));
  XOR2_X1   g265(.A(G71gat), .B(G78gat), .Z(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  OR2_X1    g267(.A1(new_n466_), .A2(new_n467_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT70), .B(KEYINPUT12), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n415_), .A2(new_n402_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n399_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n433_), .A2(new_n427_), .A3(new_n434_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT67), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n426_), .A2(KEYINPUT67), .A3(new_n427_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n475_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n410_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(KEYINPUT8), .A3(new_n407_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n412_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n471_), .B(new_n472_), .C1(new_n480_), .C2(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n470_), .B1(new_n413_), .B2(new_n436_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT12), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n487_), .A2(KEYINPUT70), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n485_), .B1(new_n486_), .B2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n413_), .A2(new_n436_), .A3(new_n470_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G230gat), .A2(G233gat), .ZN(new_n492_));
  AND3_X1   g291(.A1(new_n491_), .A2(KEYINPUT71), .A3(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(KEYINPUT71), .B1(new_n491_), .B2(new_n492_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n490_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT72), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n491_), .ZN(new_n498_));
  OAI211_X1 g297(.A(G230gat), .B(G233gat), .C1(new_n498_), .C2(new_n486_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n490_), .B(KEYINPUT72), .C1(new_n493_), .C2(new_n494_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n497_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G120gat), .B(G148gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT5), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G176gat), .B(G204gat), .ZN(new_n504_));
  XOR2_X1   g303(.A(new_n503_), .B(new_n504_), .Z(new_n505_));
  NAND2_X1  g304(.A1(new_n501_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n505_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n497_), .A2(new_n499_), .A3(new_n500_), .A4(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n506_), .A2(KEYINPUT13), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT13), .B1(new_n506_), .B2(new_n508_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G1gat), .B(G8gat), .ZN(new_n513_));
  OR2_X1    g312(.A1(new_n513_), .A2(KEYINPUT77), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(KEYINPUT77), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G15gat), .B(G22gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G1gat), .A2(G8gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT14), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n516_), .A2(new_n520_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n514_), .A2(new_n519_), .A3(new_n517_), .A4(new_n515_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(new_n440_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G229gat), .A2(G233gat), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(G113gat), .B(G141gat), .Z(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT81), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT82), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G169gat), .B(G197gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n441_), .A2(new_n522_), .A3(new_n521_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n523_), .A2(new_n440_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(new_n534_), .A3(new_n525_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n527_), .A2(new_n532_), .A3(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT83), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n527_), .A2(new_n535_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n532_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n537_), .B(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n512_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G231gat), .A2(G233gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n523_), .B(new_n543_), .ZN(new_n544_));
  XOR2_X1   g343(.A(new_n470_), .B(KEYINPUT78), .Z(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT17), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(G127gat), .B(G155gat), .Z(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT16), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G183gat), .B(G211gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n548_), .A2(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n553_), .B1(KEYINPUT17), .B2(new_n552_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n546_), .A2(KEYINPUT79), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NOR3_X1   g356(.A1(new_n463_), .A2(new_n542_), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n388_), .ZN(new_n560_));
  OAI21_X1  g359(.A(G1gat), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT38), .ZN(new_n562_));
  XNOR2_X1  g361(.A(KEYINPUT76), .B(KEYINPUT37), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n462_), .A2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n459_), .A2(new_n461_), .A3(new_n563_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n565_), .A2(new_n566_), .A3(new_n556_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT80), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n542_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n569_), .A2(new_n570_), .A3(new_n392_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT98), .ZN(new_n572_));
  INV_X1    g371(.A(new_n381_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n390_), .A2(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n360_), .B1(new_n352_), .B2(new_n355_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n372_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n378_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n377_), .A2(new_n374_), .ZN(new_n579_));
  AOI22_X1  g378(.A1(new_n578_), .A2(new_n579_), .B1(new_n344_), .B2(new_n367_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n574_), .B1(new_n580_), .B2(new_n310_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n390_), .A2(new_n309_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  AOI22_X1  g382(.A1(new_n581_), .A2(new_n255_), .B1(new_n583_), .B2(new_n389_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n584_), .A2(new_n542_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT98), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(new_n586_), .A3(new_n569_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n572_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(G1gat), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(new_n589_), .A3(new_n388_), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n590_), .A2(KEYINPUT99), .A3(new_n562_), .ZN(new_n591_));
  AOI21_X1  g390(.A(KEYINPUT99), .B1(new_n590_), .B2(new_n562_), .ZN(new_n592_));
  OAI221_X1 g391(.A(new_n561_), .B1(new_n562_), .B2(new_n590_), .C1(new_n591_), .C2(new_n592_), .ZN(G1324gat));
  NOR2_X1   g392(.A1(new_n390_), .A2(G8gat), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n572_), .A2(new_n587_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT39), .ZN(new_n596_));
  INV_X1    g395(.A(new_n390_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n542_), .A2(new_n557_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n392_), .A2(new_n597_), .A3(new_n462_), .A4(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n596_), .B1(new_n599_), .B2(G8gat), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n599_), .A2(new_n596_), .A3(G8gat), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n595_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT101), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT101), .ZN(new_n604_));
  OAI211_X1 g403(.A(new_n595_), .B(new_n604_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(G1325gat));
  INV_X1    g407(.A(new_n255_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n237_), .B1(new_n558_), .B2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT41), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n588_), .A2(new_n237_), .A3(new_n609_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(G1326gat));
  INV_X1    g412(.A(G22gat), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n614_), .B1(new_n558_), .B2(new_n310_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT42), .Z(new_n616_));
  NAND3_X1  g415(.A1(new_n588_), .A2(new_n614_), .A3(new_n310_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(G1327gat));
  NOR4_X1   g417(.A1(new_n584_), .A2(new_n542_), .A3(new_n462_), .A4(new_n556_), .ZN(new_n619_));
  AOI21_X1  g418(.A(G29gat), .B1(new_n619_), .B2(new_n388_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(KEYINPUT102), .B(KEYINPUT43), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n565_), .A2(new_n566_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n621_), .B1(new_n392_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT43), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n625_), .A2(KEYINPUT102), .ZN(new_n626_));
  AOI211_X1 g425(.A(new_n626_), .B(new_n622_), .C1(new_n386_), .C2(new_n391_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n624_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT44), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n570_), .A2(new_n557_), .ZN(new_n630_));
  NOR3_X1   g429(.A1(new_n628_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT103), .ZN(new_n632_));
  INV_X1    g431(.A(new_n621_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n633_), .B1(new_n584_), .B2(new_n622_), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n392_), .B(new_n623_), .C1(KEYINPUT102), .C2(new_n625_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n630_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n632_), .B1(new_n636_), .B2(KEYINPUT44), .ZN(new_n637_));
  OAI211_X1 g436(.A(KEYINPUT103), .B(new_n629_), .C1(new_n628_), .C2(new_n630_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n631_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n388_), .A2(G29gat), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n620_), .B1(new_n639_), .B2(new_n640_), .ZN(G1328gat));
  NOR2_X1   g440(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n642_));
  INV_X1    g441(.A(G36gat), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n643_), .B1(new_n639_), .B2(new_n597_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n619_), .A2(new_n643_), .A3(new_n597_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT45), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n642_), .B1(new_n644_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n642_), .ZN(new_n649_));
  AOI211_X1 g448(.A(new_n390_), .B(new_n631_), .C1(new_n637_), .C2(new_n638_), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n649_), .B(new_n646_), .C1(new_n650_), .C2(new_n643_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n648_), .A2(new_n651_), .ZN(G1329gat));
  NOR2_X1   g451(.A1(new_n387_), .A2(new_n232_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  AOI211_X1 g453(.A(new_n654_), .B(new_n631_), .C1(new_n637_), .C2(new_n638_), .ZN(new_n655_));
  AOI21_X1  g454(.A(G43gat), .B1(new_n619_), .B2(new_n609_), .ZN(new_n656_));
  OAI21_X1  g455(.A(KEYINPUT47), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n656_), .B1(new_n639_), .B2(new_n653_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT47), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n657_), .A2(new_n660_), .ZN(G1330gat));
  INV_X1    g460(.A(G50gat), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n310_), .A2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT105), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n619_), .A2(new_n664_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n639_), .A2(new_n310_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n666_), .B2(new_n662_), .ZN(G1331gat));
  INV_X1    g466(.A(new_n512_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n569_), .A2(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n669_), .A2(KEYINPUT106), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n670_), .A2(new_n541_), .A3(new_n584_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(KEYINPUT106), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(G57gat), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n674_), .A2(new_n675_), .A3(new_n388_), .ZN(new_n676_));
  NOR4_X1   g475(.A1(new_n463_), .A2(new_n541_), .A3(new_n512_), .A4(new_n557_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n677_), .A2(new_n388_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n676_), .B1(new_n675_), .B2(new_n678_), .ZN(G1332gat));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n677_), .A2(new_n597_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT48), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n681_), .A2(new_n682_), .A3(G64gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n682_), .B1(new_n681_), .B2(G64gat), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n390_), .A2(G64gat), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n673_), .A2(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n680_), .B1(new_n685_), .B2(new_n687_), .ZN(new_n688_));
  OAI221_X1 g487(.A(KEYINPUT107), .B1(new_n673_), .B2(new_n686_), .C1(new_n683_), .C2(new_n684_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1333gat));
  INV_X1    g489(.A(G71gat), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n674_), .A2(new_n691_), .A3(new_n609_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n691_), .B1(new_n677_), .B2(new_n609_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(KEYINPUT108), .B(KEYINPUT49), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n692_), .A2(new_n695_), .ZN(G1334gat));
  INV_X1    g495(.A(G78gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n697_), .B1(new_n677_), .B2(new_n310_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT50), .Z(new_n699_));
  NAND3_X1  g498(.A1(new_n674_), .A2(new_n697_), .A3(new_n310_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1335gat));
  NOR2_X1   g500(.A1(new_n584_), .A2(new_n541_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n512_), .A2(new_n462_), .A3(new_n556_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT109), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n702_), .A2(new_n706_), .A3(new_n703_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(G85gat), .B1(new_n708_), .B2(new_n388_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n541_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n668_), .A2(new_n710_), .A3(new_n557_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n711_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n713_), .A2(new_n423_), .A3(new_n560_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n709_), .A2(new_n714_), .ZN(G1336gat));
  NAND3_X1  g514(.A1(new_n708_), .A2(new_n418_), .A3(new_n597_), .ZN(new_n716_));
  OAI21_X1  g515(.A(G92gat), .B1(new_n713_), .B2(new_n390_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1337gat));
  INV_X1    g517(.A(new_n387_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n415_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n720_), .B1(new_n705_), .B2(new_n707_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n401_), .B1(new_n712_), .B2(new_n609_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT111), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  AND2_X1   g524(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n726_));
  OAI21_X1  g525(.A(KEYINPUT111), .B1(new_n721_), .B2(new_n722_), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n725_), .A2(new_n726_), .A3(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n726_), .B1(new_n725_), .B2(new_n727_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1338gat));
  NAND3_X1  g529(.A1(new_n708_), .A2(new_n402_), .A3(new_n310_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n712_), .A2(new_n310_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n732_), .A2(G106gat), .A3(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n732_), .B2(G106gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n731_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g536(.A(KEYINPUT120), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT54), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n739_), .A2(KEYINPUT113), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n565_), .A2(new_n710_), .A3(new_n566_), .A4(new_n556_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(KEYINPUT113), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  OR3_X1    g542(.A1(new_n741_), .A2(new_n668_), .A3(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(new_n741_), .B2(new_n668_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n740_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n508_), .A2(new_n541_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT114), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n747_), .B(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT56), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n490_), .B(KEYINPUT55), .C1(new_n493_), .C2(new_n494_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n490_), .A2(new_n491_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n752_), .B2(new_n492_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT55), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n497_), .A2(new_n754_), .A3(new_n500_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT115), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n753_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n497_), .A2(KEYINPUT115), .A3(new_n754_), .A4(new_n500_), .ZN(new_n758_));
  AOI211_X1 g557(.A(new_n750_), .B(new_n507_), .C1(new_n757_), .C2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n755_), .A2(new_n756_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n753_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(new_n758_), .A3(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(KEYINPUT56), .B1(new_n762_), .B2(new_n505_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n749_), .B1(new_n759_), .B2(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n533_), .A2(new_n534_), .A3(new_n526_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n524_), .A2(new_n525_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n539_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(new_n536_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n768_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n764_), .A2(new_n770_), .ZN(new_n771_));
  XOR2_X1   g570(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n771_), .A2(new_n462_), .A3(new_n773_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n747_), .B(KEYINPUT114), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n762_), .A2(new_n505_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n750_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n762_), .A2(KEYINPUT56), .A3(new_n505_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n775_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n462_), .B1(new_n779_), .B2(new_n769_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n768_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n508_), .A2(new_n783_), .ZN(new_n784_));
  OAI211_X1 g583(.A(KEYINPUT58), .B(new_n784_), .C1(new_n759_), .C2(new_n763_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT118), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n777_), .A2(new_n778_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n788_), .A2(KEYINPUT118), .A3(KEYINPUT58), .A4(new_n784_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n787_), .A2(new_n789_), .A3(new_n623_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(KEYINPUT117), .B(KEYINPUT58), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n784_), .B1(new_n759_), .B2(new_n763_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  OAI211_X1 g594(.A(KEYINPUT116), .B(new_n784_), .C1(new_n759_), .C2(new_n763_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n792_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n774_), .B(new_n782_), .C1(new_n790_), .C2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n746_), .B1(new_n798_), .B2(new_n557_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n582_), .A2(new_n560_), .A3(new_n387_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n738_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT116), .B1(new_n788_), .B2(new_n784_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n796_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n791_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n622_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n789_), .A3(new_n806_), .ZN(new_n807_));
  AOI22_X1  g606(.A1(new_n771_), .A2(new_n462_), .B1(KEYINPUT119), .B2(KEYINPUT57), .ZN(new_n808_));
  INV_X1    g607(.A(new_n462_), .ZN(new_n809_));
  AOI211_X1 g608(.A(new_n809_), .B(new_n772_), .C1(new_n764_), .C2(new_n770_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n808_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n556_), .B1(new_n807_), .B2(new_n811_), .ZN(new_n812_));
  OAI211_X1 g611(.A(KEYINPUT120), .B(new_n800_), .C1(new_n812_), .C2(new_n746_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n802_), .A2(new_n541_), .A3(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(G113gat), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT59), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n816_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n817_));
  OAI211_X1 g616(.A(KEYINPUT59), .B(new_n800_), .C1(new_n812_), .C2(new_n746_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n815_), .B1(new_n541_), .B2(KEYINPUT121), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n820_), .B1(KEYINPUT121), .B2(new_n815_), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n814_), .A2(new_n815_), .B1(new_n819_), .B2(new_n821_), .ZN(G1340gat));
  INV_X1    g621(.A(KEYINPUT60), .ZN(new_n823_));
  AOI21_X1  g622(.A(G120gat), .B1(new_n668_), .B2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n824_), .B1(new_n823_), .B2(G120gat), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n802_), .A2(new_n813_), .A3(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n512_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT122), .ZN(new_n828_));
  OAI21_X1  g627(.A(G120gat), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  AOI211_X1 g628(.A(KEYINPUT122), .B(new_n512_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n826_), .B1(new_n829_), .B2(new_n830_), .ZN(G1341gat));
  INV_X1    g630(.A(G127gat), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n802_), .A2(new_n813_), .A3(new_n832_), .A4(new_n556_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n557_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n833_), .B1(new_n834_), .B2(new_n832_), .ZN(G1342gat));
  INV_X1    g634(.A(G134gat), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n802_), .A2(new_n813_), .A3(new_n836_), .A4(new_n809_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n622_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(new_n838_), .B2(new_n836_), .ZN(G1343gat));
  NAND4_X1  g638(.A1(new_n255_), .A2(new_n388_), .A3(new_n310_), .A4(new_n390_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n799_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n541_), .ZN(new_n842_));
  XOR2_X1   g641(.A(KEYINPUT123), .B(G141gat), .Z(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(G1344gat));
  NAND2_X1  g643(.A1(new_n841_), .A2(new_n668_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g645(.A1(new_n841_), .A2(new_n556_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(KEYINPUT61), .B(G155gat), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n847_), .B(new_n848_), .ZN(G1346gat));
  INV_X1    g648(.A(G162gat), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n841_), .A2(new_n850_), .A3(new_n809_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n799_), .A2(new_n622_), .A3(new_n840_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT124), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n851_), .B(KEYINPUT124), .C1(new_n850_), .C2(new_n852_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(G1347gat));
  INV_X1    g656(.A(KEYINPUT62), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n255_), .A2(new_n388_), .A3(new_n310_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NOR4_X1   g659(.A1(new_n799_), .A2(new_n710_), .A3(new_n390_), .A4(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT22), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n858_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(G169gat), .ZN(new_n864_));
  INV_X1    g663(.A(G169gat), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n865_), .B1(new_n861_), .B2(new_n858_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n864_), .B1(new_n863_), .B2(new_n866_), .ZN(G1348gat));
  NOR2_X1   g666(.A1(new_n799_), .A2(new_n390_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n868_), .A2(new_n668_), .A3(new_n859_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g669(.A1(new_n868_), .A2(new_n556_), .A3(new_n859_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(new_n318_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n872_), .B1(new_n211_), .B2(new_n871_), .ZN(G1350gat));
  NAND2_X1  g672(.A1(new_n868_), .A2(new_n859_), .ZN(new_n874_));
  OAI21_X1  g673(.A(G190gat), .B1(new_n874_), .B2(new_n622_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n809_), .A2(new_n317_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(KEYINPUT125), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n875_), .B1(new_n874_), .B2(new_n877_), .ZN(G1351gat));
  NOR2_X1   g677(.A1(new_n609_), .A2(new_n381_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n868_), .A2(new_n541_), .A3(new_n879_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g680(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n882_));
  XOR2_X1   g681(.A(new_n882_), .B(KEYINPUT127), .Z(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n868_), .A2(new_n879_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n512_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n884_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  OAI221_X1 g687(.A(new_n883_), .B1(KEYINPUT126), .B2(G204gat), .C1(new_n885_), .C2(new_n512_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(G1353gat));
  XNOR2_X1  g689(.A(KEYINPUT63), .B(G211gat), .ZN(new_n891_));
  OR2_X1    g690(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n868_), .A2(new_n556_), .A3(new_n879_), .ZN(new_n893_));
  MUX2_X1   g692(.A(new_n891_), .B(new_n892_), .S(new_n893_), .Z(G1354gat));
  OAI21_X1  g693(.A(G218gat), .B1(new_n885_), .B2(new_n622_), .ZN(new_n895_));
  OR2_X1    g694(.A1(new_n462_), .A2(G218gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n885_), .B2(new_n896_), .ZN(G1355gat));
endmodule


