//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0 0 0 1 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n627_, new_n628_, new_n629_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n683_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n796_, new_n797_, new_n798_, new_n800_, new_n801_, new_n803_,
    new_n804_, new_n806_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n827_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n837_, new_n838_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_;
  XNOR2_X1  g000(.A(G71gat), .B(G78gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(G57gat), .B(G64gat), .Z(new_n203_));
  INV_X1    g002(.A(KEYINPUT11), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G57gat), .B(G64gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT11), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n202_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n208_));
  AND2_X1   g007(.A1(new_n207_), .A2(new_n202_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT67), .ZN(new_n211_));
  XOR2_X1   g010(.A(KEYINPUT10), .B(G99gat), .Z(new_n212_));
  INV_X1    g011(.A(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G92gat), .ZN(new_n215_));
  NOR3_X1   g014(.A1(new_n215_), .A2(KEYINPUT64), .A3(KEYINPUT9), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n215_), .A2(KEYINPUT64), .ZN(new_n217_));
  OAI21_X1  g016(.A(G85gat), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  AND3_X1   g017(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G85gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n222_), .A2(G92gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n215_), .A2(G85gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT9), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n214_), .A2(new_n218_), .A3(new_n221_), .A4(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT8), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NOR3_X1   g028(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G99gat), .A2(G106gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT6), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n235_));
  NAND3_X1  g034(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n234_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT66), .B1(new_n219_), .B2(new_n220_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n231_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n240_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n215_), .A2(G85gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n222_), .A2(G92gat), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n242_), .A2(new_n243_), .A3(KEYINPUT65), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n227_), .B1(new_n239_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT7), .ZN(new_n247_));
  INV_X1    g046(.A(G99gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n247_), .A2(new_n248_), .A3(new_n213_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n249_), .A2(new_n234_), .A3(new_n236_), .A4(new_n228_), .ZN(new_n250_));
  AND3_X1   g049(.A1(new_n242_), .A2(new_n243_), .A3(KEYINPUT65), .ZN(new_n251_));
  AOI21_X1  g050(.A(KEYINPUT65), .B1(new_n242_), .B2(new_n243_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n250_), .B(new_n227_), .C1(new_n251_), .C2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n226_), .B1(new_n246_), .B2(new_n254_), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n211_), .A2(new_n255_), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n255_), .B(KEYINPUT12), .C1(new_n208_), .C2(new_n209_), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n211_), .A2(new_n255_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n256_), .B(new_n257_), .C1(new_n258_), .C2(KEYINPUT12), .ZN(new_n259_));
  AND2_X1   g058(.A1(G230gat), .A2(G233gat), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n256_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n260_), .B1(new_n262_), .B2(new_n258_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  XOR2_X1   g063(.A(KEYINPUT5), .B(G176gat), .Z(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT68), .B(G204gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G120gat), .B(G148gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n264_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n261_), .A2(new_n263_), .A3(new_n269_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n273_), .A2(KEYINPUT13), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT13), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n275_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G225gat), .A2(G233gat), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT87), .ZN(new_n279_));
  AND2_X1   g078(.A1(G155gat), .A2(G162gat), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT1), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n279_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n281_), .ZN(new_n283_));
  OR2_X1    g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n285_), .A2(KEYINPUT87), .A3(KEYINPUT1), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .A4(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G141gat), .A2(G148gat), .ZN(new_n288_));
  NOR2_X1   g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT86), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n287_), .A2(new_n288_), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT3), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n289_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT2), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n288_), .B(new_n294_), .ZN(new_n295_));
  OAI211_X1 g094(.A(new_n285_), .B(new_n284_), .C1(new_n293_), .C2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n291_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G127gat), .B(G134gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G113gat), .B(G120gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n297_), .A2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n291_), .A2(new_n296_), .A3(new_n300_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n302_), .A2(KEYINPUT4), .A3(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n300_), .B1(new_n291_), .B2(new_n296_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT4), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n278_), .B1(new_n304_), .B2(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(G57gat), .B(G85gat), .Z(new_n309_));
  XNOR2_X1  g108(.A(G1gat), .B(G29gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n278_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n315_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n316_));
  OR3_X1    g115(.A1(new_n308_), .A2(new_n314_), .A3(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n314_), .B1(new_n308_), .B2(new_n316_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT25), .B(G183gat), .ZN(new_n320_));
  INV_X1    g119(.A(G190gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT26), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT26), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(G190gat), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT92), .ZN(new_n325_));
  AND3_X1   g124(.A1(new_n322_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n325_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n320_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT23), .ZN(new_n329_));
  INV_X1    g128(.A(G183gat), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n329_), .B1(new_n330_), .B2(new_n321_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NOR3_X1   g132(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G169gat), .A2(G176gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n328_), .A2(new_n335_), .A3(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT22), .B(G169gat), .ZN(new_n341_));
  INV_X1    g140(.A(G176gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n338_), .B(KEYINPUT81), .ZN(new_n344_));
  NOR2_X1   g143(.A1(G183gat), .A2(G190gat), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n343_), .B(new_n344_), .C1(new_n333_), .C2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n340_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G197gat), .B(G204gat), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n348_), .A2(KEYINPUT89), .A3(KEYINPUT90), .A4(KEYINPUT21), .ZN(new_n349_));
  INV_X1    g148(.A(G204gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(G197gat), .ZN(new_n351_));
  INV_X1    g150(.A(G197gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(G204gat), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(new_n353_), .A3(KEYINPUT90), .ZN(new_n354_));
  NAND2_X1  g153(.A1(KEYINPUT89), .A2(KEYINPUT21), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G211gat), .B(G218gat), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n349_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(KEYINPUT89), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT21), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n359_), .B1(new_n360_), .B2(new_n348_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n358_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n347_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n344_), .A2(new_n337_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT26), .B(G190gat), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT80), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n367_), .B1(new_n330_), .B2(KEYINPUT25), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n330_), .A2(KEYINPUT25), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT25), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(KEYINPUT80), .A3(G183gat), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n366_), .A2(new_n368_), .A3(new_n369_), .A4(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n335_), .A2(new_n365_), .A3(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n362_), .A2(new_n346_), .A3(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n364_), .A2(KEYINPUT20), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G226gat), .A2(G233gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT19), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n362_), .A2(new_n340_), .A3(new_n346_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT20), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT98), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n379_), .A2(KEYINPUT98), .A3(KEYINPUT20), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n373_), .A2(new_n346_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n363_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n382_), .A2(new_n383_), .A3(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n378_), .B1(new_n386_), .B2(new_n377_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G8gat), .B(G36gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(G92gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT18), .B(G64gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT99), .B1(new_n387_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT99), .ZN(new_n394_));
  INV_X1    g193(.A(new_n377_), .ZN(new_n395_));
  AOI22_X1  g194(.A1(new_n380_), .A2(new_n381_), .B1(new_n384_), .B2(new_n363_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n395_), .B1(new_n396_), .B2(new_n383_), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n394_), .B(new_n391_), .C1(new_n397_), .C2(new_n378_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n375_), .A2(new_n377_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n385_), .A2(new_n379_), .A3(KEYINPUT20), .A4(new_n395_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n399_), .A2(new_n392_), .A3(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n393_), .A2(new_n398_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT27), .ZN(new_n403_));
  INV_X1    g202(.A(new_n401_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n392_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n405_));
  OR3_X1    g204(.A1(new_n404_), .A2(new_n405_), .A3(KEYINPUT27), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n319_), .B1(new_n403_), .B2(new_n406_), .ZN(new_n407_));
  XOR2_X1   g206(.A(new_n300_), .B(KEYINPUT31), .Z(new_n408_));
  XOR2_X1   g207(.A(G71gat), .B(G99gat), .Z(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT83), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G227gat), .A2(G233gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT82), .B(KEYINPUT30), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n373_), .A2(new_n346_), .A3(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n414_), .B1(new_n373_), .B2(new_n346_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G15gat), .B(G43gat), .ZN(new_n418_));
  NOR3_X1   g217(.A1(new_n416_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n418_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n414_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n384_), .A2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n420_), .B1(new_n422_), .B2(new_n415_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n413_), .B1(new_n419_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT84), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n418_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n422_), .A2(new_n415_), .A3(new_n420_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n426_), .A2(new_n427_), .A3(new_n412_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n424_), .A2(new_n425_), .A3(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n408_), .B1(new_n429_), .B2(KEYINPUT85), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT84), .B1(new_n408_), .B2(KEYINPUT85), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n431_), .B1(new_n424_), .B2(new_n428_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G22gat), .B(G50gat), .ZN(new_n434_));
  AND2_X1   g233(.A1(G228gat), .A2(G233gat), .ZN(new_n435_));
  OR3_X1    g234(.A1(new_n297_), .A2(KEYINPUT29), .A3(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n437_));
  OAI21_X1  g236(.A(new_n435_), .B1(new_n297_), .B2(KEYINPUT29), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n437_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n434_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n441_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n434_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(new_n439_), .A3(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n362_), .B1(new_n297_), .B2(KEYINPUT29), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G78gat), .B(G106gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT91), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n446_), .B(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n442_), .A2(new_n445_), .A3(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n449_), .B1(new_n442_), .B2(new_n445_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n433_), .A2(new_n450_), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n450_), .ZN(new_n454_));
  OAI22_X1  g253(.A1(new_n454_), .A2(new_n451_), .B1(new_n432_), .B2(new_n430_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n454_), .A2(new_n451_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n303_), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT94), .B1(new_n458_), .B2(new_n305_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT94), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n302_), .A2(new_n460_), .A3(new_n303_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n459_), .A2(new_n461_), .A3(new_n315_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(new_n313_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT95), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n304_), .A2(new_n278_), .A3(new_n307_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT96), .ZN(new_n467_));
  OR2_X1    g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n467_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n462_), .A2(KEYINPUT95), .A3(new_n313_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n465_), .A2(new_n468_), .A3(new_n469_), .A4(new_n470_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n404_), .A2(new_n405_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT33), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n318_), .A2(new_n473_), .ZN(new_n474_));
  OAI211_X1 g273(.A(KEYINPUT33), .B(new_n314_), .C1(new_n308_), .C2(new_n316_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n471_), .A2(new_n472_), .A3(new_n474_), .A4(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n386_), .A2(new_n377_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n399_), .A2(KEYINPUT97), .A3(new_n400_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n378_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n392_), .A2(KEYINPUT32), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .A4(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n399_), .A2(new_n400_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n480_), .B1(new_n483_), .B2(KEYINPUT97), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n482_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n319_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n433_), .B1(new_n476_), .B2(new_n486_), .ZN(new_n487_));
  AOI22_X1  g286(.A1(new_n407_), .A2(new_n456_), .B1(new_n457_), .B2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G15gat), .B(G22gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G1gat), .A2(G8gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT14), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G1gat), .B(G8gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G29gat), .B(G36gat), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G43gat), .B(G50gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n497_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(new_n495_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n494_), .B(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n494_), .A2(new_n501_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT15), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n501_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n498_), .A2(new_n500_), .A3(KEYINPUT15), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n503_), .B1(new_n494_), .B2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G229gat), .A2(G233gat), .ZN(new_n509_));
  MUX2_X1   g308(.A(new_n502_), .B(new_n508_), .S(new_n509_), .Z(new_n510_));
  XNOR2_X1  g309(.A(G113gat), .B(G141gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT78), .ZN(new_n512_));
  XOR2_X1   g311(.A(G169gat), .B(G197gat), .Z(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n510_), .B(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT79), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n277_), .A2(new_n488_), .A3(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n520_));
  AND2_X1   g319(.A1(G232gat), .A2(G233gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT35), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n235_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n249_), .A2(new_n228_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  AOI22_X1  g326(.A1(new_n527_), .A2(new_n237_), .B1(new_n241_), .B2(new_n244_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n253_), .B1(new_n528_), .B2(new_n227_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n507_), .B1(new_n529_), .B2(new_n226_), .ZN(new_n530_));
  OAI211_X1 g329(.A(new_n226_), .B(new_n501_), .C1(new_n246_), .C2(new_n254_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n524_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT71), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n498_), .A2(new_n500_), .A3(KEYINPUT15), .ZN(new_n535_));
  AOI21_X1  g334(.A(KEYINPUT15), .B1(new_n498_), .B2(new_n500_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n255_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(new_n531_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT71), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n539_), .A2(new_n540_), .A3(new_n524_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n522_), .A2(KEYINPUT35), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n538_), .A2(new_n542_), .A3(new_n531_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT70), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n538_), .A2(KEYINPUT70), .A3(new_n542_), .A4(new_n531_), .ZN(new_n546_));
  AOI22_X1  g345(.A1(new_n534_), .A2(new_n541_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G190gat), .B(G218gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G134gat), .B(G162gat), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n548_), .B(new_n549_), .Z(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT36), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  OR3_X1    g351(.A1(new_n547_), .A2(KEYINPUT72), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n550_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n554_), .A2(KEYINPUT36), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n547_), .A2(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT72), .B1(new_n547_), .B2(new_n552_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n553_), .A2(KEYINPUT37), .A3(new_n556_), .A4(new_n557_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n543_), .A2(new_n544_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n546_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n540_), .B1(new_n539_), .B2(new_n524_), .ZN(new_n561_));
  AOI211_X1 g360(.A(KEYINPUT71), .B(new_n523_), .C1(new_n538_), .C2(new_n531_), .ZN(new_n562_));
  OAI22_X1  g361(.A1(new_n559_), .A2(new_n560_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT73), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n534_), .A2(new_n541_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT73), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n545_), .A2(new_n546_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n565_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n564_), .A2(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(KEYINPUT74), .B1(new_n569_), .B2(new_n551_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT74), .ZN(new_n571_));
  AOI211_X1 g370(.A(new_n571_), .B(new_n552_), .C1(new_n564_), .C2(new_n568_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n556_), .ZN(new_n573_));
  NOR3_X1   g372(.A1(new_n570_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n558_), .B1(new_n574_), .B2(KEYINPUT37), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n494_), .B(new_n576_), .Z(new_n577_));
  XNOR2_X1  g376(.A(new_n211_), .B(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(KEYINPUT75), .B(KEYINPUT16), .Z(new_n579_));
  XNOR2_X1  g378(.A(G127gat), .B(G155gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G183gat), .B(G211gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n583_), .B(KEYINPUT17), .Z(new_n584_));
  NAND2_X1  g383(.A1(new_n578_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n577_), .B(new_n210_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT76), .B(KEYINPUT17), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n583_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT77), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n586_), .A2(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n585_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n575_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n519_), .A2(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n319_), .B(KEYINPUT100), .Z(new_n595_));
  NOR3_X1   g394(.A1(new_n594_), .A2(G1gat), .A3(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n407_), .A2(new_n456_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n487_), .A2(new_n457_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  AOI221_X4 g400(.A(KEYINPUT73), .B1(new_n545_), .B2(new_n546_), .C1(new_n534_), .C2(new_n541_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n566_), .B1(new_n565_), .B2(new_n567_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n551_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(new_n571_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n569_), .A2(KEYINPUT74), .A3(new_n551_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n605_), .A2(new_n556_), .A3(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n601_), .A2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT102), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n274_), .A2(new_n276_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n609_), .A2(new_n591_), .A3(new_n515_), .A4(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n319_), .ZN(new_n612_));
  OAI21_X1  g411(.A(G1gat), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n598_), .A2(new_n613_), .ZN(G1324gat));
  NAND2_X1  g413(.A1(new_n403_), .A2(new_n406_), .ZN(new_n615_));
  OAI21_X1  g414(.A(G8gat), .B1(new_n611_), .B2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT39), .ZN(new_n617_));
  NOR3_X1   g416(.A1(new_n594_), .A2(G8gat), .A3(new_n615_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT103), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g420(.A(new_n433_), .ZN(new_n622_));
  OAI21_X1  g421(.A(G15gat), .B1(new_n611_), .B2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT41), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n594_), .A2(G15gat), .A3(new_n622_), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n624_), .A2(new_n625_), .ZN(G1326gat));
  OAI21_X1  g425(.A(G22gat), .B1(new_n611_), .B2(new_n457_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT42), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n457_), .A2(G22gat), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n628_), .B1(new_n594_), .B2(new_n629_), .ZN(G1327gat));
  NOR2_X1   g429(.A1(new_n607_), .A2(new_n591_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n519_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(G29gat), .B1(new_n633_), .B2(new_n319_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n515_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n277_), .A2(new_n591_), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT43), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n637_), .B1(new_n575_), .B2(new_n601_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n558_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT37), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n639_), .B1(new_n607_), .B2(new_n640_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n641_), .A2(new_n488_), .A3(KEYINPUT43), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n636_), .B1(new_n638_), .B2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(KEYINPUT104), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT44), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n575_), .A2(new_n637_), .A3(new_n601_), .ZN(new_n646_));
  OAI21_X1  g445(.A(KEYINPUT43), .B1(new_n641_), .B2(new_n488_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT104), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n648_), .A2(new_n649_), .A3(new_n636_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n644_), .A2(new_n645_), .A3(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n610_), .A2(new_n592_), .A3(new_n515_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n652_), .B1(new_n647_), .B2(new_n646_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(KEYINPUT44), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n651_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n595_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n634_), .B1(new_n657_), .B2(G29gat), .ZN(G1328gat));
  XOR2_X1   g457(.A(new_n615_), .B(KEYINPUT107), .Z(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n632_), .A2(G36gat), .A3(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT106), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n615_), .B1(new_n653_), .B2(KEYINPUT44), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n651_), .A2(KEYINPUT105), .A3(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT105), .B1(new_n651_), .B2(new_n665_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n664_), .B1(new_n668_), .B2(G36gat), .ZN(new_n669_));
  INV_X1    g468(.A(G36gat), .ZN(new_n670_));
  NOR4_X1   g469(.A1(new_n666_), .A2(new_n667_), .A3(KEYINPUT106), .A4(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n663_), .B1(new_n669_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT46), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  OAI211_X1 g473(.A(KEYINPUT46), .B(new_n663_), .C1(new_n669_), .C2(new_n671_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1329gat));
  NAND3_X1  g475(.A1(new_n655_), .A2(G43gat), .A3(new_n433_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n632_), .A2(new_n622_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n677_), .B1(G43gat), .B2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g479(.A(new_n457_), .ZN(new_n681_));
  AOI21_X1  g480(.A(G50gat), .B1(new_n633_), .B2(new_n681_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n655_), .A2(new_n681_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n682_), .B1(new_n683_), .B2(G50gat), .ZN(G1331gat));
  INV_X1    g483(.A(G57gat), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n610_), .A2(new_n488_), .A3(new_n515_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(new_n593_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n685_), .B1(new_n687_), .B2(new_n595_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT109), .Z(new_n689_));
  NOR2_X1   g488(.A1(new_n517_), .A2(new_n592_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n609_), .A2(new_n277_), .A3(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(KEYINPUT110), .B(G57gat), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n691_), .A2(new_n612_), .A3(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n689_), .A2(new_n693_), .ZN(G1332gat));
  OAI21_X1  g493(.A(G64gat), .B1(new_n691_), .B2(new_n660_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT48), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n660_), .A2(G64gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n696_), .B1(new_n687_), .B2(new_n697_), .ZN(G1333gat));
  OAI21_X1  g497(.A(G71gat), .B1(new_n691_), .B2(new_n622_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT49), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n622_), .A2(G71gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n700_), .B1(new_n687_), .B2(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT111), .ZN(G1334gat));
  OAI21_X1  g502(.A(G78gat), .B1(new_n691_), .B2(new_n457_), .ZN(new_n704_));
  XOR2_X1   g503(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n457_), .A2(G78gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n706_), .B1(new_n687_), .B2(new_n707_), .ZN(G1335gat));
  NAND2_X1  g507(.A1(new_n686_), .A2(new_n631_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(G85gat), .B1(new_n710_), .B2(new_n656_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n610_), .A2(new_n515_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n648_), .A2(new_n592_), .A3(new_n712_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n713_), .A2(new_n222_), .A3(new_n612_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n711_), .A2(new_n714_), .ZN(G1336gat));
  OAI21_X1  g514(.A(new_n215_), .B1(new_n709_), .B2(new_n615_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n215_), .A2(KEYINPUT64), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n659_), .B1(new_n217_), .B2(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n716_), .B1(new_n713_), .B2(new_n718_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT113), .Z(G1337gat));
  INV_X1    g519(.A(new_n713_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n248_), .B1(new_n721_), .B2(new_n433_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n433_), .A2(new_n212_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n710_), .B2(new_n723_), .ZN(new_n724_));
  XOR2_X1   g523(.A(KEYINPUT114), .B(KEYINPUT51), .Z(new_n725_));
  XNOR2_X1  g524(.A(new_n724_), .B(new_n725_), .ZN(G1338gat));
  NAND2_X1  g525(.A1(KEYINPUT115), .A2(KEYINPUT52), .ZN(new_n727_));
  OAI211_X1 g526(.A(G106gat), .B(new_n727_), .C1(new_n713_), .C2(new_n457_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(KEYINPUT115), .A2(KEYINPUT52), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n728_), .B(new_n729_), .Z(new_n730_));
  NAND3_X1  g529(.A1(new_n710_), .A2(new_n213_), .A3(new_n681_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g532(.A(KEYINPUT55), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n734_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n259_), .A2(new_n260_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n259_), .A2(new_n734_), .A3(new_n260_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n270_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT118), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT56), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n743_), .A2(new_n635_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n272_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n502_), .A2(new_n509_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n508_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n514_), .B(new_n748_), .C1(new_n749_), .C2(new_n509_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n750_), .B1(new_n510_), .B2(new_n514_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n752_));
  OAI211_X1 g551(.A(KEYINPUT57), .B(new_n607_), .C1(new_n747_), .C2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT57), .ZN(new_n754_));
  INV_X1    g553(.A(new_n751_), .ZN(new_n755_));
  AOI22_X1  g554(.A1(new_n744_), .A2(new_n746_), .B1(new_n273_), .B2(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n754_), .B1(new_n756_), .B2(new_n574_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n739_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n272_), .B1(new_n758_), .B2(new_n742_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT58), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n755_), .B1(new_n739_), .B2(KEYINPUT56), .ZN(new_n761_));
  OR3_X1    g560(.A1(new_n759_), .A2(new_n760_), .A3(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n760_), .B1(new_n759_), .B2(new_n761_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n762_), .A2(new_n575_), .A3(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n753_), .A2(new_n757_), .A3(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT116), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n690_), .A2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(KEYINPUT116), .B1(new_n517_), .B2(new_n592_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n641_), .A2(new_n610_), .A3(new_n767_), .A4(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT117), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n770_), .A2(KEYINPUT54), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n769_), .B(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(KEYINPUT54), .ZN(new_n773_));
  AOI22_X1  g572(.A1(new_n765_), .A2(new_n592_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n656_), .A2(new_n433_), .A3(new_n615_), .A4(new_n457_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT119), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n774_), .A2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(G113gat), .B1(new_n777_), .B2(new_n515_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT59), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n779_), .B1(new_n776_), .B2(KEYINPUT121), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n776_), .A2(KEYINPUT121), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n774_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT120), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(new_n777_), .B2(new_n779_), .ZN(new_n784_));
  OAI211_X1 g583(.A(KEYINPUT120), .B(KEYINPUT59), .C1(new_n774_), .C2(new_n776_), .ZN(new_n785_));
  AOI211_X1 g584(.A(new_n518_), .B(new_n782_), .C1(new_n784_), .C2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n778_), .B1(new_n786_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g586(.A(G120gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n788_), .B1(new_n610_), .B2(KEYINPUT60), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT122), .B1(new_n788_), .B2(KEYINPUT60), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT122), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n777_), .B(new_n791_), .C1(new_n792_), .C2(new_n789_), .ZN(new_n793_));
  AOI211_X1 g592(.A(new_n610_), .B(new_n782_), .C1(new_n784_), .C2(new_n785_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n793_), .B1(new_n794_), .B2(new_n788_), .ZN(G1341gat));
  AOI21_X1  g594(.A(G127gat), .B1(new_n777_), .B2(new_n591_), .ZN(new_n796_));
  INV_X1    g595(.A(G127gat), .ZN(new_n797_));
  AOI211_X1 g596(.A(new_n797_), .B(new_n782_), .C1(new_n784_), .C2(new_n785_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n796_), .B1(new_n798_), .B2(new_n591_), .ZN(G1342gat));
  AOI21_X1  g598(.A(G134gat), .B1(new_n777_), .B2(new_n574_), .ZN(new_n800_));
  AOI211_X1 g599(.A(new_n641_), .B(new_n782_), .C1(new_n784_), .C2(new_n785_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n801_), .B2(G134gat), .ZN(G1343gat));
  NOR3_X1   g601(.A1(new_n774_), .A2(new_n455_), .A3(new_n595_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n803_), .A2(new_n515_), .A3(new_n660_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g604(.A1(new_n803_), .A2(new_n277_), .A3(new_n660_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g606(.A1(new_n803_), .A2(new_n591_), .A3(new_n660_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(KEYINPUT61), .B(G155gat), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n808_), .B(new_n809_), .ZN(G1346gat));
  AND4_X1   g609(.A1(G162gat), .A2(new_n803_), .A3(new_n575_), .A4(new_n660_), .ZN(new_n811_));
  INV_X1    g610(.A(G162gat), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n803_), .A2(new_n574_), .A3(new_n660_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n811_), .B1(new_n812_), .B2(new_n813_), .ZN(G1347gat));
  NAND2_X1  g613(.A1(new_n765_), .A2(new_n592_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n772_), .A2(new_n773_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n660_), .A2(new_n453_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n595_), .A3(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(G169gat), .B1(new_n819_), .B2(new_n635_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT62), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n819_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n823_), .A2(new_n341_), .A3(new_n515_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n820_), .A2(new_n821_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n822_), .A2(new_n824_), .A3(new_n825_), .ZN(G1348gat));
  NOR2_X1   g625(.A1(new_n819_), .A2(new_n610_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(new_n342_), .ZN(G1349gat));
  OAI21_X1  g627(.A(new_n320_), .B1(KEYINPUT123), .B2(G183gat), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n823_), .A2(new_n591_), .A3(new_n829_), .ZN(new_n830_));
  OAI211_X1 g629(.A(KEYINPUT123), .B(new_n330_), .C1(new_n819_), .C2(new_n592_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT124), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT124), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n830_), .A2(new_n831_), .A3(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(G1350gat));
  OAI21_X1  g635(.A(G190gat), .B1(new_n819_), .B2(new_n641_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n823_), .B1(new_n327_), .B2(new_n326_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(new_n838_), .B2(new_n607_), .ZN(G1351gat));
  NOR2_X1   g638(.A1(new_n774_), .A2(new_n319_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n455_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n840_), .A2(new_n841_), .A3(new_n515_), .A4(new_n659_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n352_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(KEYINPUT126), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT126), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n842_), .A2(new_n845_), .A3(new_n352_), .ZN(new_n846_));
  OAI21_X1  g645(.A(KEYINPUT125), .B1(new_n842_), .B2(new_n352_), .ZN(new_n847_));
  NOR4_X1   g646(.A1(new_n774_), .A2(new_n319_), .A3(new_n455_), .A4(new_n660_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT125), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n848_), .A2(new_n849_), .A3(G197gat), .A4(new_n515_), .ZN(new_n850_));
  AOI22_X1  g649(.A1(new_n844_), .A2(new_n846_), .B1(new_n847_), .B2(new_n850_), .ZN(G1352gat));
  NAND2_X1  g650(.A1(new_n848_), .A2(new_n277_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n853_));
  XOR2_X1   g652(.A(new_n852_), .B(new_n853_), .Z(G1353gat));
  AOI211_X1 g653(.A(KEYINPUT63), .B(G211gat), .C1(new_n848_), .C2(new_n591_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n840_), .A2(new_n841_), .A3(new_n659_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n856_), .A2(new_n592_), .ZN(new_n857_));
  XOR2_X1   g656(.A(KEYINPUT63), .B(G211gat), .Z(new_n858_));
  AOI21_X1  g657(.A(new_n855_), .B1(new_n857_), .B2(new_n858_), .ZN(G1354gat));
  AOI21_X1  g658(.A(G218gat), .B1(new_n848_), .B2(new_n574_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n856_), .A2(new_n641_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(G218gat), .B2(new_n861_), .ZN(G1355gat));
endmodule


