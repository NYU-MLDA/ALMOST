//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 1 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 0 1 0 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n669_, new_n670_, new_n671_, new_n672_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n799_, new_n800_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n807_, new_n808_, new_n809_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n816_, new_n817_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n848_, new_n849_, new_n850_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_;
  INV_X1    g000(.A(KEYINPUT99), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT26), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(G190gat), .ZN(new_n204_));
  OR2_X1    g003(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n205_));
  NAND2_X1  g004(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G183gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT83), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n204_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G183gat), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n211_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n212_));
  AOI22_X1  g011(.A1(new_n212_), .A2(KEYINPUT83), .B1(KEYINPUT25), .B2(new_n211_), .ZN(new_n213_));
  INV_X1    g012(.A(G190gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n214_), .A2(KEYINPUT26), .ZN(new_n215_));
  XOR2_X1   g014(.A(new_n215_), .B(KEYINPUT84), .Z(new_n216_));
  NAND3_X1  g015(.A1(new_n210_), .A2(new_n213_), .A3(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218_));
  XOR2_X1   g017(.A(new_n218_), .B(KEYINPUT23), .Z(new_n219_));
  OR2_X1    g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n220_), .A2(KEYINPUT24), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n220_), .A2(KEYINPUT24), .A3(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT85), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n217_), .A2(new_n222_), .A3(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(KEYINPUT22), .B(G169gat), .Z(new_n227_));
  NOR2_X1   g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228_));
  OAI221_X1 g027(.A(new_n223_), .B1(G176gat), .B2(new_n227_), .C1(new_n219_), .C2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n226_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT30), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G127gat), .B(G134gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G113gat), .B(G120gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n231_), .B(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G227gat), .A2(G233gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT31), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n236_), .B(new_n238_), .ZN(new_n239_));
  XOR2_X1   g038(.A(G15gat), .B(G43gat), .Z(new_n240_));
  XOR2_X1   g039(.A(G71gat), .B(G99gat), .Z(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  XOR2_X1   g041(.A(new_n239_), .B(new_n242_), .Z(new_n243_));
  AOI21_X1  g042(.A(KEYINPUT87), .B1(G141gat), .B2(G148gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT2), .ZN(new_n245_));
  INV_X1    g044(.A(G141gat), .ZN(new_n246_));
  INV_X1    g045(.A(G148gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT86), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n248_), .B1(new_n249_), .B2(KEYINPUT3), .ZN(new_n250_));
  OR3_X1    g049(.A1(new_n248_), .A2(new_n249_), .A3(KEYINPUT3), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n245_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G155gat), .A2(G162gat), .ZN(new_n253_));
  OR2_X1    g052(.A1(G155gat), .A2(G162gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT88), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT88), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n252_), .A2(new_n257_), .A3(new_n253_), .A4(new_n254_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n253_), .A2(KEYINPUT1), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n253_), .A2(KEYINPUT1), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(new_n254_), .A3(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G141gat), .A2(G148gat), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n262_), .A2(new_n263_), .A3(new_n248_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n259_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(new_n235_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n264_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n267_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(new_n234_), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n266_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G225gat), .A2(G233gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT94), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n266_), .A2(new_n269_), .A3(KEYINPUT4), .ZN(new_n275_));
  OR3_X1    g074(.A1(new_n268_), .A2(KEYINPUT4), .A3(new_n234_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(new_n276_), .A3(new_n272_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n274_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G1gat), .B(G29gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(G85gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT0), .B(G57gat), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n280_), .B(new_n281_), .Z(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n278_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT97), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n274_), .A2(new_n277_), .A3(new_n282_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT97), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n278_), .A2(new_n287_), .A3(new_n283_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n285_), .A2(new_n286_), .A3(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n243_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT90), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G22gat), .B(G50gat), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT29), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n268_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT28), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n295_), .A2(KEYINPUT28), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n293_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n298_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n300_), .A2(new_n296_), .A3(new_n292_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n291_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G211gat), .B(G218gat), .ZN(new_n303_));
  INV_X1    g102(.A(G197gat), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n304_), .A2(G204gat), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n303_), .B(KEYINPUT21), .C1(KEYINPUT89), .C2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G197gat), .B(G204gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n303_), .A2(KEYINPUT21), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n311_), .B1(new_n265_), .B2(KEYINPUT29), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G228gat), .A2(G233gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G78gat), .B(G106gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n302_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n299_), .A2(new_n301_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n314_), .A2(new_n315_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n319_), .B1(new_n320_), .B2(new_n302_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n316_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n317_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT20), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n204_), .A2(new_n215_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT91), .ZN(new_n326_));
  XOR2_X1   g125(.A(KEYINPUT25), .B(G183gat), .Z(new_n327_));
  OAI21_X1  g126(.A(new_n224_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT92), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT92), .ZN(new_n330_));
  OAI211_X1 g129(.A(new_n330_), .B(new_n224_), .C1(new_n326_), .C2(new_n327_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n329_), .A2(new_n222_), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(new_n229_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n324_), .B1(new_n333_), .B2(new_n310_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n311_), .A2(new_n229_), .A3(new_n226_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G226gat), .A2(G233gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT19), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G8gat), .B(G36gat), .ZN(new_n340_));
  INV_X1    g139(.A(G92gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT18), .B(G64gat), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n342_), .B(new_n343_), .Z(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n333_), .A2(new_n310_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n324_), .B1(new_n230_), .B2(new_n310_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n338_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n346_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n339_), .A2(new_n345_), .A3(new_n351_), .ZN(new_n352_));
  AND3_X1   g151(.A1(new_n334_), .A2(new_n348_), .A3(new_n335_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT96), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n311_), .B1(new_n333_), .B2(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(KEYINPUT96), .B1(new_n332_), .B2(new_n229_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n347_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n353_), .B1(new_n338_), .B2(new_n357_), .ZN(new_n358_));
  OAI211_X1 g157(.A(KEYINPUT27), .B(new_n352_), .C1(new_n358_), .C2(new_n345_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT27), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n345_), .B1(new_n339_), .B2(new_n351_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n348_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n362_), .A2(new_n344_), .A3(new_n350_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n360_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n359_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n290_), .A2(new_n323_), .A3(new_n366_), .ZN(new_n367_));
  NOR3_X1   g166(.A1(new_n323_), .A2(new_n365_), .A3(new_n289_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT98), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n287_), .B1(new_n278_), .B2(new_n283_), .ZN(new_n370_));
  AOI211_X1 g169(.A(KEYINPUT97), .B(new_n282_), .C1(new_n274_), .C2(new_n277_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n286_), .ZN(new_n372_));
  NOR3_X1   g171(.A1(new_n370_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n345_), .A2(KEYINPUT32), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT95), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n339_), .A2(new_n351_), .A3(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n376_), .B1(new_n358_), .B2(new_n374_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n369_), .B1(new_n373_), .B2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n270_), .A2(new_n272_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n275_), .A2(new_n273_), .A3(new_n276_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(new_n380_), .A3(new_n283_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n286_), .B(KEYINPUT33), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n344_), .B1(new_n362_), .B2(new_n350_), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n352_), .A2(KEYINPUT93), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(KEYINPUT93), .B1(new_n352_), .B2(new_n383_), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n381_), .B(new_n382_), .C1(new_n384_), .C2(new_n385_), .ZN(new_n386_));
  OR2_X1    g185(.A1(new_n358_), .A2(new_n374_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n289_), .A2(new_n387_), .A3(KEYINPUT98), .A4(new_n376_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n378_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n368_), .B1(new_n389_), .B2(new_n323_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n243_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n367_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(G85gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(new_n341_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G85gat), .A2(G92gat), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT7), .ZN(new_n397_));
  INV_X1    g196(.A(G99gat), .ZN(new_n398_));
  INV_X1    g197(.A(G106gat), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .A4(KEYINPUT67), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT67), .ZN(new_n401_));
  OAI22_X1  g200(.A1(new_n401_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(KEYINPUT7), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n400_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT6), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n405_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n396_), .B1(new_n404_), .B2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT68), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT68), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n411_), .B(new_n396_), .C1(new_n404_), .C2(new_n408_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n410_), .A2(KEYINPUT8), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT9), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n414_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n415_));
  AOI21_X1  g214(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n416_));
  OR3_X1    g215(.A1(new_n415_), .A2(KEYINPUT66), .A3(new_n416_), .ZN(new_n417_));
  XOR2_X1   g216(.A(KEYINPUT10), .B(G99gat), .Z(new_n418_));
  NAND3_X1  g217(.A1(new_n418_), .A2(KEYINPUT65), .A3(new_n399_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT65), .ZN(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT10), .B(G99gat), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n420_), .B1(new_n421_), .B2(G106gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n419_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n408_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT66), .B1(new_n415_), .B2(new_n416_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n417_), .A2(new_n423_), .A3(new_n424_), .A4(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT8), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n409_), .A2(KEYINPUT68), .A3(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n413_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G71gat), .B(G78gat), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G57gat), .B(G64gat), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n431_), .B1(KEYINPUT11), .B2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(KEYINPUT11), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n433_), .B1(new_n434_), .B2(new_n431_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n429_), .A2(new_n436_), .ZN(new_n437_));
  XOR2_X1   g236(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G230gat), .A2(G233gat), .ZN(new_n440_));
  XOR2_X1   g239(.A(new_n440_), .B(KEYINPUT64), .Z(new_n441_));
  AND3_X1   g240(.A1(new_n413_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(new_n435_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n429_), .A2(KEYINPUT12), .A3(new_n436_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n439_), .A2(new_n441_), .A3(new_n443_), .A4(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT70), .ZN(new_n446_));
  AND4_X1   g245(.A1(new_n426_), .A2(new_n413_), .A3(new_n428_), .A4(new_n435_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n447_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT70), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n448_), .A2(new_n449_), .A3(new_n441_), .A4(new_n444_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n446_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n443_), .A2(new_n437_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n441_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n451_), .A2(new_n454_), .ZN(new_n455_));
  XOR2_X1   g254(.A(G176gat), .B(G204gat), .Z(new_n456_));
  XNOR2_X1  g255(.A(G120gat), .B(G148gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n455_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n460_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n451_), .A2(new_n454_), .A3(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT13), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n461_), .A2(KEYINPUT13), .A3(new_n463_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G1gat), .B(G8gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT75), .ZN(new_n470_));
  INV_X1    g269(.A(G15gat), .ZN(new_n471_));
  INV_X1    g270(.A(G22gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G15gat), .A2(G22gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G1gat), .A2(G8gat), .ZN(new_n475_));
  AOI22_X1  g274(.A1(new_n473_), .A2(new_n474_), .B1(KEYINPUT14), .B2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n470_), .B(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT72), .B(G43gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G29gat), .B(G36gat), .ZN(new_n479_));
  INV_X1    g278(.A(G50gat), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n480_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n478_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n481_), .A2(new_n482_), .A3(new_n478_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT15), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n485_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT15), .ZN(new_n488_));
  NOR3_X1   g287(.A1(new_n487_), .A2(new_n488_), .A3(new_n483_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n477_), .B1(new_n486_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G229gat), .A2(G233gat), .ZN(new_n491_));
  XOR2_X1   g290(.A(new_n470_), .B(new_n476_), .Z(new_n492_));
  NOR2_X1   g291(.A1(new_n487_), .A2(new_n483_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n490_), .A2(new_n491_), .A3(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT79), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n492_), .B(new_n493_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n491_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT79), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n490_), .A2(new_n500_), .A3(new_n491_), .A4(new_n494_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n496_), .A2(new_n499_), .A3(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(KEYINPUT80), .B(G113gat), .Z(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT81), .B(G141gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G169gat), .B(G197gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n502_), .A2(new_n508_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n496_), .A2(new_n499_), .A3(new_n501_), .A4(new_n507_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n468_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n392_), .A2(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n429_), .B1(new_n489_), .B2(new_n486_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT73), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G232gat), .A2(G233gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT34), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n517_), .A2(KEYINPUT35), .A3(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n442_), .A2(new_n493_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(new_n515_), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n519_), .A2(KEYINPUT35), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n520_), .A2(new_n522_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G190gat), .B(G218gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G134gat), .B(G162gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n527_), .B(new_n528_), .Z(new_n529_));
  INV_X1    g328(.A(KEYINPUT36), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n526_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n526_), .A2(new_n530_), .A3(new_n529_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(KEYINPUT74), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n535_), .A3(KEYINPUT37), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT37), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n532_), .B(new_n533_), .C1(KEYINPUT74), .C2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT78), .ZN(new_n540_));
  XOR2_X1   g339(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n541_));
  XNOR2_X1  g340(.A(G127gat), .B(G155gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G183gat), .B(G211gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n546_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G231gat), .A2(G233gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n477_), .B(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n435_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n551_), .A2(new_n435_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n549_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  OR2_X1    g354(.A1(new_n551_), .A2(new_n435_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n556_), .A2(new_n547_), .A3(new_n552_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT77), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n555_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n558_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n540_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n556_), .A2(new_n547_), .A3(new_n552_), .ZN(new_n562_));
  AOI22_X1  g361(.A1(new_n556_), .A2(new_n552_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT77), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n555_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n564_), .A2(KEYINPUT78), .A3(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n561_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n539_), .A2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n202_), .B1(new_n514_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(G1gat), .ZN(new_n570_));
  INV_X1    g369(.A(new_n568_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n392_), .A2(KEYINPUT99), .A3(new_n513_), .A4(new_n571_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n569_), .A2(new_n570_), .A3(new_n289_), .A4(new_n572_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n573_), .A2(KEYINPUT100), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(KEYINPUT100), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT38), .ZN(new_n576_));
  OR3_X1    g375(.A1(new_n574_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n559_), .A2(new_n560_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n392_), .A2(new_n534_), .A3(new_n513_), .A4(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(G1gat), .B1(new_n579_), .B2(new_n373_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n576_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n577_), .A2(new_n580_), .A3(new_n581_), .ZN(G1324gat));
  XNOR2_X1  g381(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(G8gat), .B1(new_n579_), .B2(new_n366_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT102), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(KEYINPUT39), .B1(new_n585_), .B2(KEYINPUT102), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(G8gat), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n569_), .A2(new_n590_), .A3(new_n365_), .A4(new_n572_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT101), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n584_), .B1(new_n589_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n592_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n588_), .B(new_n586_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n594_), .A2(new_n595_), .A3(new_n583_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n593_), .A2(new_n596_), .ZN(G1325gat));
  AND2_X1   g396(.A1(new_n569_), .A2(new_n572_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n598_), .A2(new_n471_), .A3(new_n391_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT104), .Z(new_n600_));
  OAI21_X1  g399(.A(G15gat), .B1(new_n579_), .B2(new_n243_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT41), .Z(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(G1326gat));
  OAI21_X1  g402(.A(G22gat), .B1(new_n579_), .B2(new_n323_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT42), .ZN(new_n605_));
  INV_X1    g404(.A(new_n323_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n598_), .A2(new_n472_), .A3(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(G1327gat));
  INV_X1    g407(.A(new_n567_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT43), .ZN(new_n610_));
  INV_X1    g409(.A(new_n539_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n392_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n610_), .B1(new_n392_), .B2(new_n611_), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n513_), .B(new_n609_), .C1(new_n612_), .C2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT44), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n392_), .A2(new_n611_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(KEYINPUT43), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n392_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n620_), .A2(KEYINPUT44), .A3(new_n513_), .A4(new_n609_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n616_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(new_n289_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(G29gat), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT105), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n534_), .A2(new_n567_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n625_), .B1(new_n514_), .B2(new_n627_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n392_), .A2(KEYINPUT105), .A3(new_n513_), .A4(new_n626_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n373_), .A2(G29gat), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT106), .Z(new_n632_));
  OAI21_X1  g431(.A(new_n624_), .B1(new_n630_), .B2(new_n632_), .ZN(G1328gat));
  NAND3_X1  g432(.A1(new_n616_), .A2(new_n621_), .A3(new_n365_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(G36gat), .ZN(new_n635_));
  INV_X1    g434(.A(G36gat), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n365_), .B(KEYINPUT107), .Z(new_n637_));
  NAND4_X1  g436(.A1(new_n628_), .A2(new_n636_), .A3(new_n629_), .A4(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT45), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n635_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT46), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n635_), .A2(KEYINPUT46), .A3(new_n639_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(G1329gat));
  NAND4_X1  g443(.A1(new_n616_), .A2(new_n621_), .A3(G43gat), .A4(new_n391_), .ZN(new_n645_));
  INV_X1    g444(.A(G43gat), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n646_), .B1(new_n630_), .B2(new_n243_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(G1330gat));
  NAND3_X1  g449(.A1(new_n622_), .A2(G50gat), .A3(new_n606_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n480_), .B1(new_n630_), .B2(new_n323_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(G1331gat));
  INV_X1    g452(.A(new_n468_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n654_), .A2(new_n511_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n392_), .A2(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n656_), .A2(new_n568_), .ZN(new_n657_));
  AOI21_X1  g456(.A(G57gat), .B1(new_n657_), .B2(new_n289_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT109), .ZN(new_n659_));
  INV_X1    g458(.A(new_n534_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n656_), .A2(new_n660_), .A3(new_n609_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n289_), .A2(G57gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n659_), .B1(new_n661_), .B2(new_n662_), .ZN(G1332gat));
  INV_X1    g462(.A(G64gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n664_), .B1(new_n661_), .B2(new_n637_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT48), .Z(new_n666_));
  NAND3_X1  g465(.A1(new_n657_), .A2(new_n664_), .A3(new_n637_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1333gat));
  INV_X1    g467(.A(G71gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n669_), .B1(new_n661_), .B2(new_n391_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT49), .Z(new_n671_));
  NAND3_X1  g470(.A1(new_n657_), .A2(new_n669_), .A3(new_n391_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1334gat));
  INV_X1    g472(.A(G78gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n661_), .B2(new_n606_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT50), .Z(new_n676_));
  NOR2_X1   g475(.A1(new_n323_), .A2(G78gat), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT110), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n657_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n676_), .A2(new_n679_), .ZN(G1335gat));
  OAI211_X1 g479(.A(new_n609_), .B(new_n655_), .C1(new_n612_), .C2(new_n613_), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT111), .Z(new_n682_));
  OAI21_X1  g481(.A(G85gat), .B1(new_n682_), .B2(new_n373_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n656_), .A2(new_n627_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(new_n393_), .A3(new_n289_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(G1336gat));
  INV_X1    g485(.A(new_n637_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G92gat), .B1(new_n682_), .B2(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n684_), .A2(new_n341_), .A3(new_n365_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1337gat));
  OAI21_X1  g489(.A(G99gat), .B1(new_n681_), .B2(new_n243_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n684_), .A2(new_n418_), .A3(new_n391_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT112), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT51), .ZN(new_n694_));
  AOI22_X1  g493(.A1(new_n691_), .A2(new_n692_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n693_), .A2(new_n694_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n695_), .B(new_n696_), .ZN(G1338gat));
  OAI21_X1  g496(.A(G106gat), .B1(new_n681_), .B2(new_n323_), .ZN(new_n698_));
  XOR2_X1   g497(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n684_), .A2(new_n399_), .A3(new_n606_), .ZN(new_n702_));
  OAI211_X1 g501(.A(G106gat), .B(new_n699_), .C1(new_n681_), .C2(new_n323_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n701_), .A2(new_n702_), .A3(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g504(.A1(new_n466_), .A2(new_n567_), .A3(new_n512_), .A4(new_n467_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT114), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n706_), .B(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT54), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n708_), .A2(new_n709_), .A3(new_n539_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n708_), .B2(new_n539_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT57), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT115), .ZN(new_n714_));
  AOI21_X1  g513(.A(KEYINPUT55), .B1(new_n446_), .B2(new_n450_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n448_), .A2(new_n444_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(new_n453_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n448_), .A2(KEYINPUT55), .A3(new_n441_), .A4(new_n444_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n460_), .B1(new_n715_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT56), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  OAI211_X1 g521(.A(KEYINPUT56), .B(new_n460_), .C1(new_n715_), .C2(new_n719_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n463_), .A2(new_n511_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n714_), .B1(new_n724_), .B2(new_n726_), .ZN(new_n727_));
  AOI211_X1 g526(.A(KEYINPUT115), .B(new_n725_), .C1(new_n722_), .C2(new_n723_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n497_), .A2(new_n491_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n490_), .A2(new_n498_), .A3(new_n494_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n729_), .A2(new_n508_), .A3(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n464_), .A2(new_n510_), .A3(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n727_), .A2(new_n728_), .A3(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n713_), .B1(new_n734_), .B2(new_n660_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT116), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n724_), .A2(new_n726_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT115), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n724_), .A2(new_n714_), .A3(new_n726_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(new_n732_), .A3(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n741_), .A2(KEYINPUT57), .A3(new_n534_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT117), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n722_), .A2(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n720_), .A2(KEYINPUT117), .A3(new_n721_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n744_), .A2(new_n723_), .A3(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n463_), .A2(new_n510_), .A3(new_n731_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT58), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n746_), .A2(KEYINPUT58), .A3(new_n748_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(new_n611_), .A3(new_n752_), .ZN(new_n753_));
  OAI211_X1 g552(.A(KEYINPUT116), .B(new_n713_), .C1(new_n734_), .C2(new_n660_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n737_), .A2(new_n742_), .A3(new_n753_), .A4(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n578_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n712_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  NOR4_X1   g556(.A1(new_n243_), .A2(new_n606_), .A3(new_n373_), .A4(new_n365_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(KEYINPUT118), .B1(new_n757_), .B2(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n754_), .A2(new_n742_), .A3(new_n753_), .ZN(new_n761_));
  AOI21_X1  g560(.A(KEYINPUT57), .B1(new_n741_), .B2(new_n534_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n762_), .A2(KEYINPUT116), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n756_), .B1(new_n761_), .B2(new_n763_), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n710_), .A2(new_n711_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT118), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n766_), .A2(new_n767_), .A3(new_n758_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n760_), .A2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(G113gat), .B1(new_n769_), .B2(new_n511_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n766_), .A2(new_n758_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n753_), .A2(new_n742_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n609_), .B1(new_n772_), .B2(new_n762_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT120), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT120), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n775_), .B(new_n609_), .C1(new_n772_), .C2(new_n762_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n774_), .A2(new_n765_), .A3(new_n776_), .ZN(new_n777_));
  XOR2_X1   g576(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n778_));
  NOR2_X1   g577(.A1(new_n759_), .A2(new_n778_), .ZN(new_n779_));
  AOI22_X1  g578(.A1(new_n771_), .A2(KEYINPUT59), .B1(new_n777_), .B2(new_n779_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n780_), .A2(new_n511_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n770_), .B1(new_n781_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g581(.A(G120gat), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(new_n780_), .B2(new_n468_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(KEYINPUT60), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n783_), .B1(new_n654_), .B2(KEYINPUT60), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  AOI211_X1 g586(.A(new_n785_), .B(new_n787_), .C1(new_n760_), .C2(new_n768_), .ZN(new_n788_));
  OAI21_X1  g587(.A(KEYINPUT121), .B1(new_n784_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n777_), .A2(new_n779_), .ZN(new_n790_));
  OAI21_X1  g589(.A(KEYINPUT59), .B1(new_n757_), .B2(new_n759_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(new_n791_), .A3(new_n468_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(G120gat), .ZN(new_n793_));
  INV_X1    g592(.A(new_n785_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n769_), .A2(new_n794_), .A3(new_n786_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT121), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n793_), .A2(new_n795_), .A3(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n789_), .A2(new_n797_), .ZN(G1341gat));
  AOI21_X1  g597(.A(G127gat), .B1(new_n769_), .B2(new_n567_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n578_), .A2(G127gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n780_), .B2(new_n800_), .ZN(G1342gat));
  AOI21_X1  g600(.A(G134gat), .B1(new_n769_), .B2(new_n660_), .ZN(new_n802_));
  XOR2_X1   g601(.A(KEYINPUT122), .B(G134gat), .Z(new_n803_));
  NAND2_X1  g602(.A1(new_n611_), .A2(new_n803_), .ZN(new_n804_));
  XOR2_X1   g603(.A(new_n804_), .B(KEYINPUT123), .Z(new_n805_));
  AOI21_X1  g604(.A(new_n802_), .B1(new_n780_), .B2(new_n805_), .ZN(G1343gat));
  NOR3_X1   g605(.A1(new_n757_), .A2(new_n323_), .A3(new_n391_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n637_), .A2(new_n373_), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n807_), .A2(new_n511_), .A3(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(new_n246_), .ZN(G1344gat));
  AND2_X1   g609(.A1(new_n807_), .A2(new_n808_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n468_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(G148gat), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n811_), .A2(new_n247_), .A3(new_n468_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(G1345gat));
  NAND3_X1  g614(.A1(new_n807_), .A2(new_n567_), .A3(new_n808_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(KEYINPUT61), .B(G155gat), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n816_), .B(new_n817_), .ZN(G1346gat));
  NAND4_X1  g617(.A1(new_n807_), .A2(G162gat), .A3(new_n611_), .A4(new_n808_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n391_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n820_), .A2(new_n660_), .A3(new_n606_), .A4(new_n808_), .ZN(new_n821_));
  INV_X1    g620(.A(G162gat), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n819_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT124), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT124), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n819_), .A2(new_n823_), .A3(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(G1347gat));
  NAND3_X1  g627(.A1(new_n637_), .A2(new_n323_), .A3(new_n290_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n777_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n511_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(G169gat), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT62), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  OR2_X1    g634(.A1(new_n832_), .A2(new_n227_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n832_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n835_), .A2(new_n836_), .A3(new_n837_), .ZN(G1348gat));
  AOI21_X1  g637(.A(G176gat), .B1(new_n831_), .B2(new_n468_), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n766_), .A2(G176gat), .A3(new_n468_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n839_), .B1(new_n830_), .B2(new_n840_), .ZN(G1349gat));
  NAND3_X1  g640(.A1(new_n831_), .A2(new_n327_), .A3(new_n578_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n842_), .A2(KEYINPUT125), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n842_), .A2(KEYINPUT125), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n829_), .A2(new_n609_), .ZN(new_n845_));
  AOI21_X1  g644(.A(G183gat), .B1(new_n766_), .B2(new_n845_), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n843_), .A2(new_n844_), .A3(new_n846_), .ZN(G1350gat));
  INV_X1    g646(.A(new_n326_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n831_), .A2(new_n660_), .A3(new_n848_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n831_), .A2(new_n611_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(new_n214_), .ZN(G1351gat));
  NOR3_X1   g650(.A1(new_n687_), .A2(new_n289_), .A3(new_n323_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n820_), .A2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(KEYINPUT126), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT126), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n820_), .A2(new_n855_), .A3(new_n852_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n512_), .B1(new_n854_), .B2(new_n856_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(new_n304_), .ZN(G1352gat));
  NAND2_X1  g657(.A1(new_n854_), .A2(new_n856_), .ZN(new_n859_));
  AND3_X1   g658(.A1(new_n859_), .A2(G204gat), .A3(new_n468_), .ZN(new_n860_));
  AOI21_X1  g659(.A(G204gat), .B1(new_n859_), .B2(new_n468_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1353gat));
  NAND2_X1  g661(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n863_));
  AND4_X1   g662(.A1(new_n855_), .A2(new_n766_), .A3(new_n243_), .A4(new_n852_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n855_), .B1(new_n820_), .B2(new_n852_), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n578_), .B(new_n863_), .C1(new_n864_), .C2(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(KEYINPUT127), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n866_), .B(new_n868_), .ZN(G1354gat));
  NAND2_X1  g668(.A1(new_n859_), .A2(new_n660_), .ZN(new_n870_));
  INV_X1    g669(.A(G218gat), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n871_), .B1(new_n854_), .B2(new_n856_), .ZN(new_n872_));
  AOI22_X1  g671(.A1(new_n870_), .A2(new_n871_), .B1(new_n872_), .B2(new_n611_), .ZN(G1355gat));
endmodule


