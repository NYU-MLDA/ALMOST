//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 1 1 0 0 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0 1 1 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 1 1 1 1 1 1 0 1 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n677_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n813_, new_n815_, new_n816_, new_n818_,
    new_n819_, new_n820_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n838_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n847_, new_n848_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G230gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G57gat), .B(G64gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT11), .ZN(new_n205_));
  XOR2_X1   g004(.A(G71gat), .B(G78gat), .Z(new_n206_));
  OR2_X1    g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n204_), .A2(KEYINPUT11), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n205_), .A2(new_n206_), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n207_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G85gat), .ZN(new_n211_));
  INV_X1    g010(.A(G92gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT9), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G85gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n214_), .B1(new_n215_), .B2(new_n212_), .ZN(new_n216_));
  AND2_X1   g015(.A1(G85gat), .A2(G92gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT9), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  AND2_X1   g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT66), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n222_), .A2(KEYINPUT6), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT6), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n224_), .A2(KEYINPUT66), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n221_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(KEYINPUT66), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n222_), .A2(KEYINPUT6), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n228_), .A3(new_n220_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n226_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT10), .B(G99gat), .ZN(new_n231_));
  OR3_X1    g030(.A1(new_n231_), .A2(KEYINPUT64), .A3(G106gat), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT64), .B1(new_n231_), .B2(G106gat), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n219_), .A2(new_n230_), .A3(new_n232_), .A4(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT7), .ZN(new_n235_));
  INV_X1    g034(.A(G99gat), .ZN(new_n236_));
  INV_X1    g035(.A(G106gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n240_), .B1(new_n226_), .B2(new_n229_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n242_));
  NOR2_X1   g041(.A1(G85gat), .A2(G92gat), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n242_), .B1(new_n217_), .B2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G85gat), .A2(G92gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n213_), .A2(KEYINPUT67), .A3(new_n245_), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  NOR3_X1   g046(.A1(new_n241_), .A2(new_n247_), .A3(KEYINPUT8), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT8), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n238_), .A2(new_n239_), .ZN(new_n250_));
  AND3_X1   g049(.A1(new_n227_), .A2(new_n228_), .A3(new_n220_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n220_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n250_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n244_), .A2(new_n246_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n249_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n210_), .B(new_n234_), .C1(new_n248_), .C2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT12), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT8), .B1(new_n241_), .B2(new_n247_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n253_), .A2(new_n249_), .A3(new_n254_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n210_), .B1(new_n260_), .B2(new_n234_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n257_), .A2(new_n261_), .ZN(new_n262_));
  AOI211_X1 g061(.A(KEYINPUT12), .B(new_n210_), .C1(new_n260_), .C2(new_n234_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n203_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT68), .ZN(new_n265_));
  INV_X1    g064(.A(new_n256_), .ZN(new_n266_));
  OAI211_X1 g065(.A(G230gat), .B(G233gat), .C1(new_n266_), .C2(new_n261_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n268_), .B(new_n203_), .C1(new_n262_), .C2(new_n263_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n265_), .A2(new_n267_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT69), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n265_), .A2(new_n272_), .A3(new_n267_), .A4(new_n269_), .ZN(new_n273_));
  XOR2_X1   g072(.A(G120gat), .B(G148gat), .Z(new_n274_));
  XNOR2_X1  g073(.A(G176gat), .B(G204gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n276_), .B(new_n277_), .Z(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  AND4_X1   g078(.A1(new_n202_), .A2(new_n271_), .A3(new_n273_), .A4(new_n279_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n265_), .A2(new_n267_), .A3(new_n269_), .A4(new_n278_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT71), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n278_), .B1(new_n270_), .B2(KEYINPUT69), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n282_), .B1(new_n283_), .B2(new_n273_), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT72), .B1(new_n280_), .B2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n271_), .A2(new_n273_), .A3(new_n279_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n282_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT72), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n283_), .A2(new_n202_), .A3(new_n273_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n285_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT13), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n285_), .A2(new_n291_), .A3(KEYINPUT13), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT37), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT34), .ZN(new_n299_));
  XOR2_X1   g098(.A(G29gat), .B(G36gat), .Z(new_n300_));
  XOR2_X1   g099(.A(G43gat), .B(G50gat), .Z(new_n301_));
  XOR2_X1   g100(.A(new_n300_), .B(new_n301_), .Z(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT15), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n260_), .A2(new_n234_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n260_), .A2(new_n302_), .A3(new_n234_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT73), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n299_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  AOI211_X1 g108(.A(KEYINPUT73), .B(KEYINPUT34), .C1(new_n305_), .C2(new_n306_), .ZN(new_n310_));
  OAI211_X1 g109(.A(G232gat), .B(G233gat), .C1(new_n309_), .C2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n307_), .A2(new_n308_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT34), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G232gat), .A2(G233gat), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n307_), .A2(new_n308_), .A3(new_n299_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n311_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT35), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n307_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n317_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n311_), .A2(new_n316_), .A3(KEYINPUT35), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G190gat), .B(G218gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT74), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G134gat), .B(G162gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT36), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT75), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n321_), .A2(new_n322_), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT76), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n298_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n326_), .B(KEYINPUT36), .ZN(new_n333_));
  INV_X1    g132(.A(new_n322_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n319_), .B1(new_n311_), .B2(new_n316_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n333_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n330_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n332_), .A2(new_n337_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n336_), .B(new_n330_), .C1(new_n331_), .C2(new_n298_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G231gat), .A2(G233gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n210_), .B(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT77), .B(G1gat), .ZN(new_n343_));
  INV_X1    g142(.A(G8gat), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT14), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G15gat), .B(G22gat), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G1gat), .B(G8gat), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n347_), .A2(new_n348_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  XOR2_X1   g150(.A(new_n342_), .B(new_n351_), .Z(new_n352_));
  XOR2_X1   g151(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT79), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G127gat), .B(G155gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(G183gat), .B(G211gat), .Z(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n358_), .A2(KEYINPUT17), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n352_), .A2(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n358_), .A2(KEYINPUT17), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n352_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n340_), .A2(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n297_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n302_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n351_), .B(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G229gat), .A2(G233gat), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n303_), .A2(new_n351_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n369_), .B1(new_n351_), .B2(new_n366_), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n367_), .A2(new_n369_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G113gat), .B(G141gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT80), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G169gat), .B(G197gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n372_), .B(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT86), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G71gat), .B(G99gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(G43gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(KEYINPUT82), .B(G15gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G227gat), .A2(G233gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT25), .B(G183gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT26), .B(G190gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  OR2_X1    g187(.A1(G169gat), .A2(G176gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G169gat), .A2(G176gat), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n389_), .A2(KEYINPUT24), .A3(new_n390_), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n388_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT81), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G183gat), .A2(G190gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT23), .ZN(new_n395_));
  OR2_X1    g194(.A1(new_n389_), .A2(KEYINPUT24), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n388_), .A2(new_n391_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT81), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n393_), .A2(new_n397_), .A3(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n395_), .B1(G183gat), .B2(G190gat), .ZN(new_n402_));
  INV_X1    g201(.A(new_n390_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT22), .B(G169gat), .ZN(new_n404_));
  INV_X1    g203(.A(G176gat), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n403_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n402_), .A2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n401_), .A2(KEYINPUT30), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(KEYINPUT30), .B1(new_n401_), .B2(new_n407_), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT83), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n410_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT83), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n412_), .A2(new_n413_), .A3(new_n408_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n385_), .A2(new_n411_), .A3(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT85), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n384_), .A2(new_n413_), .A3(new_n412_), .A4(new_n408_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT84), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G127gat), .B(G134gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G113gat), .B(G120gat), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n419_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n420_), .B(new_n421_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n422_), .B1(new_n423_), .B2(new_n419_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT31), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n418_), .A2(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n416_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  AOI211_X1 g227(.A(new_n416_), .B(new_n425_), .C1(new_n415_), .C2(new_n417_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n378_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G22gat), .B(G50gat), .ZN(new_n431_));
  OR2_X1    g230(.A1(G141gat), .A2(G148gat), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT2), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G141gat), .A2(G148gat), .ZN(new_n434_));
  AOI22_X1  g233(.A1(new_n432_), .A2(KEYINPUT3), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n435_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(G141gat), .A2(G148gat), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n437_), .A2(KEYINPUT88), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT3), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n439_), .B1(new_n437_), .B2(KEYINPUT88), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT89), .ZN(new_n441_));
  OR3_X1    g240(.A1(new_n438_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n441_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n436_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(G155gat), .ZN(new_n445_));
  INV_X1    g244(.A(G162gat), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(G155gat), .A2(G162gat), .ZN(new_n448_));
  OR2_X1    g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  OR2_X1    g248(.A1(new_n444_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT1), .ZN(new_n451_));
  AOI211_X1 g250(.A(KEYINPUT87), .B(new_n448_), .C1(new_n447_), .C2(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n452_), .B1(new_n451_), .B2(new_n447_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n447_), .A2(KEYINPUT87), .A3(new_n451_), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n432_), .A2(new_n434_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n453_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n450_), .A2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n431_), .B1(new_n457_), .B2(KEYINPUT29), .ZN(new_n458_));
  XOR2_X1   g257(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n459_));
  INV_X1    g258(.A(KEYINPUT29), .ZN(new_n460_));
  INV_X1    g259(.A(new_n431_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n450_), .A2(new_n460_), .A3(new_n456_), .A4(new_n461_), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n458_), .A2(new_n459_), .A3(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n459_), .B1(new_n458_), .B2(new_n462_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G78gat), .B(G106gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT95), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT92), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(G233gat), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n468_), .A2(G233gat), .ZN(new_n471_));
  OAI21_X1  g270(.A(G228gat), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(G197gat), .B(G204gat), .Z(new_n474_));
  INV_X1    g273(.A(KEYINPUT94), .ZN(new_n475_));
  OR3_X1    g274(.A1(new_n474_), .A2(new_n475_), .A3(KEYINPUT21), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n475_), .B1(new_n474_), .B2(KEYINPUT21), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n474_), .A2(KEYINPUT21), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G211gat), .B(G218gat), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .A4(new_n479_), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n478_), .A2(new_n479_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT93), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n444_), .A2(new_n449_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n456_), .ZN(new_n487_));
  OAI211_X1 g286(.A(KEYINPUT91), .B(KEYINPUT29), .C1(new_n486_), .C2(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n473_), .B1(new_n485_), .B2(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT91), .B1(new_n472_), .B2(new_n484_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n482_), .A2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n491_), .B1(new_n457_), .B2(KEYINPUT29), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n467_), .B1(new_n489_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT96), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n465_), .A2(new_n494_), .ZN(new_n495_));
  OR3_X1    g294(.A1(new_n489_), .A2(new_n492_), .A3(new_n467_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(new_n493_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n465_), .A2(new_n494_), .A3(new_n493_), .A4(new_n496_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n427_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n501_), .A2(new_n418_), .A3(new_n425_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n429_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(KEYINPUT86), .A3(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n430_), .A2(new_n500_), .A3(new_n504_), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n498_), .A2(new_n499_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n428_), .A2(new_n429_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n505_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n392_), .A2(new_n397_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n402_), .A2(KEYINPUT98), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(new_n406_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n402_), .A2(KEYINPUT98), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n510_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(new_n482_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT99), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n401_), .A2(new_n407_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(new_n483_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n514_), .A2(KEYINPUT99), .A3(new_n482_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n517_), .A2(new_n520_), .A3(KEYINPUT20), .A4(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G226gat), .A2(G233gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n522_), .A2(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(G8gat), .B(G36gat), .Z(new_n527_));
  XNOR2_X1  g326(.A(G64gat), .B(G92gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  XOR2_X1   g328(.A(KEYINPUT100), .B(KEYINPUT18), .Z(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n519_), .A2(new_n483_), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT20), .B1(new_n514_), .B2(new_n482_), .ZN(new_n533_));
  OR3_X1    g332(.A1(new_n532_), .A2(new_n525_), .A3(new_n533_), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n526_), .A2(new_n531_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n520_), .A2(KEYINPUT20), .ZN(new_n537_));
  INV_X1    g336(.A(new_n525_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n537_), .A2(new_n517_), .A3(new_n538_), .A4(new_n521_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n525_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n531_), .B(KEYINPUT102), .Z(new_n542_));
  OAI211_X1 g341(.A(new_n536_), .B(KEYINPUT27), .C1(new_n541_), .C2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT103), .B(KEYINPUT27), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n531_), .B1(new_n526_), .B2(new_n534_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n544_), .B1(new_n535_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G1gat), .B(G29gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(G85gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(KEYINPUT0), .B(G57gat), .ZN(new_n550_));
  XOR2_X1   g349(.A(new_n549_), .B(new_n550_), .Z(new_n551_));
  NAND2_X1  g350(.A1(G225gat), .A2(G233gat), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT4), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n450_), .A2(new_n423_), .A3(new_n456_), .ZN(new_n555_));
  AOI22_X1  g354(.A1(new_n555_), .A2(KEYINPUT101), .B1(new_n457_), .B2(new_n424_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT101), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n450_), .A2(new_n557_), .A3(new_n423_), .A4(new_n456_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n554_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(KEYINPUT4), .B1(new_n457_), .B2(new_n424_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n553_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n556_), .A2(new_n558_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(new_n552_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n551_), .B1(new_n561_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n561_), .A2(new_n551_), .A3(new_n564_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n547_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n509_), .A2(new_n569_), .ZN(new_n570_));
  AND3_X1   g369(.A1(new_n506_), .A2(new_n430_), .A3(new_n504_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT33), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n567_), .A2(new_n572_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n561_), .A2(new_n564_), .A3(KEYINPUT33), .A4(new_n551_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n551_), .B1(new_n563_), .B2(new_n553_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n552_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n535_), .A2(new_n545_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n573_), .A2(new_n574_), .A3(new_n577_), .A4(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n531_), .A2(KEYINPUT32), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n580_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n526_), .A2(new_n534_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n581_), .B1(new_n582_), .B2(new_n580_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n567_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n583_), .B1(new_n584_), .B2(new_n565_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n579_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n571_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n570_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n365_), .A2(new_n377_), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n590_), .A2(new_n568_), .A3(new_n343_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(KEYINPUT105), .A2(KEYINPUT38), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n593_), .B1(new_n594_), .B2(new_n591_), .ZN(new_n595_));
  AOI22_X1  g394(.A1(new_n509_), .A2(new_n569_), .B1(new_n571_), .B2(new_n586_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n337_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n363_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n596_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n377_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n600_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT104), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(new_n568_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n595_), .B1(G1gat), .B2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT106), .ZN(G1324gat));
  INV_X1    g405(.A(new_n547_), .ZN(new_n607_));
  OAI21_X1  g406(.A(G8gat), .B1(new_n602_), .B2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT39), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n590_), .A2(new_n344_), .A3(new_n547_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT40), .Z(G1325gat));
  NAND2_X1  g411(.A1(new_n430_), .A2(new_n504_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n603_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(G15gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT41), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n616_), .A2(KEYINPUT107), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(KEYINPUT107), .ZN(new_n618_));
  INV_X1    g417(.A(new_n613_), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n589_), .A2(G15gat), .A3(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT108), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n617_), .A2(new_n618_), .A3(new_n621_), .ZN(G1326gat));
  INV_X1    g421(.A(G22gat), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n623_), .B1(new_n603_), .B2(new_n500_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT42), .Z(new_n625_));
  NAND3_X1  g424(.A1(new_n590_), .A2(new_n623_), .A3(new_n500_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(G1327gat));
  NOR3_X1   g426(.A1(new_n596_), .A2(new_n337_), .A3(new_n363_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(new_n601_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n568_), .ZN(new_n630_));
  OR3_X1    g429(.A1(new_n629_), .A2(G29gat), .A3(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n338_), .A2(new_n339_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT43), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n588_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(KEYINPUT43), .B1(new_n596_), .B2(new_n340_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n363_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  AOI211_X1 g435(.A(KEYINPUT109), .B(KEYINPUT44), .C1(new_n636_), .C2(new_n601_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT109), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n634_), .A2(new_n635_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n639_), .A2(new_n601_), .A3(new_n598_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT44), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n638_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n637_), .A2(new_n642_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n639_), .A2(KEYINPUT44), .A3(new_n601_), .A4(new_n598_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT110), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n636_), .A2(KEYINPUT110), .A3(KEYINPUT44), .A4(new_n601_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n643_), .A2(new_n568_), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT111), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n649_), .A2(new_n650_), .A3(G29gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n649_), .B2(G29gat), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n631_), .B1(new_n651_), .B2(new_n652_), .ZN(G1328gat));
  NAND2_X1  g452(.A1(new_n640_), .A2(new_n641_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT109), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n640_), .A2(new_n638_), .A3(new_n641_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n648_), .A2(new_n655_), .A3(new_n547_), .A4(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT112), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n643_), .A2(KEYINPUT112), .A3(new_n547_), .A4(new_n648_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n659_), .A2(G36gat), .A3(new_n660_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n629_), .A2(G36gat), .A3(new_n607_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT45), .Z(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT46), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n661_), .A2(KEYINPUT46), .A3(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1329gat));
  NAND3_X1  g467(.A1(new_n643_), .A2(new_n507_), .A3(new_n648_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(G43gat), .ZN(new_n670_));
  OR3_X1    g469(.A1(new_n629_), .A2(G43gat), .A3(new_n619_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT47), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n672_), .B(new_n673_), .ZN(G1330gat));
  NAND4_X1  g473(.A1(new_n643_), .A2(G50gat), .A3(new_n500_), .A4(new_n648_), .ZN(new_n675_));
  INV_X1    g474(.A(G50gat), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n676_), .B1(new_n629_), .B2(new_n506_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n675_), .A2(new_n677_), .ZN(G1331gat));
  NOR2_X1   g477(.A1(new_n296_), .A2(new_n377_), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n679_), .A2(new_n599_), .A3(G57gat), .A4(new_n568_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n296_), .A2(new_n364_), .ZN(new_n681_));
  AOI211_X1 g480(.A(new_n377_), .B(new_n596_), .C1(new_n681_), .C2(KEYINPUT113), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n682_), .B1(KEYINPUT113), .B2(new_n681_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n683_), .A2(KEYINPUT114), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n568_), .B1(new_n683_), .B2(KEYINPUT114), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n680_), .B1(new_n686_), .B2(G57gat), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT115), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  OAI211_X1 g488(.A(KEYINPUT115), .B(new_n680_), .C1(new_n686_), .C2(G57gat), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1332gat));
  NAND2_X1  g490(.A1(new_n679_), .A2(new_n599_), .ZN(new_n692_));
  OAI21_X1  g491(.A(G64gat), .B1(new_n692_), .B2(new_n607_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT48), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n607_), .A2(G64gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n694_), .B1(new_n683_), .B2(new_n695_), .ZN(G1333gat));
  OAI21_X1  g495(.A(G71gat), .B1(new_n692_), .B2(new_n619_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT49), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n619_), .A2(G71gat), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n698_), .B1(new_n683_), .B2(new_n699_), .ZN(G1334gat));
  OAI21_X1  g499(.A(G78gat), .B1(new_n692_), .B2(new_n506_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT50), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n506_), .A2(G78gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n683_), .B2(new_n703_), .ZN(G1335gat));
  NAND2_X1  g503(.A1(new_n636_), .A2(new_n679_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n705_), .A2(new_n630_), .A3(new_n215_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n679_), .A2(new_n628_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT116), .Z(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(new_n568_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n706_), .B1(new_n709_), .B2(new_n211_), .ZN(G1336gat));
  NAND3_X1  g509(.A1(new_n708_), .A2(new_n212_), .A3(new_n547_), .ZN(new_n711_));
  OAI21_X1  g510(.A(G92gat), .B1(new_n705_), .B2(new_n607_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1337gat));
  NOR3_X1   g512(.A1(new_n428_), .A2(new_n231_), .A3(new_n429_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n636_), .A2(new_n613_), .A3(new_n679_), .ZN(new_n715_));
  AOI22_X1  g514(.A1(new_n708_), .A2(new_n714_), .B1(G99gat), .B2(new_n715_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g516(.A1(new_n708_), .A2(new_n237_), .A3(new_n500_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n636_), .A2(new_n500_), .A3(new_n679_), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n719_), .A2(KEYINPUT117), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT52), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n237_), .B1(new_n719_), .B2(KEYINPUT117), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n720_), .A2(new_n721_), .A3(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n721_), .B1(new_n720_), .B2(new_n722_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n718_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g525(.A(KEYINPUT122), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n508_), .A2(new_n630_), .A3(new_n547_), .ZN(new_n728_));
  XOR2_X1   g527(.A(new_n728_), .B(KEYINPUT119), .Z(new_n729_));
  INV_X1    g528(.A(KEYINPUT59), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n296_), .A2(new_n600_), .A3(new_n363_), .A4(new_n340_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n732_), .B(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n376_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n368_), .B1(new_n351_), .B2(new_n366_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n370_), .A2(new_n737_), .ZN(new_n738_));
  AOI22_X1  g537(.A1(new_n372_), .A2(new_n376_), .B1(new_n736_), .B2(new_n738_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n281_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT55), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n264_), .A2(new_n741_), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n262_), .A2(new_n203_), .A3(new_n263_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n265_), .A2(new_n741_), .A3(new_n269_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n746_), .A2(KEYINPUT56), .A3(new_n279_), .ZN(new_n747_));
  AOI21_X1  g546(.A(KEYINPUT56), .B1(new_n746_), .B2(new_n279_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n740_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT58), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  OAI211_X1 g550(.A(KEYINPUT58), .B(new_n740_), .C1(new_n747_), .C2(new_n748_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n338_), .A2(new_n751_), .A3(new_n339_), .A4(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n285_), .A2(new_n291_), .A3(new_n739_), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n377_), .B(new_n281_), .C1(new_n747_), .C2(new_n748_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n597_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n753_), .B1(new_n756_), .B2(KEYINPUT57), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT120), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT57), .ZN(new_n760_));
  AOI211_X1 g559(.A(new_n760_), .B(new_n597_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  OAI211_X1 g561(.A(KEYINPUT120), .B(new_n753_), .C1(new_n756_), .C2(KEYINPUT57), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n759_), .A2(new_n762_), .A3(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n598_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n735_), .B1(new_n765_), .B2(KEYINPUT121), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n761_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n363_), .B1(new_n767_), .B2(new_n763_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT121), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n731_), .B1(new_n766_), .B2(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n732_), .B(new_n733_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n757_), .A2(new_n761_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n772_), .B1(new_n363_), .B2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n730_), .B1(new_n774_), .B2(new_n729_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n727_), .B1(new_n771_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n731_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n770_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n772_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n777_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n773_), .A2(new_n363_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n735_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n729_), .ZN(new_n783_));
  OAI21_X1  g582(.A(KEYINPUT59), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n780_), .A2(KEYINPUT122), .A3(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n776_), .A2(new_n377_), .A3(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(G113gat), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n782_), .A2(new_n783_), .ZN(new_n788_));
  INV_X1    g587(.A(G113gat), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(new_n789_), .A3(new_n377_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n787_), .A2(new_n790_), .ZN(G1340gat));
  NOR2_X1   g590(.A1(new_n296_), .A2(KEYINPUT60), .ZN(new_n792_));
  MUX2_X1   g591(.A(new_n792_), .B(KEYINPUT60), .S(G120gat), .Z(new_n793_));
  NAND2_X1  g592(.A1(new_n788_), .A2(new_n793_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n771_), .A2(new_n296_), .A3(new_n775_), .ZN(new_n795_));
  INV_X1    g594(.A(G120gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n794_), .B1(new_n795_), .B2(new_n796_), .ZN(G1341gat));
  NAND3_X1  g596(.A1(new_n776_), .A2(new_n363_), .A3(new_n785_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(G127gat), .ZN(new_n799_));
  INV_X1    g598(.A(G127gat), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n788_), .A2(new_n800_), .A3(new_n363_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(G1342gat));
  NAND3_X1  g601(.A1(new_n776_), .A2(new_n632_), .A3(new_n785_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(G134gat), .ZN(new_n804_));
  INV_X1    g603(.A(G134gat), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n788_), .A2(new_n805_), .A3(new_n597_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(G1343gat));
  NOR3_X1   g606(.A1(new_n505_), .A2(new_n630_), .A3(new_n547_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT123), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n782_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n377_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n297_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g613(.A1(new_n810_), .A2(new_n363_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(KEYINPUT61), .B(G155gat), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n815_), .B(new_n816_), .ZN(G1346gat));
  INV_X1    g616(.A(new_n810_), .ZN(new_n818_));
  OAI21_X1  g617(.A(G162gat), .B1(new_n818_), .B2(new_n340_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n810_), .A2(new_n446_), .A3(new_n597_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(G1347gat));
  NAND3_X1  g620(.A1(new_n613_), .A2(new_n630_), .A3(new_n547_), .ZN(new_n822_));
  AOI211_X1 g621(.A(new_n500_), .B(new_n822_), .C1(new_n766_), .C2(new_n770_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n823_), .A2(new_n377_), .A3(new_n404_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n822_), .A2(new_n500_), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n377_), .B(new_n825_), .C1(new_n778_), .C2(new_n779_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(G169gat), .ZN(new_n827_));
  XNOR2_X1  g626(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT125), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n827_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n829_), .A2(new_n830_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n827_), .A2(new_n832_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n824_), .B1(new_n835_), .B2(new_n836_), .ZN(G1348gat));
  AOI21_X1  g636(.A(G176gat), .B1(new_n823_), .B2(new_n297_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n782_), .A2(new_n500_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n296_), .A2(new_n405_), .A3(new_n822_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n838_), .B1(new_n839_), .B2(new_n840_), .ZN(G1349gat));
  NOR2_X1   g640(.A1(new_n822_), .A2(new_n598_), .ZN(new_n842_));
  AOI21_X1  g641(.A(G183gat), .B1(new_n839_), .B2(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n598_), .A2(new_n386_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n843_), .B1(new_n823_), .B2(new_n844_), .ZN(G1350gat));
  NAND2_X1  g644(.A1(new_n823_), .A2(new_n632_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(G190gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n823_), .A2(new_n387_), .A3(new_n597_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(G1351gat));
  NOR4_X1   g648(.A1(new_n782_), .A2(new_n568_), .A3(new_n505_), .A4(new_n607_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n377_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n297_), .ZN(new_n853_));
  INV_X1    g652(.A(G204gat), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(KEYINPUT126), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n853_), .B(new_n855_), .ZN(G1353gat));
  NAND2_X1  g655(.A1(new_n850_), .A2(new_n363_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n858_));
  AND2_X1   g657(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n857_), .A2(new_n858_), .A3(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n860_), .B1(new_n857_), .B2(new_n858_), .ZN(G1354gat));
  INV_X1    g660(.A(G218gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n850_), .A2(new_n862_), .A3(new_n597_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n850_), .A2(new_n632_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(new_n862_), .ZN(G1355gat));
endmodule


