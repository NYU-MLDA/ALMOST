//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 0 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 0 0 0 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n785_, new_n786_, new_n787_, new_n789_, new_n790_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n797_, new_n799_,
    new_n800_, new_n802_, new_n803_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n823_, new_n824_, new_n825_, new_n827_, new_n828_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(KEYINPUT6), .ZN(new_n202_));
  AND2_X1   g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  OR3_X1    g003(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(G85gat), .B(G92gat), .Z(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n207_), .A2(KEYINPUT65), .A3(new_n208_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n211_), .A2(KEYINPUT8), .A3(new_n212_), .ZN(new_n213_));
  XOR2_X1   g012(.A(KEYINPUT10), .B(G99gat), .Z(new_n214_));
  INV_X1    g013(.A(G106gat), .ZN(new_n215_));
  AOI22_X1  g014(.A1(KEYINPUT9), .A2(new_n208_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G85gat), .ZN(new_n217_));
  INV_X1    g016(.A(G92gat), .ZN(new_n218_));
  OR3_X1    g017(.A1(new_n217_), .A2(new_n218_), .A3(KEYINPUT9), .ZN(new_n219_));
  AND3_X1   g018(.A1(new_n204_), .A2(new_n216_), .A3(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(KEYINPUT65), .B1(new_n207_), .B2(new_n208_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT8), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n220_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n213_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G29gat), .B(G36gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G43gat), .B(G50gat), .ZN(new_n226_));
  XOR2_X1   g025(.A(new_n225_), .B(new_n226_), .Z(new_n227_));
  XOR2_X1   g026(.A(new_n227_), .B(KEYINPUT15), .Z(new_n228_));
  NAND2_X1  g027(.A1(new_n224_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n227_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n213_), .A2(new_n230_), .A3(new_n223_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G232gat), .A2(G233gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT34), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n232_), .A2(KEYINPUT35), .A3(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT70), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(KEYINPUT35), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n234_), .A2(KEYINPUT35), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n229_), .A2(new_n237_), .A3(new_n238_), .A4(new_n231_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n235_), .A2(new_n236_), .A3(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G190gat), .B(G218gat), .ZN(new_n241_));
  INV_X1    g040(.A(G162gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT69), .B(G134gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n245_), .A2(KEYINPUT36), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n240_), .A2(new_n247_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n235_), .A2(new_n236_), .A3(new_n239_), .A4(new_n246_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT36), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n251_), .B1(new_n235_), .B2(new_n239_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(new_n245_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n250_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT71), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n254_), .A2(new_n255_), .A3(KEYINPUT37), .ZN(new_n256_));
  AOI22_X1  g055(.A1(new_n248_), .A2(new_n249_), .B1(new_n245_), .B2(new_n252_), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n255_), .A2(KEYINPUT37), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n255_), .A2(KEYINPUT37), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n257_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n256_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G57gat), .B(G64gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT66), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n263_), .A2(KEYINPUT11), .ZN(new_n264_));
  XOR2_X1   g063(.A(G71gat), .B(G78gat), .Z(new_n265_));
  OR2_X1    g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n263_), .A2(KEYINPUT11), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n265_), .B1(new_n264_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G15gat), .B(G22gat), .ZN(new_n270_));
  INV_X1    g069(.A(G1gat), .ZN(new_n271_));
  INV_X1    g070(.A(G8gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT14), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G1gat), .B(G8gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G231gat), .A2(G233gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n269_), .B(new_n278_), .Z(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(G183gat), .B(G211gat), .Z(new_n281_));
  XNOR2_X1  g080(.A(G127gat), .B(G155gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT17), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n286_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n280_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  AND2_X1   g088(.A1(new_n280_), .A2(new_n287_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n261_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT73), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n276_), .A2(new_n227_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT74), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n276_), .A2(new_n227_), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G229gat), .A2(G233gat), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n228_), .A2(new_n276_), .ZN(new_n301_));
  AND3_X1   g100(.A1(new_n301_), .A2(new_n296_), .A3(new_n299_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G113gat), .B(G141gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G169gat), .B(G197gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  OR3_X1    g104(.A1(new_n300_), .A2(new_n302_), .A3(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n305_), .B1(new_n300_), .B2(new_n302_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n224_), .A2(new_n269_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT67), .ZN(new_n311_));
  INV_X1    g110(.A(new_n269_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n312_), .A2(new_n223_), .A3(new_n213_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n311_), .B(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(G230gat), .ZN(new_n315_));
  INV_X1    g114(.A(G233gat), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n314_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n310_), .A2(new_n313_), .A3(KEYINPUT12), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT12), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n224_), .A2(new_n320_), .A3(new_n269_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G230gat), .A2(G233gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(G176gat), .B(G204gat), .Z(new_n325_));
  XNOR2_X1  g124(.A(G120gat), .B(G148gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n318_), .A2(new_n324_), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n329_), .B1(new_n318_), .B2(new_n324_), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT13), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n332_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT13), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(new_n335_), .A3(new_n330_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n309_), .B1(new_n333_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G228gat), .A2(G233gat), .ZN(new_n338_));
  XOR2_X1   g137(.A(G197gat), .B(G204gat), .Z(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT21), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G211gat), .B(G218gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G197gat), .B(G204gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT21), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n340_), .A2(new_n341_), .A3(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n342_), .A2(new_n343_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n341_), .ZN(new_n347_));
  AOI21_X1  g146(.A(KEYINPUT83), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT83), .ZN(new_n349_));
  NOR4_X1   g148(.A1(new_n342_), .A2(new_n341_), .A3(new_n349_), .A4(new_n343_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n345_), .B1(new_n348_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(G141gat), .ZN(new_n352_));
  INV_X1    g151(.A(G148gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G141gat), .A2(G148gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(G155gat), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n358_), .A2(new_n242_), .A3(KEYINPUT79), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n360_), .B1(G155gat), .B2(G162gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G155gat), .A2(G162gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT1), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT80), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n362_), .A2(KEYINPUT80), .A3(new_n364_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n363_), .A2(KEYINPUT1), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n357_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n352_), .A2(new_n353_), .A3(KEYINPUT3), .ZN(new_n372_));
  AOI21_X1  g171(.A(KEYINPUT3), .B1(new_n352_), .B2(new_n353_), .ZN(new_n373_));
  OAI22_X1  g172(.A1(new_n372_), .A2(new_n373_), .B1(KEYINPUT81), .B2(KEYINPUT2), .ZN(new_n374_));
  NAND2_X1  g173(.A1(KEYINPUT81), .A2(KEYINPUT2), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n355_), .B(new_n375_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n363_), .B(new_n362_), .C1(new_n374_), .C2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n371_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT29), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n338_), .B(new_n351_), .C1(new_n379_), .C2(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n380_), .B1(new_n371_), .B2(new_n377_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n351_), .ZN(new_n383_));
  OAI211_X1 g182(.A(G228gat), .B(G233gat), .C1(new_n382_), .C2(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(G78gat), .B(G106gat), .Z(new_n385_));
  NAND3_X1  g184(.A1(new_n381_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT84), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n381_), .A2(new_n384_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n385_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n387_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  AOI211_X1 g189(.A(KEYINPUT84), .B(new_n385_), .C1(new_n381_), .C2(new_n384_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n386_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G22gat), .B(G50gat), .ZN(new_n393_));
  XOR2_X1   g192(.A(KEYINPUT82), .B(KEYINPUT28), .Z(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n395_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n379_), .A2(new_n380_), .A3(new_n395_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n393_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n398_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n393_), .ZN(new_n401_));
  NOR3_X1   g200(.A1(new_n400_), .A2(new_n401_), .A3(new_n396_), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n399_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n392_), .A2(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n399_), .A2(new_n402_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n386_), .A2(KEYINPUT86), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT86), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n381_), .A2(new_n384_), .A3(new_n407_), .A4(new_n385_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n388_), .A2(new_n389_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT85), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT85), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n388_), .A2(new_n412_), .A3(new_n389_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n405_), .A2(new_n409_), .A3(new_n411_), .A4(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n404_), .A2(new_n414_), .ZN(new_n415_));
  NOR3_X1   g214(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n416_));
  AND3_X1   g215(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n417_));
  AOI21_X1  g216(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n418_));
  NOR3_X1   g217(.A1(new_n416_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(G190gat), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT26), .B1(new_n420_), .B2(KEYINPUT75), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT75), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT26), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(new_n423_), .A3(G190gat), .ZN(new_n424_));
  NOR2_X1   g223(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n425_));
  AND2_X1   g224(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n421_), .B(new_n424_), .C1(new_n425_), .C2(new_n426_), .ZN(new_n427_));
  OR2_X1    g226(.A1(G169gat), .A2(G176gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G169gat), .A2(G176gat), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(KEYINPUT24), .A3(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n419_), .A2(new_n427_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n418_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n433_));
  OR2_X1    g232(.A1(G183gat), .A2(G190gat), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n432_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(G176gat), .ZN(new_n436_));
  AND2_X1   g235(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n437_));
  NOR2_X1   g236(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n436_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n435_), .A2(new_n439_), .A3(new_n429_), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n431_), .A2(KEYINPUT76), .A3(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(KEYINPUT76), .B1(new_n431_), .B2(new_n440_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT78), .B(KEYINPUT31), .ZN(new_n444_));
  XOR2_X1   g243(.A(new_n444_), .B(KEYINPUT30), .Z(new_n445_));
  XNOR2_X1  g244(.A(new_n443_), .B(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G127gat), .B(G134gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G113gat), .B(G120gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G227gat), .A2(G233gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n446_), .B(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G15gat), .B(G43gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT77), .ZN(new_n454_));
  XOR2_X1   g253(.A(G71gat), .B(G99gat), .Z(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n452_), .B(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n415_), .A2(new_n457_), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n362_), .A2(KEYINPUT80), .A3(new_n364_), .ZN(new_n459_));
  AOI21_X1  g258(.A(KEYINPUT80), .B1(new_n362_), .B2(new_n364_), .ZN(new_n460_));
  NOR3_X1   g259(.A1(new_n459_), .A2(new_n460_), .A3(new_n370_), .ZN(new_n461_));
  OAI211_X1 g260(.A(KEYINPUT90), .B(new_n377_), .C1(new_n461_), .C2(new_n356_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n449_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n371_), .A2(KEYINPUT90), .A3(new_n377_), .A4(new_n449_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(KEYINPUT4), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G225gat), .A2(G233gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT91), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT4), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n378_), .A2(new_n469_), .A3(new_n463_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n466_), .A2(new_n468_), .A3(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n464_), .A2(new_n467_), .A3(new_n465_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G1gat), .B(G29gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(G85gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT0), .B(G57gat), .ZN(new_n476_));
  XOR2_X1   g275(.A(new_n475_), .B(new_n476_), .Z(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n473_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT95), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n471_), .A2(new_n472_), .A3(new_n477_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n473_), .A2(KEYINPUT95), .A3(new_n478_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT27), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n351_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n349_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n346_), .A2(KEYINPUT83), .A3(new_n347_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT88), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n432_), .A2(new_n433_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n490_), .B1(new_n491_), .B2(new_n416_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT26), .B(G190gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n493_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n416_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n495_), .A2(new_n432_), .A3(KEYINPUT88), .A4(new_n433_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n492_), .A2(new_n494_), .A3(new_n430_), .A4(new_n496_), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n489_), .A2(new_n497_), .A3(new_n345_), .A4(new_n440_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n486_), .A2(KEYINPUT20), .A3(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G226gat), .A2(G233gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n499_), .A2(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(KEYINPUT89), .B(KEYINPUT18), .Z(new_n505_));
  XNOR2_X1  g304(.A(G8gat), .B(G36gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G64gat), .B(G92gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n442_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n431_), .A2(KEYINPUT76), .A3(new_n440_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n383_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n497_), .A2(new_n440_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(new_n351_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n512_), .A2(KEYINPUT20), .A3(new_n514_), .A4(new_n502_), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n504_), .A2(new_n509_), .A3(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n509_), .B1(new_n504_), .B2(new_n515_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n485_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n517_), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n499_), .A2(new_n502_), .ZN(new_n520_));
  AND4_X1   g319(.A1(KEYINPUT20), .A2(new_n512_), .A3(new_n503_), .A4(new_n514_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n509_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n519_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n518_), .B1(new_n524_), .B2(new_n485_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n458_), .A2(new_n484_), .A3(new_n526_), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n523_), .A2(KEYINPUT32), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n528_), .B(KEYINPUT94), .Z(new_n529_));
  NAND2_X1  g328(.A1(new_n504_), .A2(new_n515_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n528_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n482_), .A2(new_n483_), .A3(new_n531_), .A4(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(KEYINPUT92), .B(KEYINPUT33), .Z(new_n534_));
  NAND2_X1  g333(.A1(new_n481_), .A2(new_n534_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n471_), .A2(KEYINPUT33), .A3(new_n472_), .A4(new_n477_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n516_), .A2(new_n517_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n466_), .A2(new_n467_), .A3(new_n470_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n464_), .A2(new_n465_), .A3(new_n468_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n538_), .A2(new_n478_), .A3(new_n539_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .A4(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT93), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n504_), .A2(new_n515_), .A3(new_n509_), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n540_), .A2(new_n519_), .A3(new_n544_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n545_), .A2(KEYINPUT93), .A3(new_n536_), .A4(new_n535_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n533_), .A2(new_n543_), .A3(new_n546_), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n404_), .A2(new_n414_), .ZN(new_n548_));
  AOI22_X1  g347(.A1(new_n404_), .A2(new_n414_), .B1(new_n483_), .B2(new_n482_), .ZN(new_n549_));
  AOI22_X1  g348(.A1(new_n547_), .A2(new_n548_), .B1(new_n549_), .B2(new_n526_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n457_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n527_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n337_), .A2(new_n552_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n294_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n484_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n554_), .A2(new_n271_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT38), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n558_), .B(KEYINPUT97), .Z(new_n559_));
  NOR2_X1   g358(.A1(new_n254_), .A2(new_n291_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n553_), .A2(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(G1gat), .B1(new_n561_), .B2(new_n484_), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n554_), .A2(KEYINPUT38), .A3(new_n271_), .A4(new_n555_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT96), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n559_), .A2(new_n562_), .A3(new_n564_), .ZN(G1324gat));
  NAND3_X1  g364(.A1(new_n554_), .A2(new_n272_), .A3(new_n525_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT98), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(G8gat), .B1(new_n561_), .B2(new_n526_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT39), .ZN(new_n570_));
  XNOR2_X1  g369(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n568_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n571_), .B1(new_n568_), .B2(new_n570_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(G1325gat));
  INV_X1    g373(.A(G15gat), .ZN(new_n575_));
  INV_X1    g374(.A(new_n561_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n575_), .B1(new_n576_), .B2(new_n551_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT100), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT41), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n577_), .A2(new_n578_), .ZN(new_n582_));
  OR3_X1    g381(.A1(new_n580_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n581_), .B1(new_n580_), .B2(new_n582_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n554_), .A2(new_n575_), .A3(new_n551_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n583_), .A2(new_n584_), .A3(new_n585_), .ZN(G1326gat));
  OAI21_X1  g385(.A(G22gat), .B1(new_n561_), .B2(new_n548_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT42), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n548_), .A2(G22gat), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n589_), .B(KEYINPUT101), .Z(new_n590_));
  NAND2_X1  g389(.A1(new_n554_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n588_), .A2(new_n591_), .ZN(G1327gat));
  NOR2_X1   g391(.A1(new_n257_), .A2(new_n292_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n553_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(G29gat), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n594_), .A2(new_n595_), .A3(new_n555_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT43), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n256_), .A2(new_n260_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n547_), .A2(new_n548_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n549_), .A2(new_n526_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n551_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  NOR4_X1   g400(.A1(new_n415_), .A2(new_n555_), .A3(new_n525_), .A4(new_n457_), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n597_), .B(new_n598_), .C1(new_n601_), .C2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT102), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n599_), .A2(new_n600_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n602_), .B1(new_n605_), .B2(new_n457_), .ZN(new_n606_));
  OAI21_X1  g405(.A(KEYINPUT43), .B1(new_n606_), .B2(new_n261_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT102), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n552_), .A2(new_n608_), .A3(new_n597_), .A4(new_n598_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n604_), .A2(new_n607_), .A3(new_n609_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n337_), .A2(new_n291_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n610_), .A2(KEYINPUT44), .A3(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(KEYINPUT44), .B1(new_n610_), .B2(new_n611_), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n612_), .A2(new_n613_), .A3(new_n484_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n596_), .B1(new_n614_), .B2(new_n595_), .ZN(G1328gat));
  INV_X1    g414(.A(KEYINPUT105), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT46), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT103), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n612_), .A2(new_n613_), .A3(new_n526_), .ZN(new_n621_));
  INV_X1    g420(.A(G36gat), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n620_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n613_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n610_), .A2(KEYINPUT44), .A3(new_n611_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n624_), .A2(new_n525_), .A3(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n626_), .A2(KEYINPUT103), .A3(G36gat), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n623_), .A2(new_n627_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n337_), .A2(new_n552_), .A3(new_n622_), .A4(new_n593_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n629_), .A2(KEYINPUT104), .A3(new_n526_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT45), .ZN(new_n632_));
  OAI21_X1  g431(.A(KEYINPUT104), .B1(new_n629_), .B2(new_n526_), .ZN(new_n633_));
  AND3_X1   g432(.A1(new_n631_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n632_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n635_));
  OAI22_X1  g434(.A1(new_n634_), .A2(new_n635_), .B1(KEYINPUT105), .B2(KEYINPUT46), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n619_), .B1(new_n628_), .B2(new_n637_), .ZN(new_n638_));
  AOI211_X1 g437(.A(new_n618_), .B(new_n636_), .C1(new_n623_), .C2(new_n627_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(G1329gat));
  NAND4_X1  g439(.A1(new_n624_), .A2(G43gat), .A3(new_n551_), .A4(new_n625_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n594_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n642_), .A2(new_n457_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n641_), .B1(G43gat), .B2(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g444(.A1(new_n624_), .A2(new_n415_), .A3(new_n625_), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n646_), .A2(KEYINPUT106), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(KEYINPUT106), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n647_), .A2(G50gat), .A3(new_n648_), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n548_), .A2(G50gat), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n649_), .B1(new_n642_), .B2(new_n650_), .ZN(G1331gat));
  INV_X1    g450(.A(G57gat), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT109), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n652_), .B1(new_n555_), .B2(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n606_), .A2(new_n308_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n333_), .A2(new_n336_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n655_), .A2(new_n657_), .A3(new_n560_), .ZN(new_n658_));
  AOI211_X1 g457(.A(new_n654_), .B(new_n658_), .C1(new_n653_), .C2(new_n652_), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n655_), .B(KEYINPUT107), .Z(new_n660_));
  NOR2_X1   g459(.A1(new_n660_), .A2(new_n656_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(new_n294_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT108), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(new_n555_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n659_), .B1(new_n665_), .B2(new_n652_), .ZN(G1332gat));
  OAI21_X1  g465(.A(G64gat), .B1(new_n658_), .B2(new_n526_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT48), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n526_), .A2(G64gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(new_n662_), .B2(new_n669_), .ZN(G1333gat));
  OAI21_X1  g469(.A(G71gat), .B1(new_n658_), .B2(new_n457_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT110), .Z(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT49), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n662_), .A2(G71gat), .A3(new_n457_), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1334gat));
  OAI21_X1  g474(.A(G78gat), .B1(new_n658_), .B2(new_n548_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT50), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n548_), .A2(G78gat), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT111), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n677_), .B1(new_n662_), .B2(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT112), .ZN(G1335gat));
  AND2_X1   g480(.A1(new_n661_), .A2(new_n593_), .ZN(new_n682_));
  AOI21_X1  g481(.A(G85gat), .B1(new_n682_), .B2(new_n555_), .ZN(new_n683_));
  AND4_X1   g482(.A1(new_n309_), .A2(new_n610_), .A3(new_n657_), .A4(new_n291_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n684_), .A2(G85gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n683_), .B1(new_n555_), .B2(new_n685_), .ZN(G1336gat));
  AOI21_X1  g485(.A(G92gat), .B1(new_n682_), .B2(new_n525_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n684_), .A2(new_n525_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(G92gat), .B2(new_n688_), .ZN(G1337gat));
  NAND3_X1  g488(.A1(new_n682_), .A2(new_n551_), .A3(new_n214_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT113), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n684_), .A2(new_n551_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n691_), .B1(new_n692_), .B2(G99gat), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n692_), .A2(new_n691_), .A3(G99gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n690_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(KEYINPUT51), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT51), .ZN(new_n697_));
  OAI211_X1 g496(.A(new_n690_), .B(new_n697_), .C1(new_n693_), .C2(new_n694_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(G1338gat));
  NAND3_X1  g498(.A1(new_n682_), .A2(new_n215_), .A3(new_n415_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT52), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n684_), .A2(new_n415_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n702_), .B2(G106gat), .ZN(new_n703_));
  AOI211_X1 g502(.A(KEYINPUT52), .B(new_n215_), .C1(new_n684_), .C2(new_n415_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n700_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n700_), .B(new_n706_), .C1(new_n703_), .C2(new_n704_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1339gat));
  INV_X1    g509(.A(KEYINPUT57), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n331_), .A2(new_n332_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n299_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n301_), .A2(new_n296_), .A3(new_n713_), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n305_), .B(new_n714_), .C1(new_n298_), .C2(new_n713_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n306_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT118), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n716_), .B(new_n717_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n712_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT116), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT55), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n324_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n319_), .A2(new_n317_), .A3(new_n321_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n317_), .B1(new_n319_), .B2(new_n321_), .ZN(new_n724_));
  OAI21_X1  g523(.A(KEYINPUT55), .B1(new_n724_), .B2(KEYINPUT116), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n722_), .A2(new_n723_), .A3(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n329_), .ZN(new_n727_));
  AOI21_X1  g526(.A(KEYINPUT117), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n330_), .B1(new_n728_), .B2(KEYINPUT56), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n309_), .B1(new_n728_), .B2(KEYINPUT56), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n719_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n711_), .B1(new_n732_), .B2(new_n254_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n726_), .A2(new_n727_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT117), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT56), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n308_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n738_), .A2(new_n729_), .ZN(new_n739_));
  OAI211_X1 g538(.A(KEYINPUT57), .B(new_n257_), .C1(new_n739_), .C2(new_n719_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n718_), .B1(KEYINPUT56), .B2(new_n734_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n726_), .A2(new_n737_), .A3(new_n727_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(new_n330_), .A3(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT58), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n741_), .A2(KEYINPUT58), .A3(new_n330_), .A4(new_n742_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n745_), .A2(new_n598_), .A3(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n733_), .A2(new_n740_), .A3(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(KEYINPUT115), .B1(new_n292_), .B2(new_n309_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n333_), .B2(new_n336_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n292_), .A2(KEYINPUT115), .A3(new_n309_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(new_n261_), .A3(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT54), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n752_), .A2(KEYINPUT54), .ZN(new_n754_));
  AOI22_X1  g553(.A1(new_n748_), .A2(new_n291_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n458_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n756_), .A2(new_n525_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(new_n555_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n755_), .A2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(G113gat), .B1(new_n759_), .B2(new_n308_), .ZN(new_n760_));
  OAI21_X1  g559(.A(KEYINPUT59), .B1(new_n755_), .B2(new_n758_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT120), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n758_), .A2(KEYINPUT119), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n748_), .A2(new_n291_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n754_), .A2(new_n753_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n764_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT59), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n768_), .B1(new_n758_), .B2(KEYINPUT119), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n763_), .B1(new_n767_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NOR4_X1   g571(.A1(new_n755_), .A2(KEYINPUT120), .A3(new_n769_), .A4(new_n764_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n762_), .B1(new_n772_), .B2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n308_), .A2(G113gat), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n776_), .B(KEYINPUT121), .Z(new_n777_));
  AOI21_X1  g576(.A(new_n760_), .B1(new_n775_), .B2(new_n777_), .ZN(G1340gat));
  OAI211_X1 g577(.A(new_n657_), .B(new_n761_), .C1(new_n771_), .C2(new_n773_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(G120gat), .ZN(new_n780_));
  INV_X1    g579(.A(G120gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n781_), .B1(new_n656_), .B2(KEYINPUT60), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n759_), .B(new_n782_), .C1(KEYINPUT60), .C2(new_n781_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n780_), .A2(new_n783_), .ZN(G1341gat));
  AOI21_X1  g583(.A(G127gat), .B1(new_n759_), .B2(new_n292_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n292_), .A2(G127gat), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT122), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n785_), .B1(new_n775_), .B2(new_n787_), .ZN(G1342gat));
  AOI21_X1  g587(.A(G134gat), .B1(new_n759_), .B2(new_n254_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n598_), .A2(G134gat), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n775_), .B2(new_n790_), .ZN(G1343gat));
  NOR3_X1   g590(.A1(new_n755_), .A2(new_n484_), .A3(new_n551_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n548_), .A2(new_n525_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(new_n308_), .A3(new_n793_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(KEYINPUT123), .B(G141gat), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n794_), .B(new_n795_), .ZN(G1344gat));
  NAND3_X1  g595(.A1(new_n792_), .A2(new_n657_), .A3(new_n793_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g597(.A1(new_n792_), .A2(new_n292_), .A3(new_n793_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(KEYINPUT61), .B(G155gat), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n799_), .B(new_n800_), .ZN(G1346gat));
  AND4_X1   g600(.A1(G162gat), .A2(new_n792_), .A3(new_n598_), .A4(new_n793_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n792_), .A2(new_n254_), .A3(new_n793_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n242_), .B2(new_n803_), .ZN(G1347gat));
  AOI21_X1  g603(.A(new_n526_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(new_n484_), .A3(new_n458_), .ZN(new_n806_));
  OAI21_X1  g605(.A(G169gat), .B1(new_n806_), .B2(new_n309_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT62), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NOR4_X1   g608(.A1(new_n755_), .A2(new_n555_), .A3(new_n526_), .A4(new_n756_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n810_), .B(new_n308_), .C1(new_n438_), .C2(new_n437_), .ZN(new_n811_));
  OAI211_X1 g610(.A(KEYINPUT62), .B(G169gat), .C1(new_n806_), .C2(new_n309_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n809_), .A2(new_n811_), .A3(new_n812_), .ZN(G1348gat));
  NAND4_X1  g612(.A1(new_n805_), .A2(new_n484_), .A3(new_n458_), .A4(new_n657_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n436_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT124), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT124), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n814_), .A2(new_n817_), .A3(new_n436_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT125), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n819_), .B1(new_n814_), .B2(new_n436_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n810_), .A2(KEYINPUT125), .A3(G176gat), .A4(new_n657_), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n816_), .A2(new_n818_), .B1(new_n820_), .B2(new_n821_), .ZN(G1349gat));
  NAND2_X1  g621(.A1(new_n810_), .A2(new_n292_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(G183gat), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n426_), .A2(new_n425_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n825_), .B2(new_n823_), .ZN(G1350gat));
  OAI21_X1  g625(.A(G190gat), .B1(new_n806_), .B2(new_n261_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n810_), .A2(new_n493_), .A3(new_n254_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(G1351gat));
  INV_X1    g628(.A(new_n549_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n830_), .A2(new_n551_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n805_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n308_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n657_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(G204gat), .ZN(G1353gat));
  XOR2_X1   g635(.A(KEYINPUT63), .B(G211gat), .Z(new_n837_));
  AND3_X1   g636(.A1(new_n832_), .A2(new_n292_), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n832_), .A2(new_n292_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n838_), .B1(new_n839_), .B2(new_n840_), .ZN(G1354gat));
  NAND3_X1  g640(.A1(new_n832_), .A2(KEYINPUT126), .A3(new_n254_), .ZN(new_n842_));
  XOR2_X1   g641(.A(KEYINPUT127), .B(G218gat), .Z(new_n843_));
  NAND3_X1  g642(.A1(new_n805_), .A2(new_n254_), .A3(new_n831_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT126), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n843_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n598_), .A2(new_n843_), .ZN(new_n847_));
  AOI22_X1  g646(.A1(new_n842_), .A2(new_n846_), .B1(new_n832_), .B2(new_n847_), .ZN(G1355gat));
endmodule


