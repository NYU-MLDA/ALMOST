//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 0 0 0 0 1 1 0 0 1 1 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n602_, new_n603_, new_n604_, new_n605_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n786_, new_n787_, new_n788_,
    new_n790_, new_n791_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n804_,
    new_n806_, new_n807_, new_n809_, new_n810_, new_n811_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n828_, new_n829_, new_n830_, new_n831_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n858_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G190gat), .B(G218gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT71), .ZN(new_n204_));
  INV_X1    g003(.A(G134gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G162gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT72), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G29gat), .B(G36gat), .ZN(new_n211_));
  INV_X1    g010(.A(G43gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G50gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT15), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n217_));
  XOR2_X1   g016(.A(G85gat), .B(G92gat), .Z(new_n218_));
  NOR2_X1   g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT7), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n219_), .B(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G99gat), .A2(G106gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT6), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n217_), .B(new_n218_), .C1(new_n221_), .C2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT8), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n224_), .B1(KEYINPUT9), .B2(new_n218_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G85gat), .A2(G92gat), .ZN(new_n228_));
  XOR2_X1   g027(.A(KEYINPUT10), .B(G99gat), .Z(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT64), .ZN(new_n230_));
  OAI221_X1 g029(.A(new_n227_), .B1(KEYINPUT9), .B2(new_n228_), .C1(new_n230_), .C2(G106gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n226_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n216_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT70), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G232gat), .A2(G233gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT34), .ZN(new_n237_));
  XOR2_X1   g036(.A(new_n237_), .B(KEYINPUT35), .Z(new_n238_));
  NAND3_X1  g037(.A1(new_n226_), .A2(new_n231_), .A3(new_n215_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n216_), .A2(KEYINPUT70), .A3(new_n232_), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n235_), .A2(new_n238_), .A3(new_n239_), .A4(new_n240_), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n235_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n237_), .A2(KEYINPUT35), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n210_), .B(new_n241_), .C1(new_n242_), .C2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n242_), .A2(KEYINPUT72), .A3(new_n238_), .ZN(new_n245_));
  AOI211_X1 g044(.A(KEYINPUT36), .B(new_n209_), .C1(new_n244_), .C2(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n209_), .A2(KEYINPUT36), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n209_), .A2(KEYINPUT36), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n244_), .A2(new_n248_), .A3(new_n249_), .A4(new_n245_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n202_), .B1(new_n246_), .B2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G230gat), .A2(G233gat), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G57gat), .B(G64gat), .ZN(new_n255_));
  AND2_X1   g054(.A1(new_n255_), .A2(KEYINPUT11), .ZN(new_n256_));
  XOR2_X1   g055(.A(G71gat), .B(G78gat), .Z(new_n257_));
  OR2_X1    g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n255_), .A2(KEYINPUT11), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n256_), .A2(new_n257_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n258_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n254_), .B1(new_n232_), .B2(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n263_), .B1(new_n262_), .B2(new_n232_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT66), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n232_), .A2(new_n265_), .A3(KEYINPUT12), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n266_), .B(new_n261_), .C1(KEYINPUT12), .C2(new_n232_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n232_), .A2(new_n265_), .A3(KEYINPUT12), .A4(new_n262_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n264_), .B1(new_n269_), .B2(new_n253_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G176gat), .B(G204gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(G148gat), .ZN(new_n272_));
  XOR2_X1   g071(.A(KEYINPUT67), .B(KEYINPUT5), .Z(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT68), .B(G120gat), .ZN(new_n275_));
  XOR2_X1   g074(.A(new_n274_), .B(new_n275_), .Z(new_n276_));
  XNOR2_X1  g075(.A(new_n270_), .B(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n278_));
  OR2_X1    g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n277_), .B1(KEYINPUT69), .B2(KEYINPUT13), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G127gat), .B(G155gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT16), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(G183gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(G211gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT17), .ZN(new_n286_));
  INV_X1    g085(.A(G211gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n284_), .B(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT17), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n286_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT73), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G231gat), .A2(G233gat), .ZN(new_n293_));
  XOR2_X1   g092(.A(new_n261_), .B(new_n293_), .Z(new_n294_));
  XNOR2_X1  g093(.A(G15gat), .B(G22gat), .ZN(new_n295_));
  INV_X1    g094(.A(G1gat), .ZN(new_n296_));
  INV_X1    g095(.A(G8gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT14), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n295_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G1gat), .B(G8gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n294_), .B(new_n301_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n292_), .B(new_n302_), .C1(new_n265_), .C2(new_n286_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n286_), .A2(KEYINPUT66), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT74), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT74), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n303_), .A2(new_n308_), .A3(new_n305_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n244_), .A2(new_n249_), .A3(new_n245_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n247_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n312_), .A2(KEYINPUT37), .A3(new_n250_), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n252_), .A2(new_n281_), .A3(new_n310_), .A4(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT75), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G57gat), .B(G85gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G1gat), .B(G29gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT91), .B(KEYINPUT0), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G225gat), .A2(G233gat), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT83), .ZN(new_n324_));
  INV_X1    g123(.A(G155gat), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n324_), .A2(new_n325_), .A3(new_n207_), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT83), .B1(G155gat), .B2(G162gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G155gat), .A2(G162gat), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n326_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT84), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G141gat), .A2(G148gat), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT2), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n330_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n332_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(KEYINPUT84), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n333_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  OR3_X1    g135(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n329_), .B1(new_n336_), .B2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n328_), .A2(KEYINPUT1), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT1), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(G155gat), .A3(G162gat), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n326_), .A2(new_n341_), .A3(new_n343_), .A4(new_n327_), .ZN(new_n344_));
  OR2_X1    g143(.A1(G141gat), .A2(G148gat), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n344_), .A2(new_n331_), .A3(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n340_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(G120gat), .ZN(new_n348_));
  INV_X1    g147(.A(G127gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(new_n205_), .ZN(new_n350_));
  INV_X1    g149(.A(G113gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G127gat), .A2(G134gat), .ZN(new_n352_));
  AND3_X1   g151(.A1(new_n350_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n351_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n348_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n350_), .A2(new_n352_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(G113gat), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n350_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n357_), .A2(G120gat), .A3(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n355_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n347_), .A2(new_n360_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n340_), .A2(new_n355_), .A3(new_n359_), .A4(new_n346_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n361_), .A2(KEYINPUT4), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT4), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n347_), .A2(new_n360_), .A3(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n323_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n323_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n367_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n322_), .B1(new_n366_), .B2(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT33), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G226gat), .A2(G233gat), .ZN(new_n371_));
  XOR2_X1   g170(.A(new_n371_), .B(KEYINPUT88), .Z(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT19), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G211gat), .B(G218gat), .ZN(new_n375_));
  XOR2_X1   g174(.A(G197gat), .B(G204gat), .Z(new_n376_));
  OAI21_X1  g175(.A(new_n375_), .B1(new_n376_), .B2(KEYINPUT21), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(KEYINPUT21), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(G169gat), .A2(G176gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(KEYINPUT76), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G169gat), .A2(G176gat), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n381_), .A2(KEYINPUT24), .A3(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT25), .B(G183gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT26), .B(G190gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n383_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G183gat), .A2(G190gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AND2_X1   g189(.A1(KEYINPUT78), .A2(KEYINPUT23), .ZN(new_n391_));
  NOR2_X1   g190(.A1(KEYINPUT78), .A2(KEYINPUT23), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n390_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT81), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n389_), .A2(KEYINPUT23), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT80), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n389_), .A2(KEYINPUT80), .A3(KEYINPUT23), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  OAI211_X1 g199(.A(KEYINPUT81), .B(new_n390_), .C1(new_n391_), .C2(new_n392_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n395_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT89), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT76), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n380_), .B(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT24), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n402_), .A2(new_n403_), .A3(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n403_), .B1(new_n402_), .B2(new_n407_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n388_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n391_), .A2(new_n392_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(new_n389_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n389_), .A2(KEYINPUT23), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(G183gat), .A2(G190gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT79), .B(G176gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT22), .B(G169gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n382_), .B(KEYINPUT77), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n417_), .A2(KEYINPUT90), .A3(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT90), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n415_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n425_), .B1(new_n426_), .B2(new_n422_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n424_), .A2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n379_), .B1(new_n410_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n402_), .A2(new_n416_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n423_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n381_), .A2(new_n421_), .A3(KEYINPUT24), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n432_), .A2(new_n407_), .A3(new_n386_), .A4(new_n414_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n379_), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT20), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n374_), .B1(new_n429_), .B2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G8gat), .B(G36gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT18), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(G64gat), .ZN(new_n440_));
  INV_X1    g239(.A(G92gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n410_), .A2(new_n379_), .A3(new_n428_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT20), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n444_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n443_), .A2(new_n445_), .A3(new_n373_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n437_), .A2(new_n442_), .A3(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n363_), .A2(new_n365_), .ZN(new_n448_));
  OR3_X1    g247(.A1(new_n448_), .A2(KEYINPUT93), .A3(new_n367_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT92), .ZN(new_n450_));
  INV_X1    g249(.A(new_n361_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n362_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n450_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n361_), .A2(KEYINPUT92), .A3(new_n362_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n453_), .A2(new_n367_), .A3(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT93), .B1(new_n448_), .B2(new_n367_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n449_), .A2(new_n321_), .A3(new_n455_), .A4(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n442_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n402_), .A2(new_n407_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT89), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n402_), .A2(new_n403_), .A3(new_n407_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n387_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n428_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n435_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n432_), .A2(new_n386_), .A3(new_n414_), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n465_), .A2(new_n407_), .B1(new_n430_), .B2(new_n423_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n444_), .B1(new_n466_), .B2(new_n379_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n373_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n443_), .A2(new_n445_), .A3(new_n373_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n458_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n370_), .A2(new_n447_), .A3(new_n457_), .A4(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n442_), .A2(KEYINPUT32), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n437_), .A2(new_n446_), .A3(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n448_), .A2(new_n367_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n368_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(new_n321_), .A3(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(new_n369_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n473_), .A2(new_n477_), .ZN(new_n478_));
  OR2_X1    g277(.A1(new_n426_), .A2(new_n422_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n410_), .A2(new_n379_), .A3(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n445_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(new_n374_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n464_), .A2(new_n467_), .A3(new_n373_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n472_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT94), .B1(new_n478_), .B2(new_n484_), .ZN(new_n485_));
  NOR3_X1   g284(.A1(new_n429_), .A2(new_n436_), .A3(new_n374_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n373_), .B1(new_n480_), .B2(new_n445_), .ZN(new_n487_));
  OAI211_X1 g286(.A(KEYINPUT32), .B(new_n442_), .C1(new_n486_), .C2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT94), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n488_), .A2(new_n489_), .A3(new_n477_), .A4(new_n473_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n471_), .A2(new_n485_), .A3(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n379_), .B1(KEYINPUT29), .B2(new_n347_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G22gat), .B(G50gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(G78gat), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n492_), .A2(new_n494_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G228gat), .A2(G233gat), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT86), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n498_), .B1(new_n379_), .B2(new_n499_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n500_), .A2(G106gat), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(G106gat), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n497_), .A2(new_n503_), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n495_), .B(new_n496_), .C1(new_n501_), .C2(new_n502_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n347_), .A2(KEYINPUT29), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n507_), .A2(KEYINPUT87), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(KEYINPUT87), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AND3_X1   g310(.A1(new_n508_), .A2(new_n509_), .A3(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n511_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n506_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n514_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n491_), .A2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n458_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n521_), .A2(KEYINPUT27), .A3(new_n447_), .ZN(new_n522_));
  AOI21_X1  g321(.A(KEYINPUT27), .B1(new_n470_), .B2(new_n447_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n477_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n520_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT95), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n466_), .B(KEYINPUT30), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(new_n360_), .ZN(new_n530_));
  XOR2_X1   g329(.A(KEYINPUT82), .B(KEYINPUT31), .Z(new_n531_));
  NAND2_X1  g330(.A1(G227gat), .A2(G233gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G71gat), .B(G99gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G15gat), .B(G43gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n533_), .B(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n530_), .B(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n527_), .A2(new_n528_), .A3(new_n538_), .ZN(new_n539_));
  AOI22_X1  g338(.A1(new_n491_), .A2(new_n519_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n538_), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT95), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT96), .ZN(new_n543_));
  INV_X1    g342(.A(new_n523_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n521_), .A2(KEYINPUT27), .A3(new_n447_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n543_), .B1(new_n546_), .B2(new_n518_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n477_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n519_), .A2(new_n524_), .A3(KEYINPUT96), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n547_), .A2(new_n548_), .A3(new_n549_), .A4(new_n541_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n539_), .A2(new_n542_), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n215_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n552_), .A2(new_n301_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n553_), .B1(new_n216_), .B2(new_n301_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G229gat), .A2(G233gat), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n215_), .B(new_n301_), .Z(new_n557_));
  NAND3_X1  g356(.A1(new_n557_), .A2(G229gat), .A3(G233gat), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(G113gat), .B(G141gat), .Z(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(G169gat), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n561_), .B(G197gat), .Z(new_n562_));
  OR2_X1    g361(.A1(new_n559_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n559_), .A2(new_n562_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n316_), .A2(new_n551_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT97), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n548_), .A2(G1gat), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT99), .ZN(new_n570_));
  XOR2_X1   g369(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n571_));
  OAI211_X1 g370(.A(new_n568_), .B(new_n569_), .C1(new_n570_), .C2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n570_), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT100), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n575_), .B1(new_n246_), .B2(new_n251_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n312_), .A2(KEYINPUT100), .A3(new_n250_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n551_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n281_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n565_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n579_), .A2(new_n306_), .A3(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(G1gat), .B1(new_n583_), .B2(new_n548_), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n584_), .B(KEYINPUT101), .Z(new_n585_));
  NAND2_X1  g384(.A1(new_n572_), .A2(new_n573_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n574_), .A2(new_n585_), .A3(new_n586_), .ZN(G1324gat));
  NAND3_X1  g386(.A1(new_n568_), .A2(new_n297_), .A3(new_n546_), .ZN(new_n588_));
  OAI21_X1  g387(.A(G8gat), .B1(new_n583_), .B2(new_n524_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT39), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT40), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(G1325gat));
  OAI21_X1  g392(.A(G15gat), .B1(new_n583_), .B2(new_n538_), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT41), .Z(new_n595_));
  INV_X1    g394(.A(G15gat), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n568_), .A2(new_n596_), .A3(new_n541_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT102), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n597_), .A2(new_n598_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n595_), .B1(new_n599_), .B2(new_n600_), .ZN(G1326gat));
  INV_X1    g400(.A(G22gat), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n568_), .A2(new_n602_), .A3(new_n518_), .ZN(new_n603_));
  OAI21_X1  g402(.A(G22gat), .B1(new_n583_), .B2(new_n519_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT42), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n605_), .ZN(G1327gat));
  OR3_X1    g405(.A1(new_n578_), .A2(KEYINPUT106), .A3(new_n310_), .ZN(new_n607_));
  OAI21_X1  g406(.A(KEYINPUT106), .B1(new_n578_), .B2(new_n310_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n609_), .A2(new_n551_), .A3(new_n582_), .ZN(new_n610_));
  OR3_X1    g409(.A1(new_n610_), .A2(G29gat), .A3(new_n548_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n252_), .A2(new_n313_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n551_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(KEYINPUT43), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT103), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n613_), .A2(KEYINPUT43), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n613_), .A2(KEYINPUT103), .A3(KEYINPUT43), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n616_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n310_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(new_n582_), .A3(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT104), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n624_), .A2(KEYINPUT44), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n619_), .A2(new_n582_), .A3(new_n620_), .A4(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n623_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n477_), .ZN(new_n628_));
  AOI21_X1  g427(.A(KEYINPUT105), .B1(new_n628_), .B2(G29gat), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT105), .ZN(new_n630_));
  INV_X1    g429(.A(G29gat), .ZN(new_n631_));
  AOI211_X1 g430(.A(new_n630_), .B(new_n631_), .C1(new_n627_), .C2(new_n477_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n611_), .B1(new_n629_), .B2(new_n632_), .ZN(G1328gat));
  XNOR2_X1  g432(.A(new_n546_), .B(KEYINPUT107), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n610_), .A2(G36gat), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT45), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n524_), .B1(new_n623_), .B2(new_n626_), .ZN(new_n639_));
  INV_X1    g438(.A(G36gat), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n638_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT46), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n638_), .B(KEYINPUT46), .C1(new_n639_), .C2(new_n640_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(G1329gat));
  OR3_X1    g444(.A1(new_n610_), .A2(G43gat), .A3(new_n538_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n538_), .B1(new_n623_), .B2(new_n626_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n646_), .B1(new_n647_), .B2(new_n212_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n649_), .B(new_n646_), .C1(new_n647_), .C2(new_n212_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(G1330gat));
  AOI21_X1  g452(.A(new_n519_), .B1(new_n623_), .B2(new_n626_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n518_), .A2(new_n214_), .ZN(new_n655_));
  OAI22_X1  g454(.A1(new_n654_), .A2(new_n214_), .B1(new_n610_), .B2(new_n655_), .ZN(G1331gat));
  NOR2_X1   g455(.A1(new_n281_), .A2(new_n565_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n551_), .A2(new_n657_), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n252_), .A2(new_n310_), .A3(new_n313_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(G57gat), .B1(new_n661_), .B2(new_n477_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n579_), .A2(new_n310_), .A3(new_n657_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT109), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n663_), .B(new_n664_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n477_), .A2(G57gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n662_), .B1(new_n665_), .B2(new_n666_), .ZN(G1332gat));
  INV_X1    g466(.A(G64gat), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n661_), .A2(new_n668_), .A3(new_n634_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n663_), .B(KEYINPUT109), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n670_), .A2(new_n635_), .ZN(new_n671_));
  OAI21_X1  g470(.A(KEYINPUT110), .B1(new_n671_), .B2(new_n668_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT110), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n673_), .B(G64gat), .C1(new_n670_), .C2(new_n635_), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n672_), .A2(KEYINPUT48), .A3(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(KEYINPUT48), .B1(new_n672_), .B2(new_n674_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n669_), .B1(new_n675_), .B2(new_n676_), .ZN(G1333gat));
  OAI21_X1  g476(.A(G71gat), .B1(new_n670_), .B2(new_n538_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT49), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n538_), .A2(G71gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n679_), .B1(new_n660_), .B2(new_n680_), .ZN(G1334gat));
  OAI21_X1  g480(.A(G78gat), .B1(new_n670_), .B2(new_n519_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT50), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n519_), .A2(G78gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n683_), .B1(new_n660_), .B2(new_n684_), .ZN(G1335gat));
  AND2_X1   g484(.A1(new_n609_), .A2(new_n658_), .ZN(new_n686_));
  AOI21_X1  g485(.A(G85gat), .B1(new_n686_), .B2(new_n477_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT111), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n619_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(new_n657_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n620_), .B1(new_n619_), .B2(new_n688_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n477_), .A2(G85gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n687_), .B1(new_n692_), .B2(new_n693_), .ZN(G1336gat));
  AOI21_X1  g493(.A(G92gat), .B1(new_n686_), .B2(new_n546_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n635_), .A2(new_n441_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n692_), .B2(new_n696_), .ZN(G1337gat));
  NOR2_X1   g496(.A1(new_n538_), .A2(new_n230_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n686_), .A2(new_n698_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n690_), .A2(new_n691_), .A3(new_n538_), .ZN(new_n700_));
  INV_X1    g499(.A(G99gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n699_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT51), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n703_), .A2(KEYINPUT112), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  OAI221_X1 g504(.A(new_n699_), .B1(KEYINPUT112), .B2(new_n703_), .C1(new_n700_), .C2(new_n701_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1338gat));
  NOR3_X1   g506(.A1(new_n281_), .A2(new_n519_), .A3(new_n565_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n619_), .A2(new_n620_), .A3(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n709_), .A2(G106gat), .A3(new_n710_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(G106gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n686_), .A2(new_n714_), .A3(new_n518_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n712_), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n709_), .A2(G106gat), .A3(new_n710_), .A4(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n713_), .A2(new_n715_), .A3(new_n717_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n713_), .A2(new_n719_), .A3(new_n715_), .A4(new_n717_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1339gat));
  XNOR2_X1  g522(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n659_), .A2(new_n581_), .A3(new_n281_), .A4(new_n725_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n724_), .B1(new_n314_), .B2(new_n565_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n267_), .A2(new_n268_), .A3(new_n254_), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT116), .Z(new_n731_));
  AND3_X1   g530(.A1(new_n269_), .A2(KEYINPUT55), .A3(new_n253_), .ZN(new_n732_));
  AOI21_X1  g531(.A(KEYINPUT55), .B1(new_n269_), .B2(new_n253_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n731_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n276_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT56), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT117), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n730_), .B(KEYINPUT116), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n740_), .A2(new_n733_), .A3(new_n732_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n739_), .B1(new_n741_), .B2(new_n276_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT56), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n735_), .A2(KEYINPUT117), .A3(new_n743_), .A4(new_n736_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n581_), .B1(new_n270_), .B2(new_n276_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n738_), .A2(new_n742_), .A3(new_n744_), .A4(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n557_), .A2(new_n555_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n554_), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n562_), .B(new_n747_), .C1(new_n748_), .C2(new_n555_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n277_), .A2(new_n563_), .A3(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n746_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(new_n578_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT57), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n741_), .A2(new_n276_), .ZN(new_n755_));
  AOI22_X1  g554(.A1(new_n755_), .A2(new_n743_), .B1(new_n270_), .B2(new_n276_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n563_), .A2(new_n749_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n757_), .B1(new_n737_), .B2(KEYINPUT56), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT118), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n760_), .A2(KEYINPUT58), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n756_), .B(new_n758_), .C1(new_n760_), .C2(KEYINPUT58), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n762_), .A2(new_n763_), .A3(new_n612_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n751_), .A2(KEYINPUT57), .A3(new_n578_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n754_), .A2(new_n764_), .A3(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n306_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n729_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n547_), .A2(new_n477_), .A3(new_n549_), .A4(new_n541_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(G113gat), .B1(new_n770_), .B2(new_n565_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT59), .ZN(new_n772_));
  XOR2_X1   g571(.A(new_n769_), .B(KEYINPUT119), .Z(new_n773_));
  AND3_X1   g572(.A1(new_n751_), .A2(KEYINPUT57), .A3(new_n578_), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT57), .B1(new_n751_), .B2(new_n578_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n310_), .B1(new_n776_), .B2(new_n764_), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n772_), .B(new_n773_), .C1(new_n777_), .C2(new_n729_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT59), .B1(new_n768_), .B2(new_n769_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT120), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n778_), .A2(new_n779_), .A3(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n581_), .A2(new_n351_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n771_), .B1(new_n783_), .B2(new_n784_), .ZN(G1340gat));
  OAI21_X1  g584(.A(new_n348_), .B1(new_n281_), .B2(KEYINPUT60), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n770_), .B(new_n786_), .C1(KEYINPUT60), .C2(new_n348_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n778_), .A2(new_n779_), .A3(new_n580_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n787_), .B1(new_n788_), .B2(new_n348_), .ZN(G1341gat));
  AOI21_X1  g588(.A(G127gat), .B1(new_n770_), .B2(new_n310_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n767_), .A2(new_n349_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n783_), .B2(new_n791_), .ZN(G1342gat));
  INV_X1    g591(.A(new_n578_), .ZN(new_n793_));
  AOI21_X1  g592(.A(G134gat), .B1(new_n770_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n612_), .A2(G134gat), .ZN(new_n795_));
  XOR2_X1   g594(.A(new_n795_), .B(KEYINPUT121), .Z(new_n796_));
  AOI21_X1  g595(.A(new_n794_), .B1(new_n783_), .B2(new_n796_), .ZN(G1343gat));
  NOR2_X1   g596(.A1(new_n541_), .A2(new_n519_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n635_), .A2(new_n477_), .A3(new_n798_), .ZN(new_n799_));
  XOR2_X1   g598(.A(new_n799_), .B(KEYINPUT122), .Z(new_n800_));
  NOR2_X1   g599(.A1(new_n768_), .A2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n565_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n580_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g604(.A1(new_n801_), .A2(new_n310_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(KEYINPUT61), .B(G155gat), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n806_), .B(new_n807_), .ZN(G1346gat));
  AOI21_X1  g607(.A(G162gat), .B1(new_n801_), .B2(new_n793_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n612_), .A2(G162gat), .ZN(new_n810_));
  XOR2_X1   g609(.A(new_n810_), .B(KEYINPUT123), .Z(new_n811_));
  AOI21_X1  g610(.A(new_n809_), .B1(new_n801_), .B2(new_n811_), .ZN(G1347gat));
  NOR2_X1   g611(.A1(new_n635_), .A2(new_n477_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n813_), .A2(new_n541_), .A3(new_n519_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n565_), .B(new_n815_), .C1(new_n777_), .C2(new_n729_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT124), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n766_), .A2(new_n620_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n814_), .B1(new_n818_), .B2(new_n728_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT124), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n820_), .A3(new_n565_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n817_), .A2(G169gat), .A3(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT62), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n819_), .A2(new_n419_), .A3(new_n565_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n817_), .A2(new_n821_), .A3(KEYINPUT62), .A4(G169gat), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n824_), .A2(new_n825_), .A3(new_n826_), .ZN(G1348gat));
  NAND2_X1  g626(.A1(new_n766_), .A2(new_n767_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n728_), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n829_), .A2(G176gat), .A3(new_n580_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n819_), .A2(new_n580_), .ZN(new_n831_));
  AOI22_X1  g630(.A1(new_n830_), .A2(new_n815_), .B1(new_n831_), .B2(new_n418_), .ZN(G1349gat));
  INV_X1    g631(.A(new_n384_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n819_), .A2(new_n306_), .A3(new_n833_), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n768_), .A2(new_n620_), .A3(new_n814_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(G183gat), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT125), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n836_), .B(new_n837_), .ZN(G1350gat));
  NAND2_X1  g637(.A1(new_n793_), .A2(new_n385_), .ZN(new_n839_));
  XOR2_X1   g638(.A(new_n839_), .B(KEYINPUT126), .Z(new_n840_));
  NAND2_X1  g639(.A1(new_n819_), .A2(new_n840_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n819_), .A2(new_n612_), .ZN(new_n842_));
  INV_X1    g641(.A(G190gat), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n841_), .B1(new_n842_), .B2(new_n843_), .ZN(G1351gat));
  AND3_X1   g643(.A1(new_n829_), .A2(new_n798_), .A3(new_n813_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n565_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n580_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT127), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(G204gat), .ZN(new_n850_));
  XNOR2_X1  g649(.A(KEYINPUT127), .B(G204gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n848_), .B2(new_n851_), .ZN(G1353gat));
  NAND2_X1  g651(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n845_), .A2(new_n306_), .A3(new_n853_), .ZN(new_n854_));
  OR2_X1    g653(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n854_), .B(new_n855_), .ZN(G1354gat));
  AOI21_X1  g655(.A(G218gat), .B1(new_n845_), .B2(new_n793_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n612_), .A2(G218gat), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n857_), .B1(new_n845_), .B2(new_n858_), .ZN(G1355gat));
endmodule


