//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 1 0 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 0 1 0 0 1 1 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n924_, new_n926_, new_n928_, new_n929_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n957_, new_n958_, new_n959_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n968_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_;
  INV_X1    g000(.A(KEYINPUT12), .ZN(new_n202_));
  XOR2_X1   g001(.A(G71gat), .B(G78gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(G57gat), .B(G64gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(new_n203_), .B1(KEYINPUT11), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT65), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT65), .ZN(new_n207_));
  OAI211_X1 g006(.A(new_n203_), .B(new_n207_), .C1(KEYINPUT11), .C2(new_n204_), .ZN(new_n208_));
  AND2_X1   g007(.A1(new_n204_), .A2(KEYINPUT11), .ZN(new_n209_));
  AND3_X1   g008(.A1(new_n206_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n209_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n202_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT6), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT6), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(G99gat), .A3(G106gat), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT64), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n216_), .A2(new_n218_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G99gat), .A2(G106gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT7), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n220_), .A2(new_n223_), .A3(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(G85gat), .B(G92gat), .Z(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n228_), .A2(KEYINPUT8), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT7), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n224_), .B(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n227_), .B1(new_n231_), .B2(new_n219_), .ZN(new_n232_));
  AOI22_X1  g031(.A1(new_n226_), .A2(new_n229_), .B1(new_n232_), .B2(KEYINPUT8), .ZN(new_n233_));
  XOR2_X1   g032(.A(KEYINPUT10), .B(G99gat), .Z(new_n234_));
  INV_X1    g033(.A(G106gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n227_), .A2(KEYINPUT9), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G85gat), .A2(G92gat), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n236_), .B(new_n237_), .C1(KEYINPUT9), .C2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n220_), .A2(new_n223_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n233_), .A2(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n210_), .A2(new_n211_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n214_), .B1(new_n213_), .B2(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n202_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n242_), .A2(new_n243_), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G230gat), .A2(G233gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n245_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n249_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n247_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n251_), .B1(new_n252_), .B2(new_n244_), .ZN(new_n253_));
  XOR2_X1   g052(.A(G120gat), .B(G148gat), .Z(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G176gat), .B(G204gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n250_), .A2(new_n253_), .A3(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n250_), .A2(KEYINPUT68), .A3(new_n253_), .A4(new_n259_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n250_), .A2(new_n253_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(new_n258_), .ZN(new_n266_));
  AND2_X1   g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  XOR2_X1   g066(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n264_), .A2(new_n266_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n270_), .B1(KEYINPUT69), .B2(KEYINPUT13), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n239_), .A2(new_n240_), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n226_), .A2(new_n229_), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n232_), .A2(KEYINPUT8), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n273_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G29gat), .B(G36gat), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  XOR2_X1   g077(.A(G43gat), .B(G50gat), .Z(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G43gat), .B(G50gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n277_), .A2(new_n281_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT70), .B(KEYINPUT15), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n276_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n283_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n242_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G232gat), .A2(G233gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT34), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n290_), .A2(KEYINPUT35), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n286_), .A2(new_n288_), .A3(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(KEYINPUT35), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G190gat), .B(G218gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G134gat), .B(G162gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n298_), .A2(KEYINPUT36), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n286_), .A2(new_n288_), .A3(new_n293_), .A4(new_n291_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n295_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT71), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n295_), .A2(KEYINPUT71), .A3(new_n299_), .A4(new_n300_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n295_), .A2(new_n300_), .ZN(new_n305_));
  XOR2_X1   g104(.A(new_n298_), .B(KEYINPUT36), .Z(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT72), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  AOI22_X1  g107(.A1(new_n303_), .A2(new_n304_), .B1(new_n305_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT73), .ZN(new_n310_));
  AND3_X1   g109(.A1(new_n309_), .A2(new_n310_), .A3(KEYINPUT37), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n310_), .A2(KEYINPUT37), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(KEYINPUT37), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NOR3_X1   g113(.A1(new_n309_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n311_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G231gat), .A2(G233gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n243_), .B(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT74), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G15gat), .B(G22gat), .ZN(new_n320_));
  INV_X1    g119(.A(G1gat), .ZN(new_n321_));
  INV_X1    g120(.A(G8gat), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT14), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n320_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G1gat), .B(G8gat), .ZN(new_n325_));
  XOR2_X1   g124(.A(new_n324_), .B(new_n325_), .Z(new_n326_));
  XNOR2_X1  g125(.A(new_n319_), .B(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G127gat), .B(G155gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT16), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G183gat), .B(G211gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT76), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n334_), .A2(KEYINPUT66), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n327_), .A2(new_n335_), .ZN(new_n336_));
  XOR2_X1   g135(.A(new_n331_), .B(KEYINPUT17), .Z(new_n337_));
  AOI21_X1  g136(.A(new_n337_), .B1(new_n334_), .B2(new_n213_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n327_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n336_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n316_), .A2(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n272_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n324_), .B(new_n325_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n285_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n326_), .A2(new_n287_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G229gat), .A2(G233gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n346_), .B(KEYINPUT78), .Z(new_n347_));
  NAND3_X1  g146(.A1(new_n344_), .A2(new_n345_), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n343_), .A2(new_n283_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n345_), .A2(KEYINPUT77), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT77), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n343_), .A2(new_n351_), .A3(new_n283_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n350_), .A2(G229gat), .A3(G233gat), .A4(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G113gat), .B(G141gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT79), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G169gat), .B(G197gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n348_), .A2(new_n353_), .A3(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT80), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT80), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n348_), .A2(new_n353_), .A3(new_n360_), .A4(new_n357_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n348_), .A2(new_n353_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n357_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n362_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT81), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT81), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n362_), .A2(new_n368_), .A3(new_n365_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G183gat), .A2(G190gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT23), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT23), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n374_), .A2(G183gat), .A3(G190gat), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT24), .ZN(new_n376_));
  NOR2_X1   g175(.A1(G169gat), .A2(G176gat), .ZN(new_n377_));
  AOI22_X1  g176(.A1(new_n373_), .A2(new_n375_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(G183gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT25), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT25), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(G183gat), .ZN(new_n382_));
  INV_X1    g181(.A(G190gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT26), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT26), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(G190gat), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n380_), .A2(new_n382_), .A3(new_n384_), .A4(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G169gat), .A2(G176gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n378_), .A2(new_n387_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT82), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n372_), .A2(new_n374_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n379_), .A2(new_n383_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n398_));
  OR3_X1    g197(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n392_), .A2(new_n393_), .A3(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n393_), .B1(new_n392_), .B2(new_n400_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT83), .B(KEYINPUT30), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n392_), .A2(new_n400_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT82), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n392_), .A2(new_n393_), .A3(new_n400_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n404_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n405_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT86), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT86), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n405_), .A2(new_n411_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G15gat), .B(G43gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT84), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G227gat), .A2(G233gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT85), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n418_), .B(new_n420_), .ZN(new_n421_));
  XOR2_X1   g220(.A(G71gat), .B(G99gat), .Z(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n416_), .A2(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n423_), .B1(new_n412_), .B2(KEYINPUT86), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(G134gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(G127gat), .ZN(new_n428_));
  INV_X1    g227(.A(G127gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(G134gat), .ZN(new_n430_));
  INV_X1    g229(.A(G120gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(G113gat), .ZN(new_n432_));
  INV_X1    g231(.A(G113gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(G120gat), .ZN(new_n434_));
  AND4_X1   g233(.A1(new_n428_), .A2(new_n430_), .A3(new_n432_), .A4(new_n434_), .ZN(new_n435_));
  AOI22_X1  g234(.A1(new_n428_), .A2(new_n430_), .B1(new_n432_), .B2(new_n434_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT31), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n424_), .A2(new_n426_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n438_), .ZN(new_n440_));
  XOR2_X1   g239(.A(new_n421_), .B(new_n422_), .Z(new_n441_));
  AOI21_X1  g240(.A(new_n441_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n440_), .B1(new_n442_), .B2(new_n425_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n439_), .A2(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(G155gat), .A2(G162gat), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G155gat), .A2(G162gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NOR3_X1   g249(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n448_), .B1(new_n452_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n447_), .ZN(new_n458_));
  NOR3_X1   g257(.A1(new_n458_), .A2(new_n445_), .A3(KEYINPUT1), .ZN(new_n459_));
  INV_X1    g258(.A(G141gat), .ZN(new_n460_));
  INV_X1    g259(.A(G148gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G141gat), .A2(G148gat), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT1), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n462_), .B(new_n463_), .C1(new_n464_), .C2(new_n447_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n459_), .A2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n437_), .B1(new_n457_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT3), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT2), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n463_), .A2(new_n470_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n469_), .A2(new_n471_), .A3(new_n453_), .A4(new_n449_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n472_), .A2(new_n447_), .A3(new_n446_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n428_), .A2(new_n430_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n432_), .A2(new_n434_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n428_), .A2(new_n430_), .A3(new_n432_), .A4(new_n434_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n446_), .A2(new_n464_), .A3(new_n447_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n458_), .A2(KEYINPUT1), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n479_), .A2(new_n480_), .A3(new_n463_), .A4(new_n462_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n473_), .A2(new_n478_), .A3(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n467_), .A2(KEYINPUT4), .A3(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT97), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n467_), .A2(KEYINPUT97), .A3(new_n482_), .A4(KEYINPUT4), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G225gat), .A2(G233gat), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n489_), .B1(new_n467_), .B2(KEYINPUT4), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n487_), .A2(new_n491_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n467_), .A2(new_n482_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n488_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G1gat), .B(G29gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(G85gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT0), .B(G57gat), .ZN(new_n497_));
  XOR2_X1   g296(.A(new_n496_), .B(new_n497_), .Z(new_n498_));
  NAND3_X1  g297(.A1(new_n492_), .A2(new_n494_), .A3(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT98), .ZN(new_n500_));
  INV_X1    g299(.A(new_n498_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n490_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n494_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n501_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n499_), .A2(new_n500_), .A3(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n500_), .B1(new_n499_), .B2(new_n504_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n444_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n473_), .A2(new_n481_), .ZN(new_n509_));
  OR3_X1    g308(.A1(new_n509_), .A2(KEYINPUT87), .A3(KEYINPUT29), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT87), .B1(new_n509_), .B2(KEYINPUT29), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G22gat), .B(G50gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT28), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n510_), .A2(new_n511_), .A3(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n513_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G78gat), .B(G106gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT93), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT89), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT88), .ZN(new_n520_));
  INV_X1    g319(.A(G204gat), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n520_), .B1(new_n521_), .B2(G197gat), .ZN(new_n522_));
  INV_X1    g321(.A(G197gat), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n523_), .A2(G204gat), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(KEYINPUT88), .A3(G204gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT21), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n519_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G211gat), .B(G218gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n523_), .A2(G204gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n521_), .A2(G197gat), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n531_), .A3(new_n520_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n532_), .A2(KEYINPUT89), .A3(KEYINPUT21), .A4(new_n526_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT90), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n534_), .B1(new_n521_), .B2(G197gat), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n523_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT21), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .A4(new_n531_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n528_), .A2(new_n529_), .A3(new_n533_), .A4(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n535_), .A2(new_n536_), .A3(new_n531_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT91), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT91), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n535_), .A2(new_n536_), .A3(new_n542_), .A4(new_n531_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n529_), .A2(new_n537_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n541_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n539_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT92), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n509_), .A2(KEYINPUT29), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G228gat), .A2(G233gat), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n547_), .A2(new_n549_), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT29), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n553_), .B1(new_n473_), .B2(new_n481_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n554_), .B1(new_n539_), .B2(new_n545_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT92), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n556_), .B1(new_n539_), .B2(new_n545_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n555_), .B1(new_n557_), .B2(new_n550_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n518_), .B1(new_n552_), .B2(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n516_), .B1(new_n559_), .B2(KEYINPUT94), .ZN(new_n560_));
  INV_X1    g359(.A(new_n518_), .ZN(new_n561_));
  NOR3_X1   g360(.A1(new_n555_), .A2(new_n557_), .A3(new_n550_), .ZN(new_n562_));
  AOI221_X4 g361(.A(new_n554_), .B1(new_n556_), .B2(new_n551_), .C1(new_n545_), .C2(new_n539_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n561_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n552_), .A2(new_n558_), .A3(new_n518_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n560_), .A2(new_n566_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n564_), .A2(new_n516_), .A3(KEYINPUT94), .A4(new_n565_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT99), .B(KEYINPUT27), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT20), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n571_), .B1(new_n409_), .B2(new_n546_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G226gat), .A2(G233gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT19), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT25), .B(G183gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT26), .B(G190gat), .ZN(new_n577_));
  AOI22_X1  g376(.A1(new_n576_), .A2(new_n577_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n399_), .A2(new_n398_), .ZN(new_n579_));
  AOI22_X1  g378(.A1(new_n578_), .A2(new_n378_), .B1(new_n579_), .B2(new_n397_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n539_), .A2(new_n580_), .A3(new_n545_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT95), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n539_), .A2(new_n580_), .A3(new_n545_), .A4(KEYINPUT95), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n572_), .A2(new_n575_), .A3(new_n583_), .A4(new_n584_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n407_), .A2(new_n408_), .A3(new_n545_), .A4(new_n539_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n546_), .A2(new_n406_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n586_), .A2(new_n587_), .A3(KEYINPUT20), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(new_n574_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G8gat), .B(G36gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G64gat), .B(G92gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n585_), .A2(new_n589_), .A3(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n595_), .B1(new_n585_), .B2(new_n589_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n570_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n588_), .A2(new_n574_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n575_), .B1(new_n572_), .B2(new_n581_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n594_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n585_), .A2(new_n589_), .A3(new_n595_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n601_), .A2(KEYINPUT27), .A3(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n598_), .A2(new_n603_), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n508_), .A2(new_n569_), .A3(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n595_), .A2(KEYINPUT32), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n607_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n585_), .A2(new_n589_), .A3(new_n606_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n498_), .B1(new_n492_), .B2(new_n494_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n502_), .A2(new_n503_), .A3(new_n501_), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n608_), .B(new_n609_), .C1(new_n610_), .C2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT33), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n499_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(KEYINPUT33), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n539_), .A2(new_n545_), .ZN(new_n617_));
  OAI211_X1 g416(.A(KEYINPUT20), .B(new_n575_), .C1(new_n403_), .C2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n583_), .A2(new_n584_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n571_), .B1(new_n403_), .B2(new_n617_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n575_), .B1(new_n621_), .B2(new_n587_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n594_), .B1(new_n620_), .B2(new_n622_), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n487_), .B(new_n488_), .C1(KEYINPUT4), .C2(new_n467_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n498_), .B1(new_n493_), .B2(new_n489_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n623_), .A2(new_n602_), .A3(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n612_), .B1(new_n616_), .B2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n567_), .A2(new_n568_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n623_), .A2(new_n602_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT27), .ZN(new_n632_));
  AOI211_X1 g431(.A(new_n571_), .B(new_n574_), .C1(new_n409_), .C2(new_n546_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n583_), .A2(new_n584_), .ZN(new_n634_));
  AOI22_X1  g433(.A1(new_n633_), .A2(new_n634_), .B1(new_n574_), .B2(new_n588_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n632_), .B1(new_n635_), .B2(new_n595_), .ZN(new_n636_));
  AOI22_X1  g435(.A1(new_n631_), .A2(new_n570_), .B1(new_n636_), .B2(new_n601_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n637_), .A2(new_n569_), .A3(new_n507_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n444_), .B1(new_n630_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT100), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n605_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n444_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n596_), .A2(new_n597_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n643_), .A2(new_n626_), .A3(new_n614_), .A4(new_n615_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n569_), .B1(new_n644_), .B2(new_n612_), .ZN(new_n645_));
  OAI21_X1  g444(.A(KEYINPUT98), .B1(new_n610_), .B2(new_n611_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n499_), .A2(new_n500_), .A3(new_n504_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n604_), .A2(new_n648_), .A3(new_n629_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n642_), .B1(new_n645_), .B2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(KEYINPUT100), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n371_), .B1(new_n641_), .B2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n342_), .A2(new_n652_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n653_), .A2(G1gat), .A3(new_n507_), .ZN(new_n654_));
  XOR2_X1   g453(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n655_));
  OR2_X1    g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n655_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n641_), .A2(new_n651_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n309_), .B(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n267_), .A2(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n663_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n664_), .A2(new_n370_), .A3(new_n340_), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n661_), .A2(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(G1gat), .B1(new_n666_), .B2(new_n507_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n656_), .A2(new_n657_), .A3(new_n667_), .ZN(G1324gat));
  OAI21_X1  g467(.A(G8gat), .B1(new_n666_), .B2(new_n637_), .ZN(new_n669_));
  XOR2_X1   g468(.A(KEYINPUT103), .B(KEYINPUT39), .Z(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n342_), .A2(new_n322_), .A3(new_n604_), .A4(new_n652_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(G1325gat));
  OAI21_X1  g474(.A(G15gat), .B1(new_n666_), .B2(new_n642_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT41), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n653_), .A2(G15gat), .A3(new_n642_), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1326gat));
  OAI21_X1  g478(.A(G22gat), .B1(new_n666_), .B2(new_n629_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT42), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n629_), .A2(G22gat), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT105), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n681_), .B1(new_n653_), .B2(new_n683_), .ZN(G1327gat));
  AND2_X1   g483(.A1(new_n336_), .A2(new_n339_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(new_n309_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n272_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(new_n652_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(G29gat), .B1(new_n689_), .B2(new_n648_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n664_), .A2(new_n370_), .A3(new_n685_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n311_), .A2(new_n315_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n658_), .B2(new_n694_), .ZN(new_n695_));
  AOI211_X1 g494(.A(KEYINPUT43), .B(new_n316_), .C1(new_n641_), .C2(new_n651_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n692_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  OAI211_X1 g498(.A(new_n640_), .B(new_n642_), .C1(new_n645_), .C2(new_n649_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n569_), .A2(new_n604_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n701_), .A2(new_n444_), .A3(new_n507_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n639_), .A2(new_n640_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n694_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT43), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n658_), .A2(new_n693_), .A3(new_n694_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n708_), .A2(KEYINPUT44), .A3(new_n692_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n699_), .A2(new_n709_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n648_), .A2(G29gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n690_), .B1(new_n710_), .B2(new_n711_), .ZN(G1328gat));
  NOR3_X1   g511(.A1(new_n688_), .A2(G36gat), .A3(new_n637_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT45), .Z(new_n714_));
  NAND3_X1  g513(.A1(new_n699_), .A2(new_n604_), .A3(new_n709_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT106), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n715_), .A2(new_n716_), .A3(G36gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n715_), .B2(G36gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n714_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT46), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  OAI211_X1 g520(.A(KEYINPUT46), .B(new_n714_), .C1(new_n717_), .C2(new_n718_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1329gat));
  NAND3_X1  g522(.A1(new_n710_), .A2(G43gat), .A3(new_n444_), .ZN(new_n724_));
  INV_X1    g523(.A(G43gat), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n725_), .B1(new_n688_), .B2(new_n642_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g527(.A(G50gat), .B1(new_n689_), .B2(new_n569_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n569_), .A2(G50gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n710_), .B2(new_n730_), .ZN(G1331gat));
  NAND2_X1  g530(.A1(new_n658_), .A2(new_n371_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT107), .Z(new_n733_));
  INV_X1    g532(.A(new_n341_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n733_), .A2(new_n272_), .A3(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n735_), .B(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(G57gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n737_), .A2(new_n738_), .A3(new_n648_), .ZN(new_n739_));
  OR4_X1    g538(.A1(new_n370_), .A2(new_n661_), .A3(new_n664_), .A4(new_n685_), .ZN(new_n740_));
  OAI21_X1  g539(.A(G57gat), .B1(new_n740_), .B2(new_n507_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(G1332gat));
  INV_X1    g541(.A(G64gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n737_), .A2(new_n743_), .A3(new_n604_), .ZN(new_n744_));
  OAI21_X1  g543(.A(G64gat), .B1(new_n740_), .B2(new_n637_), .ZN(new_n745_));
  XOR2_X1   g544(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n746_));
  XNOR2_X1  g545(.A(new_n745_), .B(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n744_), .A2(new_n747_), .ZN(G1333gat));
  INV_X1    g547(.A(G71gat), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n737_), .A2(new_n749_), .A3(new_n444_), .ZN(new_n750_));
  OAI21_X1  g549(.A(G71gat), .B1(new_n740_), .B2(new_n642_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT49), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1334gat));
  INV_X1    g552(.A(G78gat), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n737_), .A2(new_n754_), .A3(new_n569_), .ZN(new_n755_));
  OAI21_X1  g554(.A(G78gat), .B1(new_n740_), .B2(new_n629_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT50), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1335gat));
  INV_X1    g557(.A(KEYINPUT112), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n761_));
  INV_X1    g560(.A(new_n269_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n762_), .A2(new_n685_), .A3(new_n371_), .A4(new_n663_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n761_), .B1(new_n708_), .B2(new_n764_), .ZN(new_n765_));
  AOI211_X1 g564(.A(KEYINPUT110), .B(new_n763_), .C1(new_n706_), .C2(new_n707_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n760_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n764_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT110), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n708_), .A2(new_n761_), .A3(new_n764_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(KEYINPUT111), .A3(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n767_), .A2(new_n648_), .A3(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(G85gat), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n686_), .A2(new_n664_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n507_), .A2(G85gat), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n733_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n759_), .B1(new_n773_), .B2(new_n777_), .ZN(new_n778_));
  AOI211_X1 g577(.A(KEYINPUT112), .B(new_n776_), .C1(new_n772_), .C2(G85gat), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n778_), .A2(new_n779_), .ZN(G1336gat));
  AND2_X1   g579(.A1(new_n733_), .A2(new_n774_), .ZN(new_n781_));
  INV_X1    g580(.A(G92gat), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(new_n782_), .A3(new_n604_), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n767_), .A2(new_n604_), .A3(new_n771_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n783_), .B1(new_n784_), .B2(new_n782_), .ZN(G1337gat));
  NAND3_X1  g584(.A1(new_n781_), .A2(new_n444_), .A3(new_n234_), .ZN(new_n786_));
  INV_X1    g585(.A(G99gat), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n642_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n786_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT51), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n786_), .B(new_n791_), .C1(new_n787_), .C2(new_n788_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(G1338gat));
  OAI21_X1  g592(.A(G106gat), .B1(new_n768_), .B2(new_n629_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT52), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n781_), .A2(new_n235_), .A3(new_n569_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n795_), .A2(new_n796_), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n797_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(G1339gat));
  NOR2_X1   g600(.A1(new_n371_), .A2(new_n433_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT118), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n370_), .A2(new_n264_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n213_), .B1(new_n212_), .B2(new_n276_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT12), .B1(new_n243_), .B2(KEYINPUT66), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n247_), .B(new_n246_), .C1(new_n810_), .C2(new_n811_), .ZN(new_n812_));
  OAI211_X1 g611(.A(KEYINPUT115), .B(new_n809_), .C1(new_n812_), .C2(new_n251_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT115), .B1(new_n250_), .B2(new_n809_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n245_), .A2(new_n248_), .A3(KEYINPUT55), .A4(new_n249_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n812_), .A2(new_n251_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n814_), .A2(new_n815_), .A3(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n808_), .B1(new_n819_), .B2(new_n259_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT56), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n807_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n812_), .A2(new_n251_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n823_), .B1(new_n824_), .B2(KEYINPUT55), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n825_), .A2(new_n813_), .A3(new_n817_), .A4(new_n816_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT116), .B1(new_n826_), .B2(new_n258_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT56), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n350_), .A2(new_n352_), .A3(new_n347_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n347_), .B1(new_n326_), .B2(new_n287_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n357_), .B1(new_n344_), .B2(new_n830_), .ZN(new_n831_));
  AOI22_X1  g630(.A1(new_n359_), .A2(new_n361_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n822_), .A2(new_n828_), .B1(new_n270_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n309_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n803_), .A2(new_n804_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n806_), .B1(new_n833_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT58), .ZN(new_n838_));
  NOR2_X1   g637(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n826_), .A2(new_n258_), .A3(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n840_), .B1(new_n826_), .B2(new_n258_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(KEYINPUT117), .A2(KEYINPUT56), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n841_), .A2(new_n842_), .A3(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n264_), .A2(new_n832_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n838_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n826_), .A2(new_n258_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n844_), .B1(new_n848_), .B2(new_n839_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n826_), .A2(new_n258_), .A3(new_n840_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n846_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(KEYINPUT58), .A3(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n847_), .A2(new_n853_), .A3(new_n694_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n270_), .A2(new_n832_), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n370_), .B(new_n264_), .C1(new_n827_), .C2(KEYINPUT56), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n820_), .A2(new_n821_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n855_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n836_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n858_), .A2(new_n859_), .A3(new_n805_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n837_), .A2(new_n854_), .A3(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n685_), .ZN(new_n862_));
  XOR2_X1   g661(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n863_));
  NAND4_X1  g662(.A1(new_n734_), .A2(new_n664_), .A3(new_n371_), .A4(new_n863_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n272_), .A2(new_n370_), .A3(new_n341_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT114), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n864_), .B1(new_n865_), .B2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n862_), .A2(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n701_), .A2(new_n444_), .A3(new_n648_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(KEYINPUT59), .B1(new_n871_), .B2(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n869_), .B1(new_n861_), .B2(new_n685_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n875_), .A2(new_n876_), .A3(new_n872_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n802_), .B1(new_n874_), .B2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n871_), .A2(new_n873_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n433_), .B1(new_n879_), .B2(new_n371_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n878_), .A2(KEYINPUT119), .A3(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n882_));
  INV_X1    g681(.A(new_n802_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n858_), .A2(new_n859_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n846_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n316_), .B1(new_n885_), .B2(KEYINPUT58), .ZN(new_n886_));
  AOI22_X1  g685(.A1(new_n884_), .A2(new_n806_), .B1(new_n886_), .B2(new_n847_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n340_), .B1(new_n887_), .B2(new_n860_), .ZN(new_n888_));
  OAI211_X1 g687(.A(KEYINPUT59), .B(new_n873_), .C1(new_n888_), .C2(new_n869_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n876_), .B1(new_n875_), .B2(new_n872_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n883_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n875_), .A2(new_n872_), .ZN(new_n892_));
  AOI21_X1  g691(.A(G113gat), .B1(new_n892_), .B2(new_n370_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n882_), .B1(new_n891_), .B2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n881_), .A2(new_n894_), .ZN(G1340gat));
  AOI21_X1  g694(.A(new_n664_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n431_), .B1(new_n664_), .B2(KEYINPUT60), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(KEYINPUT120), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT60), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(G120gat), .ZN(new_n901_));
  AND3_X1   g700(.A1(new_n892_), .A2(new_n897_), .A3(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n897_), .B1(new_n892_), .B2(new_n901_), .ZN(new_n903_));
  OAI22_X1  g702(.A1(new_n896_), .A2(new_n431_), .B1(new_n902_), .B2(new_n903_), .ZN(G1341gat));
  NOR2_X1   g703(.A1(new_n685_), .A2(new_n429_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n905_), .B1(new_n874_), .B2(new_n877_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT122), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n429_), .B1(new_n879_), .B2(new_n685_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n906_), .A2(new_n907_), .A3(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n905_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n910_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n911_));
  AOI21_X1  g710(.A(G127gat), .B1(new_n892_), .B2(new_n340_), .ZN(new_n912_));
  OAI21_X1  g711(.A(KEYINPUT122), .B1(new_n911_), .B2(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n909_), .A2(new_n913_), .ZN(G1342gat));
  OAI21_X1  g713(.A(new_n427_), .B1(new_n879_), .B2(new_n660_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(KEYINPUT123), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT123), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n917_), .B(new_n427_), .C1(new_n879_), .C2(new_n660_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n889_), .A2(new_n890_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n316_), .A2(new_n427_), .ZN(new_n920_));
  AOI22_X1  g719(.A1(new_n916_), .A2(new_n918_), .B1(new_n919_), .B2(new_n920_), .ZN(G1343gat));
  NOR4_X1   g720(.A1(new_n444_), .A2(new_n604_), .A3(new_n507_), .A4(new_n629_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n871_), .A2(new_n922_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n923_), .A2(new_n371_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(new_n460_), .ZN(G1344gat));
  NOR2_X1   g724(.A1(new_n923_), .A2(new_n664_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(new_n461_), .ZN(G1345gat));
  NOR2_X1   g726(.A1(new_n923_), .A2(new_n685_), .ZN(new_n928_));
  XOR2_X1   g727(.A(KEYINPUT61), .B(G155gat), .Z(new_n929_));
  XNOR2_X1  g728(.A(new_n928_), .B(new_n929_), .ZN(G1346gat));
  INV_X1    g729(.A(G162gat), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n923_), .A2(new_n931_), .A3(new_n316_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n923_), .B2(new_n660_), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT124), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  OAI211_X1 g734(.A(KEYINPUT124), .B(new_n931_), .C1(new_n923_), .C2(new_n660_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n932_), .B1(new_n935_), .B2(new_n936_), .ZN(G1347gat));
  NOR3_X1   g736(.A1(new_n508_), .A2(new_n569_), .A3(new_n637_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n938_), .ZN(new_n939_));
  NOR4_X1   g738(.A1(new_n875_), .A2(KEYINPUT22), .A3(new_n371_), .A4(new_n939_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT62), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n940_), .A2(new_n941_), .A3(G169gat), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n875_), .A2(new_n939_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n943_), .A2(new_n941_), .A3(new_n370_), .ZN(new_n944_));
  AND2_X1   g743(.A1(new_n944_), .A2(G169gat), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n943_), .A2(new_n370_), .ZN(new_n946_));
  OAI21_X1  g745(.A(KEYINPUT62), .B1(new_n946_), .B2(KEYINPUT22), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n942_), .B1(new_n945_), .B2(new_n947_), .ZN(G1348gat));
  NAND2_X1  g747(.A1(new_n943_), .A2(new_n272_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n949_), .B(G176gat), .ZN(G1349gat));
  INV_X1    g749(.A(new_n576_), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n943_), .A2(new_n951_), .A3(new_n340_), .ZN(new_n952_));
  AND2_X1   g751(.A1(new_n952_), .A2(KEYINPUT125), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n952_), .A2(KEYINPUT125), .ZN(new_n954_));
  AOI21_X1  g753(.A(G183gat), .B1(new_n943_), .B2(new_n340_), .ZN(new_n955_));
  NOR3_X1   g754(.A1(new_n953_), .A2(new_n954_), .A3(new_n955_), .ZN(G1350gat));
  INV_X1    g755(.A(new_n660_), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n943_), .A2(new_n577_), .A3(new_n957_), .ZN(new_n958_));
  NOR3_X1   g757(.A1(new_n875_), .A2(new_n316_), .A3(new_n939_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n958_), .B1(new_n959_), .B2(new_n383_), .ZN(G1351gat));
  NOR3_X1   g759(.A1(new_n444_), .A2(new_n648_), .A3(new_n629_), .ZN(new_n961_));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n637_), .B1(new_n961_), .B2(new_n962_), .ZN(new_n963_));
  OAI21_X1  g762(.A(new_n963_), .B1(new_n962_), .B2(new_n961_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n875_), .A2(new_n964_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n965_), .A2(new_n370_), .ZN(new_n966_));
  XNOR2_X1  g765(.A(new_n966_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g766(.A1(new_n965_), .A2(new_n272_), .ZN(new_n968_));
  XNOR2_X1  g767(.A(new_n968_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g768(.A1(new_n965_), .A2(new_n340_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n971_));
  AND2_X1   g770(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n972_));
  NOR3_X1   g771(.A1(new_n970_), .A2(new_n971_), .A3(new_n972_), .ZN(new_n973_));
  AOI21_X1  g772(.A(new_n973_), .B1(new_n970_), .B2(new_n971_), .ZN(G1354gat));
  NOR4_X1   g773(.A1(new_n875_), .A2(G218gat), .A3(new_n660_), .A4(new_n964_), .ZN(new_n975_));
  INV_X1    g774(.A(new_n975_), .ZN(new_n976_));
  INV_X1    g775(.A(G218gat), .ZN(new_n977_));
  NOR3_X1   g776(.A1(new_n875_), .A2(new_n316_), .A3(new_n964_), .ZN(new_n978_));
  OAI211_X1 g777(.A(new_n976_), .B(KEYINPUT127), .C1(new_n977_), .C2(new_n978_), .ZN(new_n979_));
  INV_X1    g778(.A(KEYINPUT127), .ZN(new_n980_));
  NOR2_X1   g779(.A1(new_n978_), .A2(new_n977_), .ZN(new_n981_));
  OAI21_X1  g780(.A(new_n980_), .B1(new_n981_), .B2(new_n975_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n979_), .A2(new_n982_), .ZN(G1355gat));
endmodule


