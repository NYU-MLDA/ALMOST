//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 0 0 1 0 0 1 1 0 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 0 1 1 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n932_, new_n933_, new_n934_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n940_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n949_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n956_, new_n957_, new_n958_,
    new_n959_;
  XNOR2_X1  g000(.A(KEYINPUT25), .B(G183gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT26), .B(G190gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G169gat), .ZN(new_n205_));
  INV_X1    g004(.A(G176gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n207_), .A2(KEYINPUT24), .A3(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n204_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G183gat), .ZN(new_n211_));
  INV_X1    g010(.A(G190gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT23), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(G183gat), .A3(G190gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n207_), .A2(KEYINPUT24), .ZN(new_n218_));
  NOR3_X1   g017(.A1(new_n210_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n211_), .A2(new_n212_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n214_), .A2(KEYINPUT81), .A3(G183gat), .A4(G190gat), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n220_), .B(new_n221_), .C1(new_n216_), .C2(KEYINPUT81), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n222_), .A2(new_n208_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT80), .B(G176gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n205_), .A2(KEYINPUT22), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT78), .B(KEYINPUT22), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(KEYINPUT79), .A3(G169gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(KEYINPUT79), .B1(new_n226_), .B2(G169gat), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n224_), .B(new_n225_), .C1(new_n228_), .C2(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n219_), .B1(new_n223_), .B2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT82), .B(G15gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G227gat), .A2(G233gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n231_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(G127gat), .B(G134gat), .Z(new_n238_));
  XOR2_X1   g037(.A(G113gat), .B(G120gat), .Z(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n231_), .A2(new_n235_), .ZN(new_n242_));
  OR3_X1    g041(.A1(new_n237_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G71gat), .B(G99gat), .Z(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(G43gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT30), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT31), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n241_), .B1(new_n237_), .B2(new_n242_), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n243_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n247_), .B1(new_n243_), .B2(new_n248_), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(G197gat), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT86), .B1(new_n253_), .B2(G204gat), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT86), .ZN(new_n255_));
  INV_X1    g054(.A(G204gat), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(new_n256_), .A3(G197gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n253_), .A2(G204gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n254_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT88), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n254_), .A2(new_n257_), .A3(KEYINPUT88), .A4(new_n258_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G211gat), .B(G218gat), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT21), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n261_), .A2(new_n262_), .A3(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT89), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT89), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n261_), .A2(new_n268_), .A3(new_n262_), .A4(new_n265_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT87), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n256_), .A2(G197gat), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT85), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n256_), .A2(G197gat), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n272_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n256_), .A2(KEYINPUT85), .A3(G197gat), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n264_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n254_), .A2(new_n257_), .A3(new_n264_), .A4(new_n258_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(new_n263_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n271_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n274_), .A2(new_n273_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n281_), .A2(new_n258_), .A3(new_n276_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT21), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n283_), .A2(KEYINPUT87), .A3(new_n263_), .A4(new_n278_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n280_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n270_), .A2(new_n285_), .ZN(new_n286_));
  XOR2_X1   g085(.A(G155gat), .B(G162gat), .Z(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT3), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G155gat), .B(G162gat), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n289_), .A2(KEYINPUT1), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G141gat), .A2(G148gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT83), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(KEYINPUT83), .A2(G141gat), .A3(G148gat), .ZN(new_n294_));
  NAND3_X1  g093(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n288_), .B1(new_n290_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(G141gat), .ZN(new_n298_));
  INV_X1    g097(.A(G148gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  OR4_X1    g100(.A1(KEYINPUT84), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT2), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n293_), .A2(new_n303_), .A3(new_n294_), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT84), .B1(new_n300_), .B2(KEYINPUT3), .ZN(new_n305_));
  NAND3_X1  g104(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n302_), .A2(new_n304_), .A3(new_n305_), .A4(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n287_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n301_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT29), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n286_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n311_), .A2(G228gat), .A3(G233gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G228gat), .A2(G233gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n286_), .A2(new_n310_), .A3(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G78gat), .B(G106gat), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n312_), .A2(new_n314_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT90), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n312_), .A2(new_n314_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n315_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n309_), .A2(KEYINPUT29), .ZN(new_n321_));
  XOR2_X1   g120(.A(G22gat), .B(G50gat), .Z(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT28), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n321_), .B(new_n323_), .ZN(new_n324_));
  AND4_X1   g123(.A1(new_n317_), .A2(new_n318_), .A3(new_n320_), .A4(new_n324_), .ZN(new_n325_));
  AOI22_X1  g124(.A1(new_n318_), .A2(new_n324_), .B1(new_n320_), .B2(new_n317_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G8gat), .B(G36gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT18), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G64gat), .B(G92gat), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n330_), .B(new_n331_), .Z(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT32), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n231_), .A2(new_n270_), .A3(new_n285_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT20), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT91), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G226gat), .A2(G233gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT19), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n221_), .B1(new_n216_), .B2(KEYINPUT81), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n342_), .A2(new_n218_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n204_), .A2(KEYINPUT92), .A3(new_n209_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT92), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n210_), .A2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n343_), .A2(new_n344_), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n216_), .A2(new_n220_), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n205_), .A2(KEYINPUT22), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n224_), .A2(new_n225_), .A3(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n348_), .A2(new_n350_), .A3(new_n208_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n347_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n286_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n335_), .A2(KEYINPUT91), .A3(KEYINPUT20), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n338_), .A2(new_n341_), .A3(new_n353_), .A4(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT95), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT20), .B1(new_n286_), .B2(new_n352_), .ZN(new_n358_));
  AOI22_X1  g157(.A1(new_n267_), .A2(new_n269_), .B1(new_n280_), .B2(new_n284_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n359_), .A2(new_n231_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n340_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n356_), .B1(new_n355_), .B2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n334_), .B1(new_n357_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT96), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  OAI211_X1 g164(.A(KEYINPUT96), .B(new_n334_), .C1(new_n357_), .C2(new_n362_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT4), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n293_), .A2(new_n294_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n370_), .B(new_n295_), .C1(KEYINPUT1), .C2(new_n289_), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n371_), .A2(new_n288_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n307_), .A2(new_n287_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n241_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n301_), .A2(new_n308_), .A3(new_n240_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n374_), .A2(KEYINPUT93), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT93), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n309_), .A2(new_n377_), .A3(new_n241_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n369_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n374_), .A2(KEYINPUT4), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n368_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G1gat), .B(G29gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G57gat), .B(G85gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n376_), .A2(new_n367_), .A3(new_n378_), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n381_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n387_), .B1(new_n381_), .B2(new_n388_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n354_), .A2(new_n353_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT20), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n392_), .B1(new_n359_), .B2(new_n231_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n393_), .A2(KEYINPUT91), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n340_), .B1(new_n391_), .B2(new_n394_), .ZN(new_n395_));
  NOR3_X1   g194(.A1(new_n358_), .A2(new_n360_), .A3(new_n340_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  OAI22_X1  g197(.A1(new_n389_), .A2(new_n390_), .B1(new_n398_), .B2(new_n334_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n365_), .A2(new_n366_), .A3(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n390_), .A2(KEYINPUT33), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT33), .ZN(new_n403_));
  OR3_X1    g202(.A1(new_n379_), .A2(new_n368_), .A3(new_n380_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n376_), .A2(new_n378_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n386_), .B1(new_n405_), .B2(new_n368_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n403_), .B1(new_n404_), .B2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n402_), .B1(new_n407_), .B2(new_n390_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n332_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n398_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n395_), .A2(new_n332_), .A3(new_n397_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n408_), .A2(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n328_), .B1(new_n401_), .B2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n389_), .A2(new_n390_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n327_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  XOR2_X1   g217(.A(new_n332_), .B(KEYINPUT97), .Z(new_n419_));
  OAI21_X1  g218(.A(new_n419_), .B1(new_n357_), .B2(new_n362_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n420_), .A2(KEYINPUT27), .A3(new_n411_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT27), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n412_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n421_), .A2(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n418_), .A2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n252_), .B1(new_n414_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n251_), .A2(new_n415_), .ZN(new_n427_));
  NOR3_X1   g226(.A1(new_n424_), .A2(new_n328_), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n426_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G229gat), .A2(G233gat), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  XOR2_X1   g231(.A(KEYINPUT73), .B(G8gat), .Z(new_n433_));
  INV_X1    g232(.A(G1gat), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT14), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G15gat), .B(G22gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G1gat), .B(G8gat), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n435_), .A2(new_n436_), .A3(new_n438_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(G29gat), .B(G36gat), .Z(new_n443_));
  XOR2_X1   g242(.A(G43gat), .B(G50gat), .Z(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n442_), .A2(new_n445_), .ZN(new_n446_));
  XOR2_X1   g245(.A(new_n443_), .B(new_n444_), .Z(new_n447_));
  AOI21_X1  g246(.A(new_n447_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n432_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n448_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n447_), .A2(KEYINPUT15), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT15), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n445_), .A2(new_n452_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n451_), .A2(new_n441_), .A3(new_n440_), .A4(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n450_), .A2(new_n454_), .A3(new_n431_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n449_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT76), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n449_), .A2(new_n455_), .A3(KEYINPUT76), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G113gat), .B(G141gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G169gat), .B(G197gat), .ZN(new_n461_));
  XOR2_X1   g260(.A(new_n460_), .B(new_n461_), .Z(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n458_), .A2(new_n459_), .A3(KEYINPUT77), .A4(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n449_), .A2(new_n455_), .A3(new_n462_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n458_), .A2(new_n459_), .A3(new_n463_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT77), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n466_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n430_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT7), .ZN(new_n472_));
  INV_X1    g271(.A(G99gat), .ZN(new_n473_));
  INV_X1    g272(.A(G106gat), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT66), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G99gat), .A2(G106gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT6), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT6), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(G99gat), .A3(G106gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT66), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n475_), .A2(new_n484_), .A3(new_n476_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n478_), .A2(new_n483_), .A3(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(G85gat), .ZN(new_n487_));
  INV_X1    g286(.A(G92gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G85gat), .A2(G92gat), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n491_), .A2(KEYINPUT8), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n480_), .A2(new_n482_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n491_), .B1(new_n493_), .B2(new_n477_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT8), .ZN(new_n495_));
  AOI22_X1  g294(.A1(new_n486_), .A2(new_n492_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  OR2_X1    g295(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n497_), .A2(new_n474_), .A3(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT64), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  AND2_X1   g300(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n502_));
  NOR2_X1   g301(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n504_), .A2(KEYINPUT64), .A3(new_n474_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n501_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT65), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n489_), .A2(KEYINPUT9), .A3(new_n490_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n490_), .A2(KEYINPUT9), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n483_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n506_), .A2(new_n507_), .A3(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n507_), .B1(new_n506_), .B2(new_n510_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n496_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT68), .ZN(new_n514_));
  AOI21_X1  g313(.A(KEYINPUT64), .B1(new_n504_), .B2(new_n474_), .ZN(new_n515_));
  NOR4_X1   g314(.A1(new_n502_), .A2(new_n503_), .A3(new_n500_), .A4(G106gat), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n483_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT65), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n506_), .A2(new_n510_), .A3(new_n507_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT68), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n521_), .A2(new_n522_), .A3(new_n496_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n514_), .A2(new_n523_), .A3(new_n451_), .A4(new_n453_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n521_), .A2(new_n445_), .A3(new_n496_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G232gat), .A2(G233gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT35), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n525_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n524_), .A2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n528_), .A2(new_n529_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n532_), .B(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G190gat), .B(G218gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G134gat), .B(G162gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n538_), .B(KEYINPUT36), .Z(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT72), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n535_), .A2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n538_), .A2(KEYINPUT36), .ZN(new_n542_));
  AOI21_X1  g341(.A(KEYINPUT71), .B1(new_n535_), .B2(new_n542_), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n532_), .A2(new_n533_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n532_), .A2(new_n533_), .ZN(new_n545_));
  AND4_X1   g344(.A1(KEYINPUT71), .A2(new_n544_), .A3(new_n542_), .A4(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n541_), .B1(new_n543_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT37), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n541_), .B(KEYINPUT37), .C1(new_n543_), .C2(new_n546_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G231gat), .A2(G233gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n442_), .B(new_n552_), .ZN(new_n553_));
  XOR2_X1   g352(.A(G71gat), .B(G78gat), .Z(new_n554_));
  XNOR2_X1  g353(.A(G57gat), .B(G64gat), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n554_), .B1(KEYINPUT11), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT67), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(new_n557_), .A3(KEYINPUT11), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n557_), .B1(new_n555_), .B2(KEYINPUT11), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n556_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(G57gat), .B(G64gat), .Z(new_n562_));
  INV_X1    g361(.A(KEYINPUT11), .ZN(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT67), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n563_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n564_), .A2(new_n565_), .A3(new_n554_), .A4(new_n558_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n561_), .A2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n553_), .B(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT74), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G127gat), .B(G155gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT16), .ZN(new_n572_));
  XOR2_X1   g371(.A(G183gat), .B(G211gat), .Z(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(KEYINPUT17), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n570_), .A2(new_n576_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n568_), .A2(new_n569_), .A3(KEYINPUT17), .A4(new_n575_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  OR3_X1    g378(.A1(new_n568_), .A2(KEYINPUT17), .A3(new_n575_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT75), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT75), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n579_), .A2(new_n583_), .A3(new_n580_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n551_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n567_), .ZN(new_n587_));
  AOI21_X1  g386(.A(KEYINPUT12), .B1(new_n513_), .B2(new_n587_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n567_), .B(new_n496_), .C1(new_n511_), .C2(new_n512_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G230gat), .A2(G233gat), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT12), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n567_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n514_), .A2(new_n523_), .A3(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n591_), .A2(new_n592_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n592_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n567_), .B1(new_n521_), .B2(new_n496_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n597_), .B1(new_n590_), .B2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G120gat), .B(G148gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT5), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G176gat), .B(G204gat), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n601_), .B(new_n602_), .Z(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n596_), .A2(new_n599_), .A3(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT69), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n596_), .A2(KEYINPUT69), .A3(new_n599_), .A4(new_n604_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n596_), .A2(new_n599_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n609_), .B1(new_n610_), .B2(new_n604_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT13), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n611_), .A2(new_n612_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n586_), .A2(new_n615_), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n471_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(KEYINPUT98), .ZN(new_n618_));
  OR3_X1    g417(.A1(new_n471_), .A2(KEYINPUT98), .A3(new_n616_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(new_n434_), .A3(new_n416_), .ZN(new_n621_));
  XOR2_X1   g420(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n615_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n470_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n581_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n625_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n430_), .A2(new_n628_), .A3(new_n547_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G1gat), .B1(new_n630_), .B2(new_n415_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n620_), .A2(new_n434_), .A3(new_n416_), .A4(new_n622_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n624_), .A2(new_n631_), .A3(new_n632_), .ZN(G1324gat));
  XNOR2_X1  g432(.A(KEYINPUT101), .B(KEYINPUT39), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n430_), .A2(new_n628_), .A3(new_n424_), .A4(new_n547_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(G8gat), .B1(new_n636_), .B2(new_n637_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n635_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n629_), .A2(KEYINPUT100), .A3(new_n424_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n642_), .A2(G8gat), .A3(new_n634_), .A4(new_n638_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n618_), .A2(new_n424_), .A3(new_n433_), .A4(new_n619_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n644_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n646_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(G1325gat));
  INV_X1    g448(.A(G15gat), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n650_), .B1(new_n629_), .B2(new_n251_), .ZN(new_n651_));
  XOR2_X1   g450(.A(KEYINPUT103), .B(KEYINPUT41), .Z(new_n652_));
  OR2_X1    g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n652_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n251_), .A2(new_n650_), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n653_), .B(new_n654_), .C1(new_n617_), .C2(new_n655_), .ZN(G1326gat));
  INV_X1    g455(.A(G22gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n657_), .B1(new_n629_), .B2(new_n328_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT42), .Z(new_n659_));
  NAND2_X1  g458(.A1(new_n328_), .A2(new_n657_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT104), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n659_), .B1(new_n617_), .B2(new_n661_), .ZN(G1327gat));
  INV_X1    g461(.A(new_n585_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n663_), .A2(new_n547_), .ZN(new_n664_));
  AND4_X1   g463(.A1(new_n430_), .A2(new_n470_), .A3(new_n615_), .A4(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n415_), .A2(G29gat), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT106), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  XOR2_X1   g467(.A(KEYINPUT105), .B(KEYINPUT43), .Z(new_n669_));
  NAND3_X1  g468(.A1(new_n417_), .A2(new_n421_), .A3(new_n423_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n408_), .A2(new_n412_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n399_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n672_), .B2(new_n366_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n670_), .B1(new_n673_), .B2(new_n328_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n428_), .B1(new_n674_), .B2(new_n252_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n551_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n669_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT43), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n401_), .A2(new_n413_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(new_n327_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n251_), .B1(new_n680_), .B2(new_n670_), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n678_), .B(new_n551_), .C1(new_n681_), .C2(new_n428_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n677_), .A2(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n615_), .A2(new_n470_), .A3(new_n585_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT44), .B1(new_n683_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687_));
  AOI211_X1 g486(.A(new_n687_), .B(new_n684_), .C1(new_n677_), .C2(new_n682_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n686_), .A2(new_n688_), .A3(new_n415_), .ZN(new_n689_));
  INV_X1    g488(.A(G29gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n668_), .B1(new_n689_), .B2(new_n690_), .ZN(G1328gat));
  NOR2_X1   g490(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n692_));
  INV_X1    g491(.A(G36gat), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n686_), .A2(new_n688_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n694_), .B2(new_n424_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n665_), .A2(new_n693_), .A3(new_n424_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT45), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n696_), .B(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n692_), .B1(new_n695_), .B2(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n696_), .B(KEYINPUT45), .ZN(new_n700_));
  INV_X1    g499(.A(new_n692_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n424_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n686_), .A2(new_n688_), .A3(new_n702_), .ZN(new_n703_));
  OAI211_X1 g502(.A(new_n700_), .B(new_n701_), .C1(new_n703_), .C2(new_n693_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n699_), .A2(new_n704_), .ZN(G1329gat));
  NAND2_X1  g504(.A1(new_n251_), .A2(G43gat), .ZN(new_n706_));
  NOR3_X1   g505(.A1(new_n686_), .A2(new_n688_), .A3(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(G43gat), .B1(new_n665_), .B2(new_n251_), .ZN(new_n708_));
  OR3_X1    g507(.A1(new_n707_), .A2(KEYINPUT47), .A3(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(KEYINPUT47), .B1(new_n707_), .B2(new_n708_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1330gat));
  AOI21_X1  g510(.A(G50gat), .B1(new_n665_), .B2(new_n328_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n328_), .A2(G50gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n694_), .B2(new_n713_), .ZN(G1331gat));
  NAND2_X1  g513(.A1(new_n430_), .A2(new_n626_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n615_), .B1(new_n715_), .B2(KEYINPUT108), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT108), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n430_), .A2(new_n717_), .A3(new_n626_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n716_), .A2(new_n586_), .A3(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n415_), .A2(G57gat), .ZN(new_n721_));
  INV_X1    g520(.A(new_n547_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n675_), .A2(new_n722_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n615_), .A2(new_n470_), .A3(new_n585_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n723_), .A2(new_n416_), .A3(new_n724_), .ZN(new_n725_));
  AOI22_X1  g524(.A1(new_n720_), .A2(new_n721_), .B1(G57gat), .B2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT109), .ZN(G1332gat));
  NAND2_X1  g526(.A1(new_n723_), .A2(new_n724_), .ZN(new_n728_));
  OAI21_X1  g527(.A(G64gat), .B1(new_n728_), .B2(new_n702_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n729_), .A2(KEYINPUT48), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(KEYINPUT48), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n702_), .A2(G64gat), .ZN(new_n732_));
  OAI22_X1  g531(.A1(new_n730_), .A2(new_n731_), .B1(new_n719_), .B2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT110), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n735_));
  OAI221_X1 g534(.A(new_n735_), .B1(new_n719_), .B2(new_n732_), .C1(new_n730_), .C2(new_n731_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(G1333gat));
  OAI21_X1  g536(.A(G71gat), .B1(new_n728_), .B2(new_n252_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT49), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n252_), .A2(G71gat), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT111), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n739_), .B1(new_n719_), .B2(new_n741_), .ZN(G1334gat));
  OAI21_X1  g541(.A(G78gat), .B1(new_n728_), .B2(new_n327_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT50), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n327_), .A2(G78gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n744_), .B1(new_n719_), .B2(new_n745_), .ZN(G1335gat));
  OAI211_X1 g545(.A(new_n585_), .B(new_n626_), .C1(new_n613_), .C2(new_n614_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT112), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n683_), .A2(new_n749_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n415_), .A2(new_n487_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT113), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n750_), .A2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT108), .B1(new_n675_), .B2(new_n470_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n754_), .A2(new_n718_), .A3(new_n625_), .A4(new_n664_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n416_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n753_), .B1(new_n757_), .B2(new_n487_), .ZN(G1336gat));
  NAND3_X1  g557(.A1(new_n756_), .A2(new_n488_), .A3(new_n424_), .ZN(new_n759_));
  OAI21_X1  g558(.A(G92gat), .B1(new_n750_), .B2(new_n702_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(G1337gat));
  NAND3_X1  g560(.A1(new_n756_), .A2(new_n251_), .A3(new_n504_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n683_), .A2(new_n251_), .A3(new_n749_), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n763_), .A2(KEYINPUT114), .A3(G99gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(KEYINPUT114), .B1(new_n763_), .B2(G99gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n762_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT51), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n762_), .B(new_n768_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1338gat));
  XNOR2_X1  g569(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n771_));
  AOI211_X1 g570(.A(new_n327_), .B(new_n748_), .C1(new_n677_), .C2(new_n682_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774_));
  OAI21_X1  g573(.A(G106gat), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  OAI22_X1  g574(.A1(new_n772_), .A2(new_n775_), .B1(KEYINPUT115), .B2(KEYINPUT52), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n683_), .A2(new_n328_), .A3(new_n749_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n777_), .A2(new_n773_), .A3(new_n774_), .A4(G106gat), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n328_), .A2(new_n474_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n755_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n771_), .B1(new_n779_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n771_), .ZN(new_n784_));
  AOI211_X1 g583(.A(new_n781_), .B(new_n784_), .C1(new_n776_), .C2(new_n778_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n783_), .A2(new_n785_), .ZN(G1339gat));
  NAND2_X1  g585(.A1(new_n702_), .A2(new_n327_), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n787_), .A2(new_n415_), .A3(new_n252_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT56), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n514_), .A2(new_n523_), .A3(new_n594_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n589_), .B1(new_n598_), .B2(KEYINPUT12), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n597_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT117), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n513_), .A2(new_n587_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n593_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n595_), .A2(new_n589_), .A3(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT117), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(new_n798_), .A3(new_n597_), .ZN(new_n799_));
  AND4_X1   g598(.A1(KEYINPUT55), .A2(new_n591_), .A3(new_n592_), .A4(new_n595_), .ZN(new_n800_));
  AOI22_X1  g599(.A1(new_n794_), .A2(new_n799_), .B1(new_n800_), .B2(KEYINPUT118), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n591_), .A2(KEYINPUT55), .A3(new_n592_), .A4(new_n595_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT118), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n596_), .A2(new_n805_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n804_), .A2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n604_), .B1(new_n801_), .B2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n790_), .B1(new_n808_), .B2(KEYINPUT119), .ZN(new_n809_));
  AOI211_X1 g608(.A(KEYINPUT117), .B(new_n592_), .C1(new_n591_), .C2(new_n595_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n798_), .B1(new_n797_), .B2(new_n597_), .ZN(new_n811_));
  OAI22_X1  g610(.A1(new_n810_), .A2(new_n811_), .B1(new_n803_), .B2(new_n802_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n804_), .A2(new_n806_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n603_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT119), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n814_), .A2(new_n815_), .A3(KEYINPUT56), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n470_), .A2(new_n609_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n809_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n431_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n450_), .A2(new_n454_), .A3(new_n432_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n820_), .A3(new_n463_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT120), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n822_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n465_), .A3(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n611_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n818_), .A2(new_n827_), .ZN(new_n828_));
  AND4_X1   g627(.A1(KEYINPUT122), .A2(new_n828_), .A3(KEYINPUT57), .A4(new_n547_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n722_), .B1(new_n818_), .B2(new_n827_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT122), .B1(new_n830_), .B2(KEYINPUT57), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n829_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT58), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n790_), .B(new_n603_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n825_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n794_), .A2(new_n799_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n800_), .A2(KEYINPUT118), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n837_), .A2(new_n804_), .A3(new_n806_), .A4(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n790_), .B1(new_n839_), .B2(new_n603_), .ZN(new_n840_));
  OAI211_X1 g639(.A(KEYINPUT121), .B(new_n833_), .C1(new_n836_), .C2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n551_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n814_), .A2(KEYINPUT56), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n843_), .A2(new_n834_), .A3(new_n835_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n833_), .B1(new_n844_), .B2(KEYINPUT121), .ZN(new_n845_));
  OAI22_X1  g644(.A1(new_n830_), .A2(KEYINPUT57), .B1(new_n842_), .B2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n627_), .B1(new_n832_), .B2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT54), .B1(new_n616_), .B2(new_n470_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n586_), .A2(new_n849_), .A3(new_n626_), .A4(new_n615_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n789_), .B1(new_n847_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(G113gat), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(new_n853_), .A3(new_n470_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n828_), .A2(KEYINPUT57), .A3(new_n547_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n830_), .A2(KEYINPUT122), .A3(KEYINPUT57), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n846_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n851_), .B1(new_n860_), .B2(new_n581_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n855_), .B1(new_n861_), .B2(new_n788_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n788_), .A2(new_n855_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n585_), .B1(new_n832_), .B2(new_n846_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(new_n851_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n862_), .A2(new_n865_), .A3(new_n626_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n854_), .B1(new_n866_), .B2(new_n853_), .ZN(G1340gat));
  NOR3_X1   g666(.A1(new_n862_), .A2(new_n865_), .A3(new_n615_), .ZN(new_n868_));
  INV_X1    g667(.A(G120gat), .ZN(new_n869_));
  INV_X1    g668(.A(new_n852_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n615_), .B2(KEYINPUT60), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n871_), .B1(KEYINPUT60), .B2(new_n869_), .ZN(new_n872_));
  OAI22_X1  g671(.A1(new_n868_), .A2(new_n869_), .B1(new_n870_), .B2(new_n872_), .ZN(G1341gat));
  INV_X1    g672(.A(G127gat), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n627_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n862_), .A2(new_n865_), .A3(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(G127gat), .B1(new_n852_), .B2(new_n663_), .ZN(new_n878_));
  OAI21_X1  g677(.A(KEYINPUT123), .B1(new_n877_), .B2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n864_), .A2(new_n851_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n789_), .A2(KEYINPUT59), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n882_), .B(new_n875_), .C1(new_n855_), .C2(new_n852_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT123), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n861_), .A2(new_n663_), .A3(new_n788_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n874_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n883_), .A2(new_n884_), .A3(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n879_), .A2(new_n887_), .ZN(G1342gat));
  INV_X1    g687(.A(G134gat), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n852_), .A2(new_n889_), .A3(new_n722_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n862_), .A2(new_n865_), .A3(new_n676_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n889_), .ZN(G1343gat));
  INV_X1    g691(.A(new_n861_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n328_), .A2(new_n252_), .A3(new_n416_), .ZN(new_n894_));
  OR3_X1    g693(.A1(new_n893_), .A2(new_n424_), .A3(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(G141gat), .B1(new_n895_), .B2(new_n626_), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n893_), .A2(new_n424_), .A3(new_n894_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n897_), .A2(new_n298_), .A3(new_n470_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n896_), .A2(new_n898_), .ZN(G1344gat));
  XNOR2_X1  g698(.A(KEYINPUT124), .B(G148gat), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n901_), .B1(new_n895_), .B2(new_n615_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n897_), .A2(new_n625_), .A3(new_n900_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1345gat));
  XNOR2_X1  g703(.A(KEYINPUT61), .B(G155gat), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n905_), .B1(new_n895_), .B2(new_n585_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n905_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n897_), .A2(new_n663_), .A3(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n908_), .ZN(G1346gat));
  OAI21_X1  g708(.A(G162gat), .B1(new_n895_), .B2(new_n676_), .ZN(new_n910_));
  INV_X1    g709(.A(G162gat), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n897_), .A2(new_n911_), .A3(new_n722_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n910_), .A2(new_n912_), .ZN(G1347gat));
  NOR2_X1   g712(.A1(new_n702_), .A2(new_n427_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(new_n328_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n880_), .A2(new_n470_), .A3(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(G169gat), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n917_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n349_), .A2(new_n225_), .ZN(new_n922_));
  OAI211_X1 g721(.A(new_n920_), .B(new_n921_), .C1(new_n922_), .C2(new_n917_), .ZN(G1348gat));
  NAND3_X1  g722(.A1(new_n880_), .A2(new_n625_), .A3(new_n916_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n224_), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT125), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n925_), .A2(new_n926_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n924_), .A2(KEYINPUT125), .A3(new_n224_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n893_), .A2(new_n328_), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n915_), .A2(new_n206_), .A3(new_n615_), .ZN(new_n930_));
  AOI22_X1  g729(.A1(new_n927_), .A2(new_n928_), .B1(new_n929_), .B2(new_n930_), .ZN(G1349gat));
  NAND3_X1  g730(.A1(new_n929_), .A2(new_n663_), .A3(new_n914_), .ZN(new_n932_));
  AND2_X1   g731(.A1(new_n880_), .A2(new_n916_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n627_), .A2(new_n202_), .ZN(new_n934_));
  AOI22_X1  g733(.A1(new_n932_), .A2(new_n211_), .B1(new_n933_), .B2(new_n934_), .ZN(G1350gat));
  NAND2_X1  g734(.A1(new_n722_), .A2(new_n203_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(KEYINPUT126), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n933_), .A2(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n933_), .A2(new_n551_), .ZN(new_n939_));
  INV_X1    g738(.A(new_n939_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n938_), .B1(new_n940_), .B2(new_n212_), .ZN(G1351gat));
  NOR3_X1   g740(.A1(new_n702_), .A2(new_n418_), .A3(new_n251_), .ZN(new_n942_));
  AND2_X1   g741(.A1(new_n861_), .A2(new_n942_), .ZN(new_n943_));
  AOI21_X1  g742(.A(G197gat), .B1(new_n943_), .B2(new_n470_), .ZN(new_n944_));
  NAND4_X1  g743(.A1(new_n861_), .A2(G197gat), .A3(new_n470_), .A4(new_n942_), .ZN(new_n945_));
  AND2_X1   g744(.A1(new_n945_), .A2(KEYINPUT127), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n945_), .A2(KEYINPUT127), .ZN(new_n947_));
  NOR3_X1   g746(.A1(new_n944_), .A2(new_n946_), .A3(new_n947_), .ZN(G1352gat));
  NAND2_X1  g747(.A1(new_n943_), .A2(new_n625_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n949_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g749(.A1(new_n943_), .A2(new_n581_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(KEYINPUT63), .B(G211gat), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n951_), .A2(new_n952_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n953_), .B1(new_n951_), .B2(new_n954_), .ZN(G1354gat));
  INV_X1    g754(.A(G218gat), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n943_), .A2(new_n956_), .A3(new_n722_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n943_), .A2(new_n551_), .ZN(new_n958_));
  INV_X1    g757(.A(new_n958_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n957_), .B1(new_n959_), .B2(new_n956_), .ZN(G1355gat));
endmodule


