//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 1 1 1 0 0 0 0 1 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n772_, new_n773_, new_n774_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n804_, new_n805_, new_n806_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n821_, new_n822_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n945_, new_n946_, new_n948_, new_n949_,
    new_n951_, new_n952_, new_n953_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n974_, new_n976_, new_n978_,
    new_n979_, new_n980_, new_n982_, new_n983_, new_n985_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n992_, new_n993_, new_n994_;
  XOR2_X1   g000(.A(G29gat), .B(G36gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G43gat), .B(G50gat), .Z(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G29gat), .B(G36gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G43gat), .B(G50gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT15), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n211_));
  INV_X1    g010(.A(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G85gat), .ZN(new_n215_));
  INV_X1    g014(.A(G92gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G85gat), .A2(G92gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(KEYINPUT9), .A3(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT9), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n220_), .A2(G85gat), .A3(G92gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n214_), .A2(new_n219_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT7), .ZN(new_n223_));
  INV_X1    g022(.A(G99gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(new_n224_), .A3(new_n212_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT8), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n222_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT64), .B(KEYINPUT6), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G99gat), .A2(G106gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(KEYINPUT64), .A2(KEYINPUT6), .ZN(new_n233_));
  INV_X1    g032(.A(new_n231_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(KEYINPUT64), .A2(KEYINPUT6), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n232_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n229_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n217_), .A2(new_n218_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(new_n226_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n242_), .A2(KEYINPUT6), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT6), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n244_), .A2(KEYINPUT65), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n234_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(KEYINPUT65), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n242_), .A2(KEYINPUT6), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n247_), .A2(new_n248_), .A3(new_n231_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n246_), .A2(new_n225_), .A3(new_n227_), .A4(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n239_), .A2(new_n226_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n241_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n210_), .B1(new_n238_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n238_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n204_), .A2(new_n207_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G232gat), .A2(G233gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT34), .ZN(new_n257_));
  OAI22_X1  g056(.A1(new_n254_), .A2(new_n255_), .B1(KEYINPUT35), .B2(new_n257_), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n253_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n257_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT35), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n259_), .A2(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n253_), .A2(new_n258_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n262_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n263_), .A2(new_n266_), .ZN(new_n267_));
  XOR2_X1   g066(.A(G190gat), .B(G218gat), .Z(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT72), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G134gat), .B(G162gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  XOR2_X1   g070(.A(new_n271_), .B(KEYINPUT36), .Z(new_n272_));
  AND2_X1   g071(.A1(new_n267_), .A2(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n274_));
  NAND2_X1  g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(new_n275_), .B(KEYINPUT74), .Z(new_n276_));
  NAND3_X1  g075(.A1(new_n276_), .A2(new_n263_), .A3(new_n266_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n273_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT89), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G227gat), .A2(G233gat), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n282_), .B(KEYINPUT84), .Z(new_n283_));
  INV_X1    g082(.A(G15gat), .ZN(new_n284_));
  INV_X1    g083(.A(G43gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G15gat), .A2(G43gat), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n286_), .A2(KEYINPUT83), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(KEYINPUT83), .B1(new_n286_), .B2(new_n287_), .ZN(new_n290_));
  OAI21_X1  g089(.A(G71gat), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n286_), .A2(new_n287_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT83), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(G71gat), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(new_n295_), .A3(new_n288_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n291_), .A2(G99gat), .A3(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(G99gat), .B1(new_n291_), .B2(new_n296_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n283_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NOR3_X1   g099(.A1(new_n289_), .A2(G71gat), .A3(new_n290_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n295_), .B1(new_n294_), .B2(new_n288_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n224_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n283_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n303_), .A2(new_n304_), .A3(new_n297_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n300_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(G169gat), .ZN(new_n307_));
  INV_X1    g106(.A(G176gat), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT24), .ZN(new_n310_));
  NOR2_X1   g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311_));
  NOR3_X1   g110(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n310_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G183gat), .A2(G190gat), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT23), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n313_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n312_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT25), .B(G183gat), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT26), .ZN(new_n321_));
  INV_X1    g120(.A(G190gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT81), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT81), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(G190gat), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n321_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n320_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n323_), .A2(new_n325_), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n316_), .B(new_n317_), .C1(new_n329_), .C2(G183gat), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT22), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n308_), .B1(new_n331_), .B2(KEYINPUT82), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(new_n307_), .ZN(new_n333_));
  OAI211_X1 g132(.A(G169gat), .B(new_n308_), .C1(new_n331_), .C2(KEYINPUT82), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  AOI22_X1  g134(.A1(new_n319_), .A2(new_n328_), .B1(new_n330_), .B2(new_n335_), .ZN(new_n336_));
  OR2_X1    g135(.A1(new_n336_), .A2(KEYINPUT30), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(KEYINPUT30), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n337_), .A2(KEYINPUT85), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT85), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n336_), .A2(KEYINPUT30), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n319_), .A2(new_n328_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n330_), .A2(new_n335_), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n342_), .A2(KEYINPUT30), .A3(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n340_), .B1(new_n341_), .B2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n306_), .A2(new_n339_), .A3(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n341_), .A2(new_n344_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n347_), .A2(KEYINPUT85), .A3(new_n300_), .A4(new_n305_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT31), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G113gat), .B(G120gat), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(G134gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(G127gat), .ZN(new_n354_));
  INV_X1    g153(.A(G127gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(G134gat), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n354_), .A2(new_n356_), .A3(KEYINPUT87), .ZN(new_n357_));
  AOI21_X1  g156(.A(KEYINPUT87), .B1(new_n354_), .B2(new_n356_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n352_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT87), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n355_), .A2(G134gat), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n353_), .A2(G127gat), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n360_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n354_), .A2(new_n356_), .A3(KEYINPUT87), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n363_), .A2(new_n364_), .A3(new_n351_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n359_), .A2(new_n365_), .A3(KEYINPUT88), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(KEYINPUT88), .B1(new_n359_), .B2(new_n365_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n350_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n368_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(KEYINPUT31), .A3(new_n366_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n281_), .B1(new_n349_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT86), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n346_), .A2(new_n348_), .A3(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n372_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n375_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n374_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n349_), .A2(KEYINPUT86), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n380_), .A2(new_n281_), .A3(new_n372_), .A4(new_n376_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  XOR2_X1   g181(.A(KEYINPUT92), .B(G233gat), .Z(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(G228gat), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT94), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n384_), .A2(KEYINPUT94), .ZN(new_n388_));
  OR2_X1    g187(.A1(G197gat), .A2(G204gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G197gat), .A2(G204gat), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(G211gat), .B(G218gat), .Z(new_n392_));
  INV_X1    g191(.A(KEYINPUT93), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n391_), .A2(new_n392_), .A3(new_n393_), .A4(KEYINPUT21), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n389_), .A2(KEYINPUT21), .A3(new_n390_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G211gat), .B(G218gat), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT93), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n394_), .A2(new_n397_), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n395_), .A2(new_n396_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n389_), .A2(new_n390_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT21), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n399_), .A2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n388_), .B1(new_n398_), .B2(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(G155gat), .A2(G162gat), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G155gat), .A2(G162gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT90), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT3), .ZN(new_n411_));
  INV_X1    g210(.A(G141gat), .ZN(new_n412_));
  INV_X1    g211(.A(G148gat), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n411_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n415_));
  NAND3_X1  g214(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n414_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n408_), .B1(new_n410_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n412_), .A2(new_n413_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G141gat), .A2(G148gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n405_), .B1(KEYINPUT1), .B2(new_n407_), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n407_), .A2(KEYINPUT1), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n422_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT29), .B1(new_n419_), .B2(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n387_), .B1(new_n404_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G78gat), .B(G106gat), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n404_), .A2(new_n426_), .A3(new_n387_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n428_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n404_), .A2(new_n426_), .A3(new_n387_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n429_), .B1(new_n433_), .B2(new_n427_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT95), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT90), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n409_), .B(new_n437_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n406_), .B(new_n407_), .C1(new_n438_), .C2(new_n417_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n425_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT28), .B1(new_n441_), .B2(KEYINPUT29), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n419_), .A2(new_n425_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT28), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT29), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n443_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G22gat), .B(G50gat), .ZN(new_n447_));
  XOR2_X1   g246(.A(new_n447_), .B(KEYINPUT91), .Z(new_n448_));
  AND3_X1   g247(.A1(new_n442_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n448_), .B1(new_n442_), .B2(new_n446_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n436_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n442_), .A2(new_n446_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n448_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n442_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(KEYINPUT95), .A3(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n435_), .A2(new_n451_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n454_), .A2(new_n455_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n458_), .A2(new_n434_), .A3(new_n436_), .A4(new_n432_), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G226gat), .A2(G233gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT19), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n342_), .A2(new_n343_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n398_), .A2(new_n403_), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT20), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n397_), .A2(new_n394_), .B1(new_n399_), .B2(new_n402_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n327_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT96), .ZN(new_n468_));
  NAND2_X1  g267(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n468_), .B1(new_n467_), .B2(new_n469_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n320_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n312_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n318_), .A2(KEYINPUT97), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n316_), .A2(new_n317_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT97), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n475_), .A2(new_n476_), .A3(new_n313_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .A4(new_n477_), .ZN(new_n478_));
  XOR2_X1   g277(.A(KEYINPUT22), .B(G169gat), .Z(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n309_), .B1(new_n480_), .B2(new_n308_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n475_), .B1(G183gat), .B2(G190gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n466_), .B1(new_n478_), .B2(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n462_), .B1(new_n465_), .B2(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(G8gat), .B(G36gat), .Z(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT18), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G64gat), .B(G92gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT20), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n490_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n462_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n478_), .A2(new_n466_), .A3(new_n483_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n485_), .A2(new_n489_), .A3(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n489_), .B1(new_n485_), .B2(new_n494_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT100), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n441_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n359_), .A2(new_n365_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n443_), .A2(new_n501_), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n500_), .A2(KEYINPUT4), .A3(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(KEYINPUT98), .B(KEYINPUT4), .Z(new_n504_));
  OAI211_X1 g303(.A(new_n441_), .B(new_n504_), .C1(new_n367_), .C2(new_n368_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G225gat), .A2(G233gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n499_), .B1(new_n503_), .B2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n500_), .A2(KEYINPUT4), .A3(new_n502_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n509_), .A2(KEYINPUT100), .A3(new_n506_), .A4(new_n505_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT99), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n443_), .B1(new_n370_), .B2(new_n366_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n501_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n441_), .A2(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n511_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n500_), .A2(KEYINPUT99), .A3(new_n502_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n506_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n515_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G1gat), .B(G29gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(G85gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT0), .B(G57gat), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n520_), .B(new_n521_), .Z(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n508_), .A2(new_n510_), .A3(new_n518_), .A4(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n500_), .A2(new_n502_), .A3(new_n506_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n505_), .A2(new_n517_), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n522_), .B(new_n525_), .C1(new_n503_), .C2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT33), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n509_), .A2(new_n517_), .A3(new_n505_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n530_), .A2(KEYINPUT33), .A3(new_n522_), .A4(new_n525_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n498_), .A2(new_n524_), .A3(new_n529_), .A4(new_n531_), .ZN(new_n532_));
  NOR3_X1   g331(.A1(new_n465_), .A2(new_n484_), .A3(new_n462_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n492_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n534_));
  OAI211_X1 g333(.A(KEYINPUT32), .B(new_n489_), .C1(new_n533_), .C2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n489_), .A2(KEYINPUT32), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n485_), .A2(new_n494_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n527_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n522_), .B1(new_n530_), .B2(new_n525_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n535_), .B(new_n537_), .C1(new_n538_), .C2(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n460_), .B1(new_n532_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n530_), .A2(new_n525_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(new_n523_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n457_), .A2(new_n543_), .A3(new_n459_), .A4(new_n527_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT27), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n545_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n489_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n547_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n548_), .A2(KEYINPUT27), .A3(new_n495_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n546_), .A2(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n544_), .A2(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n382_), .B1(new_n541_), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT101), .ZN(new_n553_));
  AND3_X1   g352(.A1(new_n548_), .A2(KEYINPUT27), .A3(new_n495_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n478_), .A2(new_n483_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(new_n464_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n490_), .B1(new_n466_), .B2(new_n336_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n492_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n547_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(KEYINPUT27), .B1(new_n560_), .B2(new_n495_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n553_), .B1(new_n554_), .B2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n546_), .A2(new_n549_), .A3(KEYINPUT101), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n460_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n538_), .A2(new_n539_), .ZN(new_n565_));
  AND3_X1   g364(.A1(new_n379_), .A2(new_n565_), .A3(new_n381_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n280_), .B1(new_n552_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT13), .ZN(new_n569_));
  XOR2_X1   g368(.A(G120gat), .B(G148gat), .Z(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT71), .ZN(new_n571_));
  XOR2_X1   g370(.A(G176gat), .B(G204gat), .Z(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n573_), .B(new_n574_), .Z(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G57gat), .B(G64gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G71gat), .B(G78gat), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n577_), .A2(new_n578_), .A3(KEYINPUT11), .ZN(new_n579_));
  INV_X1    g378(.A(new_n578_), .ZN(new_n580_));
  INV_X1    g379(.A(G64gat), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(G57gat), .ZN(new_n582_));
  INV_X1    g381(.A(G57gat), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(G64gat), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n582_), .A2(new_n584_), .A3(KEYINPUT11), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n580_), .A2(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n577_), .A2(KEYINPUT11), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n579_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n247_), .A2(new_n248_), .A3(new_n231_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n231_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n225_), .A2(new_n227_), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n590_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n251_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n240_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n232_), .A2(new_n236_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n596_), .B1(new_n228_), .B2(new_n222_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n589_), .B1(new_n595_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT67), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n252_), .A2(new_n238_), .A3(new_n588_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT66), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n252_), .A2(new_n238_), .A3(KEYINPUT66), .A4(new_n588_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n254_), .A2(KEYINPUT67), .A3(new_n589_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n600_), .A2(new_n603_), .A3(new_n604_), .A4(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(G230gat), .ZN(new_n607_));
  INV_X1    g406(.A(G233gat), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n606_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT68), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n606_), .A2(KEYINPUT68), .A3(new_n609_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(KEYINPUT69), .B(KEYINPUT12), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n616_), .B1(new_n254_), .B2(new_n589_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT12), .ZN(new_n618_));
  AOI211_X1 g417(.A(new_n618_), .B(new_n588_), .C1(new_n252_), .C2(new_n238_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n609_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n601_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n620_), .A2(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n576_), .B1(new_n614_), .B2(new_n624_), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n606_), .A2(KEYINPUT68), .A3(new_n609_), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT68), .B1(new_n606_), .B2(new_n609_), .ZN(new_n627_));
  OAI211_X1 g426(.A(new_n624_), .B(new_n576_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n569_), .B1(new_n625_), .B2(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n624_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(new_n575_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(KEYINPUT13), .A3(new_n628_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n630_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(G231gat), .A2(G233gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n588_), .B(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(G1gat), .B(G8gat), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n637_), .A2(KEYINPUT76), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(KEYINPUT76), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(G15gat), .B(G22gat), .ZN(new_n641_));
  NAND2_X1  g440(.A1(G1gat), .A2(G8gat), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT14), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n640_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n644_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n638_), .A2(new_n646_), .A3(new_n639_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n636_), .B(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(G127gat), .B(G155gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(G183gat), .B(G211gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(KEYINPUT77), .A2(KEYINPUT17), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT17), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n658_), .B2(new_n655_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n650_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n649_), .A2(new_n657_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(G229gat), .A2(G233gat), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n647_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n646_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n665_), .A2(new_n666_), .A3(new_n208_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n255_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n664_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n208_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n670_));
  OAI211_X1 g469(.A(new_n670_), .B(new_n663_), .C1(new_n210_), .C2(new_n648_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n669_), .A2(new_n671_), .A3(KEYINPUT79), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n210_), .A2(new_n648_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT79), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n673_), .A2(new_n670_), .A3(new_n674_), .A4(new_n663_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n672_), .A2(new_n675_), .ZN(new_n676_));
  XOR2_X1   g475(.A(G113gat), .B(G141gat), .Z(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT80), .ZN(new_n678_));
  XNOR2_X1  g477(.A(G169gat), .B(G197gat), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n678_), .B(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n676_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n672_), .A2(new_n675_), .A3(new_n680_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n634_), .A2(new_n662_), .A3(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n568_), .A2(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G1gat), .B1(new_n687_), .B2(new_n565_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT38), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n634_), .A2(new_n685_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n552_), .A2(new_n567_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(KEYINPUT75), .B(KEYINPUT37), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n694_), .B1(new_n273_), .B2(new_n278_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n267_), .A2(new_n272_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(new_n277_), .A3(new_n693_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n699_), .A2(new_n662_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n692_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n565_), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n703_), .A2(KEYINPUT102), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(KEYINPUT102), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  OR3_X1    g505(.A1(new_n702_), .A2(G1gat), .A3(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(new_n689_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n708_), .A2(KEYINPUT103), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n708_), .A2(KEYINPUT103), .ZN(new_n710_));
  OAI221_X1 g509(.A(new_n688_), .B1(new_n689_), .B2(new_n707_), .C1(new_n709_), .C2(new_n710_), .ZN(G1324gat));
  NAND2_X1  g510(.A1(new_n562_), .A2(new_n563_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n568_), .A2(new_n686_), .A3(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(G8gat), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT39), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n712_), .A2(G8gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(new_n702_), .B2(new_n717_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n718_), .B(new_n719_), .ZN(G1325gat));
  OAI21_X1  g519(.A(G15gat), .B1(new_n687_), .B2(new_n382_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n722_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n382_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n701_), .A2(new_n284_), .A3(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n723_), .A2(new_n724_), .A3(new_n726_), .ZN(G1326gat));
  INV_X1    g526(.A(new_n460_), .ZN(new_n728_));
  OAI21_X1  g527(.A(G22gat), .B1(new_n687_), .B2(new_n728_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT42), .Z(new_n730_));
  NOR3_X1   g529(.A1(new_n702_), .A2(G22gat), .A3(new_n728_), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1327gat));
  INV_X1    g531(.A(new_n662_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n279_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n692_), .A2(new_n734_), .ZN(new_n735_));
  OR3_X1    g534(.A1(new_n735_), .A2(G29gat), .A3(new_n565_), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n634_), .A2(new_n733_), .A3(new_n685_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n738_), .B1(new_n691_), .B2(new_n699_), .ZN(new_n739_));
  AOI211_X1 g538(.A(KEYINPUT43), .B(new_n698_), .C1(new_n552_), .C2(new_n567_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n737_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  OAI211_X1 g542(.A(KEYINPUT44), .B(new_n737_), .C1(new_n739_), .C2(new_n740_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n706_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n747_), .A2(KEYINPUT106), .A3(G29gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(KEYINPUT106), .B1(new_n747_), .B2(G29gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n736_), .B1(new_n748_), .B2(new_n749_), .ZN(G1328gat));
  NAND2_X1  g549(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n743_), .A2(new_n713_), .A3(new_n744_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(G36gat), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT107), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT107), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n752_), .A2(new_n755_), .A3(G36gat), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n758_));
  INV_X1    g557(.A(new_n735_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n712_), .A2(G36gat), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT45), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n759_), .A2(new_n763_), .A3(new_n760_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n758_), .B1(new_n762_), .B2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n751_), .B1(new_n757_), .B2(new_n765_), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n752_), .A2(new_n755_), .A3(G36gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n755_), .B1(new_n752_), .B2(G36gat), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n751_), .B(new_n765_), .C1(new_n767_), .C2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n766_), .A2(new_n770_), .ZN(G1329gat));
  NAND3_X1  g570(.A1(new_n745_), .A2(G43gat), .A3(new_n725_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n285_), .B1(new_n735_), .B2(new_n382_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g574(.A1(new_n735_), .A2(G50gat), .A3(new_n728_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n745_), .A2(KEYINPUT109), .A3(new_n460_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(G50gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT109), .B1(new_n745_), .B2(new_n460_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n776_), .B1(new_n778_), .B2(new_n779_), .ZN(G1331gat));
  AND3_X1   g579(.A1(new_n632_), .A2(KEYINPUT13), .A3(new_n628_), .ZN(new_n781_));
  AOI21_X1  g580(.A(KEYINPUT13), .B1(new_n632_), .B2(new_n628_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NOR3_X1   g582(.A1(new_n783_), .A2(new_n662_), .A3(new_n684_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n568_), .ZN(new_n785_));
  OAI21_X1  g584(.A(G57gat), .B1(new_n785_), .B2(new_n565_), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n691_), .A2(new_n685_), .A3(new_n634_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n700_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n746_), .A2(new_n583_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n786_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT110), .ZN(G1332gat));
  INV_X1    g590(.A(new_n788_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n792_), .A2(new_n581_), .A3(new_n713_), .ZN(new_n793_));
  OAI21_X1  g592(.A(G64gat), .B1(new_n785_), .B2(new_n712_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(KEYINPUT111), .B(KEYINPUT48), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n795_), .A2(new_n796_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n793_), .B1(new_n797_), .B2(new_n798_), .ZN(G1333gat));
  OAI21_X1  g598(.A(G71gat), .B1(new_n785_), .B2(new_n382_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(KEYINPUT49), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n792_), .A2(new_n295_), .A3(new_n725_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(G1334gat));
  OAI21_X1  g602(.A(G78gat), .B1(new_n785_), .B2(new_n728_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT50), .ZN(new_n805_));
  OR2_X1    g604(.A1(new_n728_), .A2(G78gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n788_), .B2(new_n806_), .ZN(G1335gat));
  OR2_X1    g606(.A1(new_n739_), .A2(new_n740_), .ZN(new_n808_));
  NOR3_X1   g607(.A1(new_n783_), .A2(new_n733_), .A3(new_n684_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT112), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n810_), .A2(new_n813_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n812_), .A2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(G85gat), .B1(new_n815_), .B2(new_n565_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n787_), .A2(new_n734_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n818_), .A2(new_n215_), .A3(new_n746_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n816_), .A2(new_n819_), .ZN(G1336gat));
  OAI21_X1  g619(.A(G92gat), .B1(new_n815_), .B2(new_n712_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n818_), .A2(new_n216_), .A3(new_n713_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(G1337gat));
  NAND4_X1  g622(.A1(new_n818_), .A2(new_n211_), .A3(new_n213_), .A4(new_n725_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n382_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n825_), .B2(new_n224_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT51), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT51), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n828_), .B(new_n824_), .C1(new_n825_), .C2(new_n224_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n829_), .ZN(G1338gat));
  AOI21_X1  g629(.A(new_n212_), .B1(new_n811_), .B2(new_n460_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT52), .ZN(new_n832_));
  AND4_X1   g631(.A1(new_n212_), .A2(new_n787_), .A3(new_n460_), .A4(new_n734_), .ZN(new_n833_));
  XOR2_X1   g632(.A(new_n833_), .B(KEYINPUT113), .Z(new_n834_));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n831_), .A2(KEYINPUT52), .ZN(new_n836_));
  OAI21_X1  g635(.A(KEYINPUT53), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n836_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n838_), .A2(new_n839_), .A3(new_n832_), .A4(new_n834_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n837_), .A2(new_n840_), .ZN(G1339gat));
  XNOR2_X1  g640(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT114), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n684_), .A2(new_n662_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n843_), .B1(new_n783_), .B2(new_n844_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n630_), .A2(new_n843_), .A3(new_n633_), .A4(new_n844_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n698_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n842_), .B1(new_n845_), .B2(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n630_), .A2(new_n633_), .A3(new_n844_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT114), .ZN(new_n850_));
  INV_X1    g649(.A(new_n842_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n850_), .A2(new_n698_), .A3(new_n851_), .A4(new_n846_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n848_), .A2(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n663_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n670_), .B(new_n664_), .C1(new_n210_), .C2(new_n648_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n854_), .A2(new_n855_), .A3(new_n680_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(KEYINPUT119), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n682_), .B(new_n857_), .C1(new_n625_), .C2(new_n629_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n628_), .A2(new_n684_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n598_), .A2(new_n615_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n254_), .A2(KEYINPUT12), .A3(new_n589_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n623_), .A2(new_n862_), .A3(KEYINPUT55), .A4(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(KEYINPUT117), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT117), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n620_), .A2(new_n866_), .A3(KEYINPUT55), .A4(new_n623_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT55), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n588_), .B1(new_n252_), .B2(new_n238_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n863_), .B1(new_n869_), .B2(new_n616_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n868_), .B1(new_n870_), .B2(new_n622_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n603_), .A2(new_n604_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n609_), .B1(new_n870_), .B2(new_n872_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n865_), .A2(new_n867_), .A3(new_n871_), .A4(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(KEYINPUT56), .B1(new_n874_), .B2(new_n575_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT118), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n628_), .A2(new_n684_), .A3(KEYINPUT116), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n861_), .A2(new_n876_), .A3(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n874_), .A2(new_n575_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT56), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n874_), .A2(KEYINPUT56), .A3(new_n575_), .ZN(new_n883_));
  AND3_X1   g682(.A1(new_n881_), .A2(new_n882_), .A3(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n858_), .B1(new_n878_), .B2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n279_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT57), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n881_), .A2(new_n882_), .A3(new_n883_), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n889_), .A2(new_n876_), .A3(new_n877_), .A4(new_n861_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n280_), .B1(new_n890_), .B2(new_n858_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT57), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n628_), .A2(new_n682_), .A3(new_n857_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n883_), .B1(new_n875_), .B2(KEYINPUT120), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n895_));
  AOI211_X1 g694(.A(new_n895_), .B(KEYINPUT56), .C1(new_n874_), .C2(new_n575_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n893_), .B1(new_n894_), .B2(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT58), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  OAI211_X1 g698(.A(KEYINPUT58), .B(new_n893_), .C1(new_n894_), .C2(new_n896_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n899_), .A2(new_n699_), .A3(new_n900_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n888_), .A2(new_n892_), .A3(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n853_), .B1(new_n902_), .B2(new_n662_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n746_), .A2(new_n725_), .A3(new_n564_), .ZN(new_n904_));
  OAI21_X1  g703(.A(KEYINPUT121), .B1(new_n903_), .B2(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n906_));
  INV_X1    g705(.A(new_n904_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n698_), .B1(new_n897_), .B2(new_n898_), .ZN(new_n908_));
  AOI22_X1  g707(.A1(new_n886_), .A2(new_n887_), .B1(new_n908_), .B2(new_n900_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n733_), .B1(new_n909_), .B2(new_n892_), .ZN(new_n910_));
  OAI211_X1 g709(.A(new_n906_), .B(new_n907_), .C1(new_n910_), .C2(new_n853_), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n905_), .A2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(G113gat), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n912_), .A2(new_n913_), .A3(new_n684_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n901_), .B1(KEYINPUT57), .B2(new_n891_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n886_), .A2(new_n887_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n662_), .B1(new_n915_), .B2(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n853_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n919_), .A2(KEYINPUT59), .A3(new_n907_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n921_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n685_), .B1(new_n920_), .B2(new_n922_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n914_), .B1(new_n913_), .B2(new_n923_), .ZN(G1340gat));
  INV_X1    g723(.A(G120gat), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n925_), .B1(new_n783_), .B2(KEYINPUT60), .ZN(new_n926_));
  OAI211_X1 g725(.A(new_n912_), .B(new_n926_), .C1(KEYINPUT60), .C2(new_n925_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n783_), .B1(new_n920_), .B2(new_n922_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n927_), .B1(new_n925_), .B2(new_n928_), .ZN(G1341gat));
  AOI211_X1 g728(.A(new_n355_), .B(new_n662_), .C1(new_n920_), .C2(new_n922_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n905_), .A2(new_n733_), .A3(new_n911_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(new_n355_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(KEYINPUT122), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n931_), .A2(new_n934_), .A3(new_n355_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n930_), .B1(new_n933_), .B2(new_n935_), .ZN(G1342gat));
  NAND3_X1  g735(.A1(new_n912_), .A2(new_n353_), .A3(new_n280_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n698_), .B1(new_n920_), .B2(new_n922_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n353_), .B2(new_n938_), .ZN(G1343gat));
  NOR4_X1   g738(.A1(new_n706_), .A2(new_n713_), .A3(new_n728_), .A4(new_n725_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(KEYINPUT123), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n903_), .A2(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n942_), .A2(new_n684_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g743(.A1(new_n942_), .A2(new_n634_), .ZN(new_n945_));
  XOR2_X1   g744(.A(KEYINPUT124), .B(G148gat), .Z(new_n946_));
  XNOR2_X1  g745(.A(new_n945_), .B(new_n946_), .ZN(G1345gat));
  NAND2_X1  g746(.A1(new_n942_), .A2(new_n733_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(KEYINPUT61), .B(G155gat), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n948_), .B(new_n949_), .ZN(G1346gat));
  INV_X1    g749(.A(G162gat), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n942_), .A2(new_n951_), .A3(new_n280_), .ZN(new_n952_));
  NOR3_X1   g751(.A1(new_n903_), .A2(new_n698_), .A3(new_n941_), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n952_), .B1(new_n951_), .B2(new_n953_), .ZN(G1347gat));
  NAND4_X1  g753(.A1(new_n706_), .A2(new_n728_), .A3(new_n725_), .A4(new_n713_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n955_), .B1(new_n917_), .B2(new_n918_), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n956_), .A2(new_n684_), .A3(new_n480_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n307_), .B1(KEYINPUT125), .B2(KEYINPUT62), .ZN(new_n958_));
  INV_X1    g757(.A(new_n958_), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n959_), .B1(new_n956_), .B2(new_n684_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n961_));
  INV_X1    g760(.A(new_n961_), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n957_), .B1(new_n960_), .B2(new_n962_), .ZN(new_n963_));
  AOI211_X1 g762(.A(new_n959_), .B(new_n961_), .C1(new_n956_), .C2(new_n684_), .ZN(new_n964_));
  OAI21_X1  g763(.A(KEYINPUT126), .B1(new_n963_), .B2(new_n964_), .ZN(new_n965_));
  INV_X1    g764(.A(new_n955_), .ZN(new_n966_));
  NAND3_X1  g765(.A1(new_n919_), .A2(new_n684_), .A3(new_n966_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n967_), .A2(new_n958_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n968_), .A2(new_n961_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n960_), .A2(new_n962_), .ZN(new_n970_));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n971_));
  NAND4_X1  g770(.A1(new_n969_), .A2(new_n970_), .A3(new_n971_), .A4(new_n957_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n965_), .A2(new_n972_), .ZN(G1348gat));
  NAND2_X1  g772(.A1(new_n956_), .A2(new_n634_), .ZN(new_n974_));
  XNOR2_X1  g773(.A(new_n974_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g774(.A1(new_n956_), .A2(new_n733_), .ZN(new_n976_));
  MUX2_X1   g775(.A(new_n320_), .B(G183gat), .S(new_n976_), .Z(G1350gat));
  INV_X1    g776(.A(new_n956_), .ZN(new_n978_));
  OAI21_X1  g777(.A(G190gat), .B1(new_n978_), .B2(new_n698_), .ZN(new_n979_));
  OAI21_X1  g778(.A(new_n280_), .B1(new_n471_), .B2(new_n470_), .ZN(new_n980_));
  OAI21_X1  g779(.A(new_n979_), .B1(new_n978_), .B2(new_n980_), .ZN(G1351gat));
  NOR4_X1   g780(.A1(new_n903_), .A2(new_n544_), .A3(new_n725_), .A4(new_n712_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n982_), .A2(new_n684_), .ZN(new_n983_));
  XNOR2_X1  g782(.A(new_n983_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g783(.A1(new_n982_), .A2(new_n634_), .ZN(new_n985_));
  XNOR2_X1  g784(.A(new_n985_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g785(.A1(new_n982_), .A2(new_n733_), .ZN(new_n987_));
  XNOR2_X1  g786(.A(KEYINPUT63), .B(G211gat), .ZN(new_n988_));
  NOR2_X1   g787(.A1(new_n987_), .A2(new_n988_), .ZN(new_n989_));
  NOR2_X1   g788(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n990_));
  AOI21_X1  g789(.A(new_n989_), .B1(new_n987_), .B2(new_n990_), .ZN(G1354gat));
  NAND2_X1  g790(.A1(new_n982_), .A2(new_n280_), .ZN(new_n992_));
  XOR2_X1   g791(.A(KEYINPUT127), .B(G218gat), .Z(new_n993_));
  NOR2_X1   g792(.A1(new_n698_), .A2(new_n993_), .ZN(new_n994_));
  AOI22_X1  g793(.A1(new_n992_), .A2(new_n993_), .B1(new_n982_), .B2(new_n994_), .ZN(G1355gat));
endmodule


