//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n706_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n815_, new_n816_, new_n817_, new_n818_, new_n820_,
    new_n821_, new_n822_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n829_, new_n830_, new_n831_, new_n833_, new_n834_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT19), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G183gat), .A2(G190gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT23), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT84), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT84), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n205_), .A2(new_n208_), .A3(KEYINPUT23), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n205_), .A2(KEYINPUT23), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n207_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT22), .B(G169gat), .ZN(new_n216_));
  INV_X1    g015(.A(G176gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n214_), .A2(new_n215_), .A3(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT25), .B(G183gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT26), .B(G190gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224_));
  AOI22_X1  g023(.A1(new_n221_), .A2(new_n222_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n215_), .A2(KEYINPUT24), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n226_), .A2(new_n224_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n210_), .A2(KEYINPUT86), .A3(new_n206_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT86), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n205_), .A2(new_n230_), .A3(KEYINPUT23), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n228_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT93), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT93), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n235_), .B1(new_n228_), .B2(new_n232_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n220_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(G197gat), .A2(G204gat), .ZN(new_n238_));
  INV_X1    g037(.A(G204gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT91), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT91), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(G204gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n238_), .B1(new_n243_), .B2(G197gat), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n244_), .A2(KEYINPUT21), .ZN(new_n245_));
  XOR2_X1   g044(.A(G211gat), .B(G218gat), .Z(new_n246_));
  OR2_X1    g045(.A1(new_n243_), .A2(G197gat), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT21), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n248_), .B1(G197gat), .B2(G204gat), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n246_), .B1(new_n247_), .B2(new_n249_), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n246_), .A2(KEYINPUT21), .ZN(new_n251_));
  AOI22_X1  g050(.A1(new_n245_), .A2(new_n250_), .B1(new_n244_), .B2(new_n251_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n237_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n218_), .A2(KEYINPUT85), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT85), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n216_), .A2(new_n255_), .A3(new_n217_), .ZN(new_n256_));
  AOI22_X1  g055(.A1(new_n254_), .A2(new_n256_), .B1(G169gat), .B2(G176gat), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n229_), .A2(new_n213_), .A3(new_n231_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n228_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(new_n211_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n245_), .A2(new_n250_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n251_), .A2(new_n244_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT20), .B1(new_n262_), .B2(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n204_), .B1(new_n253_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n237_), .A2(new_n252_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n204_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT20), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n270_), .B1(new_n262_), .B2(new_n265_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n268_), .A2(new_n269_), .A3(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(G8gat), .B(G36gat), .Z(new_n273_));
  XNOR2_X1  g072(.A(G64gat), .B(G92gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n267_), .A2(new_n272_), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT96), .ZN(new_n280_));
  NOR3_X1   g079(.A1(new_n265_), .A2(new_n220_), .A3(new_n233_), .ZN(new_n281_));
  AOI22_X1  g080(.A1(new_n257_), .A2(new_n258_), .B1(new_n260_), .B2(new_n211_), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT20), .B1(new_n282_), .B2(new_n252_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n204_), .B1(new_n281_), .B2(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n270_), .B1(new_n282_), .B2(new_n252_), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n285_), .B(new_n269_), .C1(new_n237_), .C2(new_n252_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  AOI22_X1  g086(.A1(new_n279_), .A2(new_n280_), .B1(new_n287_), .B2(new_n277_), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n267_), .A2(new_n272_), .A3(KEYINPUT96), .A4(new_n278_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n202_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n267_), .A2(new_n272_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(new_n277_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n292_), .A2(new_n202_), .A3(new_n279_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n290_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G227gat), .A2(G233gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(G15gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT30), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n282_), .B(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G127gat), .B(G134gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G113gat), .B(G120gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT87), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n299_), .B(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G71gat), .B(G99gat), .ZN(new_n305_));
  INV_X1    g104(.A(G43gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT31), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n304_), .A2(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n304_), .A2(new_n308_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(G141gat), .ZN(new_n313_));
  INV_X1    g112(.A(G148gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT88), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n315_), .B1(new_n316_), .B2(KEYINPUT3), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G141gat), .A2(G148gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT89), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT2), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT2), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n318_), .A2(KEYINPUT89), .A3(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT3), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n323_), .A2(new_n313_), .A3(new_n314_), .A4(KEYINPUT88), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n317_), .A2(new_n320_), .A3(new_n322_), .A4(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(G155gat), .B(G162gat), .Z(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT1), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n329_), .A2(new_n330_), .A3(new_n315_), .A4(new_n318_), .ZN(new_n331_));
  AND2_X1   g130(.A1(new_n327_), .A2(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n303_), .A2(new_n332_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n332_), .A2(new_n302_), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT4), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G225gat), .A2(G233gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT95), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT4), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(new_n303_), .B2(new_n332_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n335_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n340_));
  OR2_X1    g139(.A1(new_n333_), .A2(new_n334_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n337_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G1gat), .B(G29gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(G85gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT0), .B(G57gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n345_), .B(new_n346_), .Z(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n340_), .A2(new_n343_), .A3(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n348_), .B1(new_n340_), .B2(new_n343_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n327_), .A2(new_n331_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n252_), .B1(KEYINPUT29), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G228gat), .A2(G233gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  XOR2_X1   g157(.A(G22gat), .B(G50gat), .Z(new_n359_));
  INV_X1    g158(.A(KEYINPUT29), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n332_), .A2(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n362_));
  NOR2_X1   g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n354_), .A2(KEYINPUT29), .ZN(new_n364_));
  INV_X1    g163(.A(new_n362_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n359_), .B1(new_n363_), .B2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G78gat), .B(G106gat), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n369_), .A2(KEYINPUT92), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n361_), .A2(new_n362_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n359_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n364_), .A2(new_n365_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n371_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n367_), .A2(new_n370_), .A3(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n369_), .B1(new_n367_), .B2(new_n374_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n358_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n374_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n372_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n368_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n367_), .A2(new_n370_), .A3(new_n374_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n380_), .A2(new_n357_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n377_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NOR4_X1   g183(.A1(new_n295_), .A2(new_n312_), .A3(new_n353_), .A4(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n340_), .A2(new_n343_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(new_n347_), .ZN(new_n387_));
  AND4_X1   g186(.A1(new_n377_), .A2(new_n387_), .A3(new_n382_), .A4(new_n349_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n388_), .B1(new_n290_), .B2(new_n294_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT97), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n287_), .A2(KEYINPUT32), .A3(new_n278_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n278_), .A2(KEYINPUT32), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n267_), .A2(new_n272_), .A3(new_n393_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n392_), .B(new_n394_), .C1(new_n350_), .C2(new_n351_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT33), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n396_), .B1(new_n386_), .B2(new_n347_), .ZN(new_n397_));
  AOI211_X1 g196(.A(KEYINPUT33), .B(new_n348_), .C1(new_n340_), .C2(new_n343_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n337_), .B1(new_n335_), .B2(new_n339_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n348_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n292_), .B(new_n279_), .C1(new_n400_), .C2(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n395_), .B1(new_n399_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(new_n383_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n388_), .B(KEYINPUT97), .C1(new_n290_), .C2(new_n294_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n391_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n385_), .B1(new_n406_), .B2(new_n312_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G15gat), .B(G22gat), .ZN(new_n408_));
  INV_X1    g207(.A(G1gat), .ZN(new_n409_));
  INV_X1    g208(.A(G8gat), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT14), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n408_), .A2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G1gat), .B(G8gat), .ZN(new_n413_));
  XOR2_X1   g212(.A(new_n412_), .B(new_n413_), .Z(new_n414_));
  XNOR2_X1  g213(.A(G29gat), .B(G36gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT74), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G43gat), .B(G50gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT15), .ZN(new_n419_));
  INV_X1    g218(.A(new_n417_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n416_), .B(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT15), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n414_), .B1(new_n419_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G229gat), .A2(G233gat), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n418_), .A2(new_n414_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NOR3_X1   g227(.A1(new_n424_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT83), .ZN(new_n430_));
  INV_X1    g229(.A(new_n414_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n421_), .A2(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n425_), .B1(new_n427_), .B2(new_n432_), .ZN(new_n433_));
  NOR3_X1   g232(.A1(new_n429_), .A2(new_n430_), .A3(new_n433_), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n429_), .A2(new_n430_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G113gat), .B(G141gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G169gat), .B(G197gat), .ZN(new_n437_));
  XOR2_X1   g236(.A(new_n436_), .B(new_n437_), .Z(new_n438_));
  OR3_X1    g237(.A1(new_n434_), .A2(new_n435_), .A3(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n438_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n407_), .A2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT98), .ZN(new_n444_));
  INV_X1    g243(.A(G230gat), .ZN(new_n445_));
  INV_X1    g244(.A(G233gat), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT66), .ZN(new_n448_));
  OAI22_X1  g247(.A1(new_n448_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT7), .ZN(new_n450_));
  INV_X1    g249(.A(G99gat), .ZN(new_n451_));
  INV_X1    g250(.A(G106gat), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .A4(KEYINPUT66), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT6), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n454_), .B1(G99gat), .B2(G106gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G99gat), .A2(G106gat), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n456_), .A2(KEYINPUT6), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n449_), .B(new_n453_), .C1(new_n455_), .C2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT8), .ZN(new_n459_));
  AND2_X1   g258(.A1(G85gat), .A2(G92gat), .ZN(new_n460_));
  NOR2_X1   g259(.A1(G85gat), .A2(G92gat), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n458_), .A2(new_n459_), .A3(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n459_), .B1(new_n458_), .B2(new_n462_), .ZN(new_n464_));
  AND2_X1   g263(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n465_));
  NOR2_X1   g264(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n456_), .A2(KEYINPUT6), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n454_), .A2(G99gat), .A3(G106gat), .ZN(new_n469_));
  AOI22_X1  g268(.A1(new_n467_), .A2(new_n452_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT9), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n471_), .A2(G85gat), .A3(G92gat), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT64), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT9), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n471_), .A2(KEYINPUT64), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n472_), .B1(new_n476_), .B2(new_n462_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n470_), .B1(new_n477_), .B2(KEYINPUT65), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT65), .ZN(new_n479_));
  AOI211_X1 g278(.A(new_n479_), .B(new_n472_), .C1(new_n476_), .C2(new_n462_), .ZN(new_n480_));
  OAI22_X1  g279(.A1(new_n463_), .A2(new_n464_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT67), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n455_), .A2(new_n457_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n453_), .A2(new_n449_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n462_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT8), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n458_), .A2(new_n459_), .A3(new_n462_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G85gat), .B(G92gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n479_), .B1(new_n492_), .B2(new_n472_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n477_), .A2(KEYINPUT65), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(new_n494_), .A3(new_n470_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n489_), .A2(KEYINPUT67), .A3(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT68), .B(G71gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(G78gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G57gat), .B(G64gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT11), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n499_), .A2(KEYINPUT11), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n498_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(G78gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n497_), .B(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(new_n500_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n503_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n483_), .A2(new_n496_), .A3(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT69), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n508_), .B1(new_n483_), .B2(new_n496_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n447_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT70), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n481_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n489_), .A2(KEYINPUT70), .A3(new_n495_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n514_), .A2(KEYINPUT12), .A3(new_n507_), .A4(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n516_), .B1(new_n511_), .B2(KEYINPUT12), .ZN(new_n517_));
  INV_X1    g316(.A(new_n447_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n509_), .A2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT71), .B1(new_n517_), .B2(new_n519_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n509_), .A2(new_n518_), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n489_), .A2(KEYINPUT67), .A3(new_n495_), .ZN(new_n522_));
  AOI21_X1  g321(.A(KEYINPUT67), .B1(new_n489_), .B2(new_n495_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n507_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT12), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT71), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n521_), .A2(new_n526_), .A3(new_n527_), .A4(new_n516_), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n512_), .A2(new_n520_), .A3(new_n528_), .ZN(new_n529_));
  XOR2_X1   g328(.A(G176gat), .B(G204gat), .Z(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT73), .ZN(new_n531_));
  XOR2_X1   g330(.A(G120gat), .B(G148gat), .Z(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n533_), .B(new_n534_), .Z(new_n535_));
  OR2_X1    g334(.A1(new_n529_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n529_), .A2(new_n535_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n538_), .A2(KEYINPUT13), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(KEYINPUT13), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n421_), .A2(new_n422_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n418_), .A2(KEYINPUT15), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n514_), .B(new_n515_), .C1(new_n542_), .C2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n483_), .A2(new_n418_), .A3(new_n496_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT75), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G232gat), .A2(G233gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n548_), .B(new_n551_), .C1(KEYINPUT35), .C2(new_n546_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n551_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n546_), .A2(new_n547_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT79), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n552_), .A2(KEYINPUT79), .A3(new_n554_), .ZN(new_n558_));
  XOR2_X1   g357(.A(G190gat), .B(G218gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(G134gat), .B(G162gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT36), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n557_), .A2(new_n558_), .A3(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT76), .B(KEYINPUT36), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT77), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n552_), .A2(new_n554_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT78), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT78), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n552_), .A2(new_n569_), .A3(new_n554_), .A4(new_n566_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n563_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT37), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n573_), .B1(new_n555_), .B2(new_n562_), .ZN(new_n574_));
  AOI22_X1  g373(.A1(new_n572_), .A2(new_n573_), .B1(new_n571_), .B2(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(G127gat), .B(G155gat), .Z(new_n576_));
  XNOR2_X1  g375(.A(G183gat), .B(G211gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT17), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT81), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(new_n431_), .ZN(new_n583_));
  AND2_X1   g382(.A1(G231gat), .A2(G233gat), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n584_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(new_n508_), .A3(new_n586_), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n580_), .A2(KEYINPUT17), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT82), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n508_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n591_));
  OR3_X1    g390(.A1(new_n589_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n590_), .B1(new_n589_), .B2(new_n591_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n541_), .A2(new_n575_), .A3(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n444_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n597_), .A2(new_n409_), .A3(new_n353_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT38), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n562_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n601_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n602_));
  AOI22_X1  g401(.A1(new_n558_), .A2(new_n602_), .B1(new_n568_), .B2(new_n570_), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n407_), .A2(new_n594_), .A3(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n442_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(G1gat), .B1(new_n606_), .B2(new_n352_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n598_), .A2(new_n599_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n600_), .A2(new_n607_), .A3(new_n608_), .ZN(G1324gat));
  NAND3_X1  g408(.A1(new_n597_), .A2(new_n410_), .A3(new_n295_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n295_), .ZN(new_n611_));
  OAI21_X1  g410(.A(G8gat), .B1(new_n606_), .B2(new_n611_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n612_), .A2(KEYINPUT39), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(KEYINPUT39), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n610_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g415(.A(G15gat), .B1(new_n606_), .B2(new_n312_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT41), .Z(new_n618_));
  INV_X1    g417(.A(G15gat), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n597_), .A2(new_n619_), .A3(new_n311_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(G1326gat));
  OAI21_X1  g420(.A(G22gat), .B1(new_n606_), .B2(new_n383_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT42), .ZN(new_n623_));
  INV_X1    g422(.A(G22gat), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n597_), .A2(new_n624_), .A3(new_n384_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(G1327gat));
  NOR2_X1   g425(.A1(new_n595_), .A2(new_n572_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n627_), .A2(new_n541_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n444_), .A2(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(G29gat), .B1(new_n629_), .B2(new_n353_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT100), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT43), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n632_), .B1(new_n407_), .B2(new_n575_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n571_), .A2(new_n574_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n634_), .B1(new_n603_), .B2(KEYINPUT37), .ZN(new_n635_));
  AOI22_X1  g434(.A1(new_n389_), .A2(new_n390_), .B1(new_n403_), .B2(new_n383_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n311_), .B1(new_n636_), .B2(new_n405_), .ZN(new_n637_));
  OAI211_X1 g436(.A(KEYINPUT43), .B(new_n635_), .C1(new_n637_), .C2(new_n385_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n633_), .A2(new_n638_), .A3(new_n594_), .A4(new_n605_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT99), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n631_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT44), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(KEYINPUT99), .B1(new_n642_), .B2(KEYINPUT100), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n639_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n353_), .A2(G29gat), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n630_), .B1(new_n646_), .B2(new_n647_), .ZN(G1328gat));
  NOR2_X1   g447(.A1(new_n611_), .A2(G36gat), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n629_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(KEYINPUT45), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT45), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n629_), .A2(new_n652_), .A3(new_n649_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT101), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n635_), .B1(new_n637_), .B2(new_n385_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n595_), .B1(new_n656_), .B2(new_n632_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n657_), .A2(KEYINPUT99), .A3(new_n605_), .A4(new_n638_), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT44), .B1(new_n658_), .B2(new_n631_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n645_), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n655_), .B(new_n295_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(G36gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n655_), .B1(new_n646_), .B2(new_n295_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n654_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT46), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n654_), .B(KEYINPUT46), .C1(new_n662_), .C2(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1329gat));
  NAND3_X1  g467(.A1(new_n629_), .A2(new_n306_), .A3(new_n311_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n312_), .B1(new_n643_), .B2(new_n645_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n669_), .B1(new_n670_), .B2(new_n306_), .ZN(new_n671_));
  XOR2_X1   g470(.A(KEYINPUT102), .B(KEYINPUT47), .Z(new_n672_));
  XNOR2_X1  g471(.A(new_n671_), .B(new_n672_), .ZN(G1330gat));
  AOI21_X1  g472(.A(G50gat), .B1(new_n629_), .B2(new_n384_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n384_), .A2(G50gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n646_), .B2(new_n675_), .ZN(G1331gat));
  NOR3_X1   g475(.A1(new_n407_), .A2(new_n541_), .A3(new_n441_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n677_), .A2(new_n595_), .A3(new_n575_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n678_), .A2(new_n352_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n541_), .A2(new_n441_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n604_), .A2(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G57gat), .B1(new_n352_), .B2(KEYINPUT103), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n682_), .B1(KEYINPUT103), .B2(G57gat), .ZN(new_n683_));
  OAI22_X1  g482(.A1(new_n679_), .A2(G57gat), .B1(new_n681_), .B2(new_n683_), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT104), .Z(G1332gat));
  OAI21_X1  g484(.A(G64gat), .B1(new_n681_), .B2(new_n611_), .ZN(new_n686_));
  XOR2_X1   g485(.A(KEYINPUT105), .B(KEYINPUT48), .Z(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n611_), .A2(G64gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(new_n678_), .B2(new_n689_), .ZN(G1333gat));
  OAI21_X1  g489(.A(G71gat), .B1(new_n681_), .B2(new_n312_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT49), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n312_), .A2(G71gat), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n692_), .B1(new_n678_), .B2(new_n693_), .ZN(G1334gat));
  OAI21_X1  g493(.A(G78gat), .B1(new_n681_), .B2(new_n383_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT50), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n384_), .A2(new_n504_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n696_), .B1(new_n678_), .B2(new_n697_), .ZN(G1335gat));
  NAND3_X1  g497(.A1(new_n657_), .A2(new_n638_), .A3(new_n680_), .ZN(new_n699_));
  OAI21_X1  g498(.A(G85gat), .B1(new_n699_), .B2(new_n352_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n677_), .A2(new_n627_), .ZN(new_n701_));
  OR3_X1    g500(.A1(new_n701_), .A2(G85gat), .A3(new_n352_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(G1336gat));
  OAI21_X1  g502(.A(G92gat), .B1(new_n699_), .B2(new_n611_), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n611_), .A2(G92gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n704_), .B1(new_n701_), .B2(new_n705_), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT106), .Z(G1337gat));
  INV_X1    g506(.A(new_n701_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n708_), .A2(new_n311_), .A3(new_n467_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n699_), .A2(new_n312_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n711_), .B2(G99gat), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n710_), .B(G99gat), .C1(new_n699_), .C2(new_n312_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n709_), .B1(new_n712_), .B2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g515(.A1(new_n708_), .A2(new_n452_), .A3(new_n384_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT52), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n699_), .A2(new_n383_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n719_), .B2(G106gat), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n718_), .B(G106gat), .C1(new_n699_), .C2(new_n383_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n717_), .B1(new_n720_), .B2(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g523(.A(KEYINPUT54), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n596_), .A2(new_n725_), .A3(new_n442_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n596_), .B2(new_n442_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT115), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n729_), .A2(KEYINPUT57), .ZN(new_n730_));
  OR3_X1    g529(.A1(new_n424_), .A2(KEYINPUT112), .A3(new_n428_), .ZN(new_n731_));
  OAI21_X1  g530(.A(KEYINPUT112), .B1(new_n424_), .B2(new_n428_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n731_), .A2(new_n426_), .A3(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT113), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n427_), .A2(new_n432_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n438_), .B1(new_n735_), .B2(new_n425_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n733_), .A2(new_n734_), .A3(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n440_), .A2(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n734_), .B1(new_n733_), .B2(new_n736_), .ZN(new_n739_));
  OAI21_X1  g538(.A(KEYINPUT114), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n739_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT114), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n741_), .A2(new_n440_), .A3(new_n742_), .A4(new_n737_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n740_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n538_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n441_), .A2(new_n537_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT56), .ZN(new_n748_));
  XOR2_X1   g547(.A(KEYINPUT108), .B(KEYINPUT55), .Z(new_n749_));
  NAND3_X1  g548(.A1(new_n520_), .A2(new_n528_), .A3(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT109), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n520_), .A2(new_n528_), .A3(new_n752_), .A4(new_n749_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n447_), .B1(new_n510_), .B2(new_n517_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n521_), .A2(new_n526_), .A3(KEYINPUT55), .A4(new_n516_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n754_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n757_), .B1(new_n751_), .B2(new_n753_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n535_), .B1(new_n762_), .B2(KEYINPUT110), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n748_), .B1(new_n761_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT111), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n747_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n761_), .A2(new_n763_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(new_n765_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n748_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n746_), .B1(new_n766_), .B2(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n730_), .B1(new_n770_), .B2(new_n603_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n746_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n754_), .A2(KEYINPUT110), .A3(new_n758_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n535_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n762_), .A2(KEYINPUT110), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n765_), .B(KEYINPUT56), .C1(new_n775_), .C2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n747_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT56), .B1(new_n767_), .B2(new_n765_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n772_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n730_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(new_n572_), .A3(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT58), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n761_), .A2(new_n763_), .A3(new_n748_), .ZN(new_n785_));
  AOI22_X1  g584(.A1(new_n740_), .A2(new_n743_), .B1(new_n529_), .B2(new_n535_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n784_), .B1(new_n787_), .B2(new_n764_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT116), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(new_n789_), .A3(new_n635_), .ZN(new_n790_));
  OR3_X1    g589(.A1(new_n787_), .A2(new_n784_), .A3(new_n764_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n789_), .B1(new_n788_), .B2(new_n635_), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n771_), .B(new_n783_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n728_), .B1(new_n794_), .B2(new_n594_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n295_), .A2(new_n384_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(new_n353_), .A3(new_n311_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n795_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(G113gat), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(new_n799_), .A3(new_n441_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n794_), .A2(new_n594_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n728_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n797_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n803_), .A2(KEYINPUT59), .A3(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT59), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n806_), .B1(new_n795_), .B2(new_n797_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n442_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n800_), .B1(new_n808_), .B2(new_n799_), .ZN(G1340gat));
  INV_X1    g608(.A(G120gat), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n810_), .B1(new_n541_), .B2(KEYINPUT60), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n798_), .B(new_n811_), .C1(KEYINPUT60), .C2(new_n810_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n541_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n812_), .B1(new_n813_), .B2(new_n810_), .ZN(G1341gat));
  AOI21_X1  g613(.A(G127gat), .B1(new_n798_), .B2(new_n595_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n805_), .A2(new_n807_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n595_), .A2(G127gat), .ZN(new_n817_));
  XOR2_X1   g616(.A(new_n817_), .B(KEYINPUT117), .Z(new_n818_));
  AOI21_X1  g617(.A(new_n815_), .B1(new_n816_), .B2(new_n818_), .ZN(G1342gat));
  INV_X1    g618(.A(G134gat), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n798_), .A2(new_n820_), .A3(new_n603_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n575_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n822_), .B2(new_n820_), .ZN(G1343gat));
  NOR4_X1   g622(.A1(new_n295_), .A2(new_n383_), .A3(new_n352_), .A4(new_n311_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n795_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n441_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g627(.A(new_n541_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n826_), .A2(new_n829_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(KEYINPUT118), .B(G148gat), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n830_), .B(new_n831_), .ZN(G1345gat));
  NAND2_X1  g631(.A1(new_n826_), .A2(new_n595_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(KEYINPUT61), .B(G155gat), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n833_), .B(new_n834_), .ZN(G1346gat));
  NAND2_X1  g634(.A1(new_n803_), .A2(new_n824_), .ZN(new_n836_));
  INV_X1    g635(.A(G162gat), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n836_), .A2(new_n837_), .A3(new_n575_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT119), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n795_), .A2(new_n572_), .A3(new_n825_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n840_), .B2(G162gat), .ZN(new_n841_));
  OAI211_X1 g640(.A(KEYINPUT119), .B(new_n837_), .C1(new_n836_), .C2(new_n572_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n838_), .B1(new_n841_), .B2(new_n842_), .ZN(G1347gat));
  NOR3_X1   g642(.A1(new_n611_), .A2(new_n353_), .A3(new_n312_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n441_), .ZN(new_n845_));
  XOR2_X1   g644(.A(new_n845_), .B(KEYINPUT120), .Z(new_n846_));
  NAND3_X1  g645(.A1(new_n803_), .A2(new_n383_), .A3(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT62), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n847_), .A2(new_n848_), .A3(G169gat), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n848_), .B1(new_n847_), .B2(G169gat), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n803_), .A2(new_n383_), .A3(new_n844_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n441_), .A2(new_n216_), .ZN(new_n852_));
  OAI22_X1  g651(.A1(new_n849_), .A2(new_n850_), .B1(new_n851_), .B2(new_n852_), .ZN(G1348gat));
  NOR2_X1   g652(.A1(new_n795_), .A2(new_n384_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n854_), .A2(new_n829_), .A3(new_n844_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT121), .B(G176gat), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(G1349gat));
  NAND3_X1  g656(.A1(new_n854_), .A2(new_n595_), .A3(new_n844_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n859_), .B2(G183gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n221_), .B1(KEYINPUT122), .B2(G183gat), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n858_), .B2(new_n861_), .ZN(G1350gat));
  OAI21_X1  g661(.A(G190gat), .B1(new_n851_), .B2(new_n575_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n603_), .A2(new_n222_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n851_), .B2(new_n864_), .ZN(G1351gat));
  NAND3_X1  g664(.A1(new_n295_), .A2(new_n312_), .A3(new_n388_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n866_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n441_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g668(.A(new_n866_), .ZN(new_n870_));
  AOI21_X1  g669(.A(KEYINPUT111), .B1(new_n761_), .B2(new_n763_), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n777_), .B(new_n778_), .C1(KEYINPUT56), .C2(new_n871_), .ZN(new_n872_));
  AOI211_X1 g671(.A(new_n603_), .B(new_n730_), .C1(new_n872_), .C2(new_n772_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n782_), .B1(new_n781_), .B2(new_n572_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n788_), .A2(new_n635_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT116), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n877_), .A2(new_n791_), .A3(new_n790_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n595_), .B1(new_n875_), .B2(new_n878_), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n829_), .B(new_n870_), .C1(new_n879_), .C2(new_n728_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(KEYINPUT123), .A2(G204gat), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT124), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT123), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n240_), .B1(new_n242_), .B2(new_n884_), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n803_), .A2(new_n829_), .A3(new_n870_), .A4(new_n885_), .ZN(new_n886_));
  AND3_X1   g685(.A1(new_n882_), .A2(new_n883_), .A3(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n883_), .B1(new_n882_), .B2(new_n886_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1353gat));
  NAND2_X1  g688(.A1(new_n867_), .A2(new_n595_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(KEYINPUT63), .B(G211gat), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n892_), .B1(new_n890_), .B2(new_n893_), .ZN(G1354gat));
  AOI21_X1  g693(.A(G218gat), .B1(new_n867_), .B2(new_n603_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n635_), .A2(G218gat), .ZN(new_n896_));
  XOR2_X1   g695(.A(new_n896_), .B(KEYINPUT125), .Z(new_n897_));
  AND3_X1   g696(.A1(new_n803_), .A2(new_n870_), .A3(new_n897_), .ZN(new_n898_));
  OAI21_X1  g697(.A(KEYINPUT126), .B1(new_n895_), .B2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n867_), .A2(new_n897_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT126), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n795_), .A2(new_n572_), .A3(new_n866_), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n900_), .B(new_n901_), .C1(new_n902_), .C2(G218gat), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n899_), .A2(new_n903_), .ZN(G1355gat));
endmodule


