//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 0 0 1 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 1 1 0 0 0 0 1 1 1 1 0 1 1 0 0 1 1 1 1 0 1 0 0 0 0 1 0 0 0 0 0 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n792_, new_n793_, new_n794_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n899_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n927_, new_n928_, new_n930_,
    new_n931_, new_n933_, new_n934_, new_n936_, new_n937_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT86), .ZN(new_n204_));
  INV_X1    g003(.A(G197gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n204_), .B1(new_n205_), .B2(G204gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(G204gat), .ZN(new_n207_));
  INV_X1    g006(.A(G204gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n208_), .A2(KEYINPUT86), .A3(G197gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n206_), .A2(new_n207_), .A3(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT21), .ZN(new_n211_));
  INV_X1    g010(.A(G218gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(G211gat), .ZN(new_n213_));
  INV_X1    g012(.A(G211gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(G218gat), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n211_), .B1(new_n213_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n210_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT88), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT88), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n210_), .A2(new_n216_), .A3(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT87), .B(KEYINPUT21), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n222_), .A2(new_n206_), .A3(new_n207_), .A4(new_n209_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n213_), .A2(new_n215_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n208_), .A2(G197gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(new_n207_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n224_), .B1(KEYINPUT21), .B2(new_n226_), .ZN(new_n227_));
  AOI22_X1  g026(.A1(new_n218_), .A2(new_n220_), .B1(new_n223_), .B2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT25), .B(G183gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT26), .B(G190gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT24), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n231_), .B1(G169gat), .B2(G176gat), .ZN(new_n232_));
  INV_X1    g031(.A(G169gat), .ZN(new_n233_));
  INV_X1    g032(.A(G176gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  AOI22_X1  g034(.A1(new_n229_), .A2(new_n230_), .B1(new_n232_), .B2(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n231_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n240_));
  AND3_X1   g039(.A1(new_n238_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G169gat), .A2(G176gat), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT22), .B(G169gat), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n243_), .B1(new_n244_), .B2(new_n234_), .ZN(new_n245_));
  INV_X1    g044(.A(G183gat), .ZN(new_n246_));
  INV_X1    g045(.A(G190gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n238_), .A2(new_n248_), .A3(new_n239_), .ZN(new_n249_));
  AOI22_X1  g048(.A1(new_n236_), .A2(new_n241_), .B1(new_n245_), .B2(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT20), .B1(new_n228_), .B2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n226_), .A2(KEYINPUT21), .ZN(new_n252_));
  INV_X1    g051(.A(new_n224_), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n252_), .B(new_n253_), .C1(new_n210_), .C2(new_n221_), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n210_), .A2(new_n216_), .A3(new_n219_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n219_), .B1(new_n210_), .B2(new_n216_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n254_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n246_), .A2(KEYINPUT25), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT25), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(G183gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n247_), .A2(KEYINPUT26), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT26), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(G190gat), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n258_), .A2(new_n260_), .A3(new_n261_), .A4(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n239_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n265_), .A2(new_n237_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n235_), .A2(KEYINPUT24), .A3(new_n242_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n264_), .A2(new_n266_), .A3(new_n240_), .A4(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n233_), .A2(KEYINPUT22), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT22), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(G169gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n271_), .A3(new_n234_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n249_), .A2(new_n272_), .A3(new_n242_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n268_), .A2(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n257_), .A2(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n203_), .B1(new_n251_), .B2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G8gat), .B(G36gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT18), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G64gat), .B(G92gat), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n279_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT20), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n284_), .B1(new_n257_), .B2(new_n274_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n228_), .A2(new_n250_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n203_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n285_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n276_), .A2(new_n283_), .A3(new_n288_), .ZN(new_n289_));
  AND2_X1   g088(.A1(new_n289_), .A2(KEYINPUT27), .ZN(new_n290_));
  AND3_X1   g089(.A1(new_n285_), .A2(new_n287_), .A3(new_n286_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n274_), .A2(KEYINPUT98), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT98), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n268_), .A2(new_n273_), .A3(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n228_), .A2(new_n292_), .A3(new_n294_), .ZN(new_n295_));
  XOR2_X1   g094(.A(KEYINPUT97), .B(KEYINPUT20), .Z(new_n296_));
  AOI21_X1  g095(.A(new_n296_), .B1(new_n257_), .B2(new_n274_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n287_), .B1(new_n295_), .B2(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n282_), .B1(new_n291_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT100), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  OAI211_X1 g100(.A(KEYINPUT100), .B(new_n282_), .C1(new_n291_), .C2(new_n298_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n290_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT101), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT101), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n290_), .A2(new_n301_), .A3(new_n305_), .A4(new_n302_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(G50gat), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT28), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G155gat), .A2(G162gat), .ZN(new_n310_));
  OR2_X1    g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(KEYINPUT82), .A2(G141gat), .A3(G148gat), .ZN(new_n312_));
  AOI21_X1  g111(.A(KEYINPUT2), .B1(new_n312_), .B2(KEYINPUT85), .ZN(new_n313_));
  NAND2_X1  g112(.A1(KEYINPUT85), .A2(KEYINPUT2), .ZN(new_n314_));
  AOI22_X1  g113(.A1(new_n314_), .A2(KEYINPUT82), .B1(G141gat), .B2(G148gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(G141gat), .A2(G148gat), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT3), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n310_), .B(new_n311_), .C1(new_n316_), .C2(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321_));
  AND2_X1   g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT1), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n321_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  AND3_X1   g123(.A1(new_n310_), .A2(KEYINPUT83), .A3(KEYINPUT1), .ZN(new_n325_));
  AOI21_X1  g124(.A(KEYINPUT83), .B1(new_n310_), .B2(KEYINPUT1), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n324_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n312_), .ZN(new_n328_));
  AOI21_X1  g127(.A(KEYINPUT82), .B1(G141gat), .B2(G148gat), .ZN(new_n329_));
  NOR3_X1   g128(.A1(new_n328_), .A2(new_n329_), .A3(new_n317_), .ZN(new_n330_));
  AND3_X1   g129(.A1(new_n327_), .A2(KEYINPUT84), .A3(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(KEYINPUT84), .B1(new_n327_), .B2(new_n330_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n320_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n309_), .B1(new_n333_), .B2(KEYINPUT29), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n311_), .A2(new_n310_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G141gat), .A2(G148gat), .ZN(new_n336_));
  AND2_X1   g135(.A1(KEYINPUT85), .A2(KEYINPUT2), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT82), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n336_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n312_), .A2(KEYINPUT85), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n339_), .B1(new_n340_), .B2(KEYINPUT2), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n317_), .B(KEYINPUT3), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n335_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT84), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n323_), .A2(G155gat), .A3(G162gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(new_n311_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT83), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n347_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n310_), .A2(KEYINPUT83), .A3(KEYINPUT1), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n346_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  OR3_X1    g149(.A1(new_n328_), .A2(new_n329_), .A3(new_n317_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n344_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n327_), .A2(KEYINPUT84), .A3(new_n330_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n343_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT29), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(KEYINPUT28), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(G22gat), .ZN(new_n357_));
  AND3_X1   g156(.A1(new_n334_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n357_), .B1(new_n334_), .B2(new_n356_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n308_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n334_), .A2(new_n356_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(G22gat), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n334_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(G50gat), .A3(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n257_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G228gat), .A2(G233gat), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n257_), .B(new_n366_), .C1(new_n354_), .C2(new_n355_), .ZN(new_n369_));
  XOR2_X1   g168(.A(G78gat), .B(G106gat), .Z(new_n370_));
  NAND3_X1  g169(.A1(new_n368_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT89), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n360_), .A2(new_n364_), .A3(new_n373_), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n368_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n370_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n376_));
  OR2_X1    g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n374_), .A2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n375_), .A2(new_n376_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n379_), .A2(new_n360_), .A3(new_n373_), .A4(new_n364_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G1gat), .B(G29gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT91), .B(G85gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT0), .B(G57gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(G134gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(G127gat), .ZN(new_n388_));
  INV_X1    g187(.A(G127gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(G134gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(G120gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(G113gat), .ZN(new_n393_));
  INV_X1    g192(.A(G113gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(G120gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n391_), .A2(new_n396_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n388_), .A2(new_n390_), .A3(new_n393_), .A4(new_n395_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n333_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n352_), .A2(new_n353_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n397_), .A2(new_n398_), .A3(KEYINPUT90), .ZN(new_n403_));
  AOI21_X1  g202(.A(KEYINPUT90), .B1(new_n397_), .B2(new_n398_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n402_), .A2(new_n405_), .A3(new_n320_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G225gat), .A2(G233gat), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n401_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n401_), .A2(KEYINPUT4), .A3(new_n406_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n407_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n410_), .B1(new_n401_), .B2(KEYINPUT4), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n386_), .B(new_n408_), .C1(new_n409_), .C2(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n399_), .B1(new_n402_), .B2(new_n320_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT4), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n407_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n401_), .A2(KEYINPUT4), .A3(new_n406_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n386_), .B1(new_n417_), .B2(new_n408_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT99), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n412_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G227gat), .A2(G233gat), .ZN(new_n421_));
  INV_X1    g220(.A(G15gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT30), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G71gat), .B(G99gat), .ZN(new_n426_));
  INV_X1    g225(.A(G43gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n250_), .A2(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n274_), .A2(new_n428_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n425_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n250_), .A2(new_n429_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n274_), .A2(new_n428_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(new_n434_), .A3(new_n424_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n432_), .A2(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(KEYINPUT81), .B1(new_n436_), .B2(KEYINPUT80), .ZN(new_n437_));
  XOR2_X1   g236(.A(new_n399_), .B(KEYINPUT31), .Z(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n436_), .A2(KEYINPUT81), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n438_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n440_), .B1(new_n442_), .B2(new_n437_), .ZN(new_n443_));
  AOI211_X1 g242(.A(KEYINPUT99), .B(new_n386_), .C1(new_n417_), .C2(new_n408_), .ZN(new_n444_));
  NOR3_X1   g243(.A1(new_n420_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n287_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n282_), .B1(new_n291_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n289_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(KEYINPUT102), .B(KEYINPUT27), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT103), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n448_), .A2(KEYINPUT103), .A3(new_n449_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n307_), .A2(new_n381_), .A3(new_n445_), .A4(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT104), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n304_), .A2(new_n306_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT104), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n457_), .A2(new_n458_), .A3(new_n381_), .A4(new_n445_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n456_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT92), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n408_), .A2(new_n386_), .ZN(new_n462_));
  AOI211_X1 g261(.A(new_n461_), .B(KEYINPUT33), .C1(new_n462_), .C2(new_n417_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT33), .ZN(new_n464_));
  AOI21_X1  g263(.A(KEYINPUT92), .B1(new_n412_), .B2(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  NOR3_X1   g265(.A1(new_n291_), .A2(new_n446_), .A3(new_n282_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n283_), .B1(new_n276_), .B2(new_n288_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n462_), .A2(KEYINPUT33), .A3(new_n417_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT93), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n402_), .A2(new_n320_), .A3(new_n405_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n471_), .B1(new_n472_), .B2(new_n413_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n401_), .A2(KEYINPUT93), .A3(new_n406_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(new_n474_), .A3(new_n410_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n410_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n386_), .B1(new_n476_), .B2(new_n416_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n469_), .A2(new_n470_), .A3(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT94), .B1(new_n466_), .B2(new_n479_), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n469_), .A2(new_n470_), .A3(new_n478_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT94), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n481_), .B(new_n482_), .C1(new_n465_), .C2(new_n463_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n417_), .A2(new_n408_), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT99), .B1(new_n484_), .B2(new_n386_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n418_), .A2(new_n419_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(new_n486_), .A3(new_n412_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n291_), .A2(new_n446_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n280_), .A2(KEYINPUT32), .A3(new_n281_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT95), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT96), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT96), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n488_), .A2(new_n493_), .A3(new_n490_), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n291_), .A2(new_n298_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n489_), .ZN(new_n496_));
  AOI22_X1  g295(.A1(new_n492_), .A2(new_n494_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n487_), .A2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n480_), .A2(new_n483_), .A3(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n381_), .A2(new_n487_), .ZN(new_n500_));
  AOI22_X1  g299(.A1(new_n499_), .A2(new_n381_), .B1(new_n457_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n443_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n460_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT15), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G29gat), .B(G36gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT73), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G43gat), .B(G50gat), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT73), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n505_), .B(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n511_), .A2(new_n507_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n504_), .B1(new_n509_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n507_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n506_), .A2(new_n508_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(new_n515_), .A3(KEYINPUT15), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n513_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT76), .B(G1gat), .ZN(new_n518_));
  INV_X1    g317(.A(G8gat), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT14), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT77), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT75), .B(G15gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(new_n357_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G1gat), .B(G8gat), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n521_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n521_), .A2(new_n523_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n524_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n517_), .A2(new_n525_), .A3(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n509_), .A2(new_n512_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n525_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n524_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n530_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G229gat), .A2(G233gat), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n529_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT79), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n529_), .A2(new_n533_), .A3(KEYINPUT79), .A4(new_n534_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n534_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n528_), .A2(new_n525_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n540_), .A2(new_n530_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n530_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n542_), .B1(new_n528_), .B2(new_n525_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n539_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n537_), .A2(new_n538_), .A3(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G113gat), .B(G141gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G169gat), .B(G197gat), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n546_), .B(new_n547_), .Z(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n545_), .A2(new_n549_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n537_), .A2(new_n544_), .A3(new_n538_), .A4(new_n548_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n503_), .A2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(KEYINPUT10), .B(G99gat), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT65), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(G106gat), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G99gat), .A2(G106gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT6), .ZN(new_n560_));
  OAI21_X1  g359(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(KEYINPUT66), .B(G92gat), .ZN(new_n562_));
  INV_X1    g361(.A(G85gat), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n561_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT67), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n565_), .A2(new_n566_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n564_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n558_), .A2(new_n560_), .A3(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(KEYINPUT68), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT68), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n558_), .A2(new_n572_), .A3(new_n560_), .A4(new_n569_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n575_));
  OR3_X1    g374(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n560_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(G85gat), .B(G92gat), .Z(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT8), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT8), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n577_), .A2(new_n581_), .A3(new_n578_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n574_), .A2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G57gat), .B(G64gat), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n585_), .A2(KEYINPUT11), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(KEYINPUT11), .ZN(new_n587_));
  XOR2_X1   g386(.A(G71gat), .B(G78gat), .Z(new_n588_));
  NAND3_X1  g387(.A1(new_n586_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n587_), .A2(new_n588_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT12), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n584_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G230gat), .A2(G233gat), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n596_), .B(KEYINPUT64), .Z(new_n597_));
  NAND3_X1  g396(.A1(new_n583_), .A2(new_n570_), .A3(new_n591_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n591_), .B1(new_n583_), .B2(new_n570_), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n599_), .A2(KEYINPUT12), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n595_), .A2(new_n597_), .A3(new_n598_), .A4(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n599_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(new_n598_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n597_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  XOR2_X1   g404(.A(G120gat), .B(G148gat), .Z(new_n606_));
  XNOR2_X1  g405(.A(G176gat), .B(G204gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n601_), .A2(new_n605_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT71), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n601_), .A2(KEYINPUT71), .A3(new_n605_), .A4(new_n610_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n601_), .A2(new_n605_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n610_), .B(KEYINPUT70), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n615_), .A2(new_n618_), .A3(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n622_), .B1(new_n615_), .B2(new_n618_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G190gat), .B(G218gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G134gat), .B(G162gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT36), .Z(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  AOI22_X1  g429(.A1(new_n571_), .A2(new_n573_), .B1(new_n580_), .B2(new_n582_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n631_), .B1(new_n516_), .B2(new_n513_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n530_), .A2(new_n583_), .A3(new_n570_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(G232gat), .A2(G233gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT34), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n633_), .B1(KEYINPUT35), .B2(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n632_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(KEYINPUT35), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  OAI211_X1 g438(.A(KEYINPUT35), .B(new_n635_), .C1(new_n632_), .C2(new_n636_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n630_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n628_), .A2(KEYINPUT36), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n639_), .A2(new_n640_), .A3(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n642_), .A2(KEYINPUT37), .A3(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n641_), .A2(KEYINPUT74), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n644_), .B1(new_n641_), .B2(KEYINPUT74), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n645_), .B1(new_n648_), .B2(KEYINPUT37), .ZN(new_n649_));
  NAND2_X1  g448(.A1(G231gat), .A2(G233gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT78), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n540_), .B(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(new_n591_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(G127gat), .B(G155gat), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT16), .ZN(new_n655_));
  XOR2_X1   g454(.A(G183gat), .B(G211gat), .Z(new_n656_));
  XNOR2_X1  g455(.A(new_n655_), .B(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n653_), .A2(KEYINPUT17), .A3(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n657_), .B(KEYINPUT17), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n659_), .B1(new_n653_), .B2(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n649_), .A2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n553_), .A2(new_n625_), .A3(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(new_n487_), .A3(new_n518_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT38), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n552_), .B1(new_n621_), .B2(new_n623_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT105), .ZN(new_n670_));
  INV_X1    g469(.A(new_n662_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT105), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n672_), .B(new_n552_), .C1(new_n621_), .C2(new_n623_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n670_), .A2(new_n671_), .A3(new_n673_), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n674_), .A2(KEYINPUT106), .ZN(new_n675_));
  INV_X1    g474(.A(new_n648_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n503_), .A2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n674_), .A2(KEYINPUT106), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n675_), .A2(new_n677_), .A3(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n487_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G1gat), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n666_), .A2(new_n667_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n668_), .A2(new_n681_), .A3(new_n682_), .ZN(G1324gat));
  INV_X1    g482(.A(new_n457_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n665_), .A2(new_n519_), .A3(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G8gat), .B1(new_n679_), .B2(new_n457_), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n686_), .A2(KEYINPUT39), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n686_), .A2(KEYINPUT39), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n685_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT40), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  OAI211_X1 g491(.A(KEYINPUT40), .B(new_n685_), .C1(new_n688_), .C2(new_n689_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1325gat));
  OAI21_X1  g493(.A(G15gat), .B1(new_n679_), .B2(new_n443_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n696_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n665_), .A2(new_n422_), .A3(new_n502_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n697_), .A2(new_n698_), .A3(new_n699_), .ZN(G1326gat));
  OAI21_X1  g499(.A(G22gat), .B1(new_n679_), .B2(new_n381_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT42), .ZN(new_n702_));
  INV_X1    g501(.A(new_n381_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n665_), .A2(new_n357_), .A3(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(G1327gat));
  AND4_X1   g504(.A1(new_n553_), .A2(new_n625_), .A3(new_n662_), .A4(new_n648_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G29gat), .B1(new_n706_), .B2(new_n487_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT110), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n670_), .A2(new_n662_), .A3(new_n673_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n499_), .A2(new_n381_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n500_), .A2(new_n457_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n502_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n456_), .A2(new_n459_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n649_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  XOR2_X1   g513(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n503_), .A2(new_n717_), .A3(new_n649_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n709_), .B1(new_n716_), .B2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n708_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n709_), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n503_), .A2(new_n717_), .A3(new_n649_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n715_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n724_), .B1(new_n503_), .B2(new_n649_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n722_), .B1(new_n723_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n720_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n726_), .A2(KEYINPUT110), .A3(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n721_), .A2(new_n728_), .ZN(new_n729_));
  OAI211_X1 g528(.A(KEYINPUT44), .B(new_n722_), .C1(new_n723_), .C2(new_n725_), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n730_), .A2(G29gat), .A3(new_n487_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n707_), .B1(new_n729_), .B2(new_n731_), .ZN(G1328gat));
  INV_X1    g531(.A(G36gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n706_), .A2(new_n733_), .A3(new_n684_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT45), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n730_), .A2(new_n684_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n736_), .B1(new_n721_), .B2(new_n728_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT111), .ZN(new_n738_));
  OAI21_X1  g537(.A(G36gat), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  AOI211_X1 g538(.A(KEYINPUT111), .B(new_n736_), .C1(new_n721_), .C2(new_n728_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n735_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT46), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  OAI211_X1 g542(.A(KEYINPUT46), .B(new_n735_), .C1(new_n739_), .C2(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1329gat));
  AOI21_X1  g544(.A(G43gat), .B1(new_n706_), .B2(new_n502_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n730_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n747_), .A2(new_n427_), .A3(new_n443_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n746_), .B1(new_n748_), .B2(new_n729_), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g549(.A(G50gat), .B1(new_n706_), .B2(new_n703_), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n747_), .A2(new_n308_), .A3(new_n381_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n752_), .B2(new_n729_), .ZN(G1331gat));
  INV_X1    g552(.A(new_n552_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n503_), .A2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n755_), .A2(new_n624_), .A3(new_n663_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT112), .ZN(new_n757_));
  AOI21_X1  g556(.A(G57gat), .B1(new_n757_), .B2(new_n487_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n624_), .A2(new_n754_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n759_), .A2(new_n662_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n677_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n680_), .A2(KEYINPUT113), .ZN(new_n763_));
  MUX2_X1   g562(.A(KEYINPUT113), .B(new_n763_), .S(G57gat), .Z(new_n764_));
  AOI21_X1  g563(.A(new_n758_), .B1(new_n762_), .B2(new_n764_), .ZN(G1332gat));
  OAI21_X1  g564(.A(G64gat), .B1(new_n761_), .B2(new_n457_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT48), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n457_), .A2(G64gat), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT114), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n757_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n767_), .A2(new_n770_), .ZN(G1333gat));
  INV_X1    g570(.A(G71gat), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n757_), .A2(new_n772_), .A3(new_n502_), .ZN(new_n773_));
  OAI21_X1  g572(.A(G71gat), .B1(new_n761_), .B2(new_n443_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT49), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1334gat));
  INV_X1    g575(.A(G78gat), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n757_), .A2(new_n777_), .A3(new_n703_), .ZN(new_n778_));
  OAI21_X1  g577(.A(G78gat), .B1(new_n761_), .B2(new_n381_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT50), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(G1335gat));
  NAND4_X1  g580(.A1(new_n755_), .A2(new_n624_), .A3(new_n662_), .A4(new_n648_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n783_), .A2(new_n563_), .A3(new_n487_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n716_), .A2(new_n718_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n759_), .A2(new_n671_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n787_), .A2(KEYINPUT115), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(KEYINPUT115), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n680_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n784_), .B1(new_n790_), .B2(new_n563_), .ZN(G1336gat));
  AOI21_X1  g590(.A(G92gat), .B1(new_n783_), .B2(new_n684_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n788_), .A2(new_n789_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n457_), .A2(new_n562_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n792_), .B1(new_n793_), .B2(new_n794_), .ZN(G1337gat));
  NAND3_X1  g594(.A1(new_n783_), .A2(new_n502_), .A3(new_n556_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n443_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n797_));
  INV_X1    g596(.A(G99gat), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n796_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g599(.A1(new_n783_), .A2(new_n557_), .A3(new_n703_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802_));
  INV_X1    g601(.A(new_n787_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n703_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n802_), .B1(new_n804_), .B2(G106gat), .ZN(new_n805_));
  AOI211_X1 g604(.A(KEYINPUT52), .B(new_n557_), .C1(new_n803_), .C2(new_n703_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n801_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g607(.A1(new_n663_), .A2(new_n754_), .A3(new_n625_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT54), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n631_), .A2(new_n593_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n598_), .B1(new_n599_), .B2(KEYINPUT12), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n811_), .A2(new_n604_), .A3(new_n812_), .ZN(new_n813_));
  XOR2_X1   g612(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n814_));
  OAI21_X1  g613(.A(KEYINPUT118), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n597_), .A2(KEYINPUT119), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n595_), .A2(new_n598_), .A3(new_n600_), .A4(new_n816_), .ZN(new_n817_));
  OAI22_X1  g616(.A1(new_n811_), .A2(new_n812_), .B1(KEYINPUT119), .B2(new_n597_), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n604_), .A2(KEYINPUT55), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n817_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT118), .ZN(new_n821_));
  INV_X1    g620(.A(new_n814_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n601_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n815_), .A2(new_n820_), .A3(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n617_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT56), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT56), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n824_), .A2(new_n827_), .A3(new_n617_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT121), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n529_), .A2(new_n829_), .A3(new_n533_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n529_), .B2(new_n533_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n830_), .A2(new_n831_), .A3(new_n534_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n534_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n549_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n551_), .B1(new_n832_), .B2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n835_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n826_), .A2(new_n828_), .A3(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT58), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n826_), .A2(KEYINPUT58), .A3(new_n836_), .A4(new_n828_), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n839_), .A2(new_n649_), .A3(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT57), .ZN(new_n843_));
  AOI21_X1  g642(.A(KEYINPUT116), .B1(new_n615_), .B2(new_n552_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n846_), .B1(new_n824_), .B2(new_n617_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n615_), .A2(new_n552_), .A3(KEYINPUT116), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n824_), .A2(new_n617_), .A3(new_n846_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n845_), .A2(new_n848_), .A3(new_n849_), .A4(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n615_), .A2(new_n618_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n835_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n851_), .A2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n843_), .B1(new_n855_), .B2(new_n676_), .ZN(new_n856_));
  AOI211_X1 g655(.A(KEYINPUT57), .B(new_n648_), .C1(new_n851_), .C2(new_n854_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n842_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n662_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n810_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n861_));
  NOR4_X1   g660(.A1(new_n684_), .A2(new_n680_), .A3(new_n703_), .A4(new_n443_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n860_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n615_), .A2(new_n552_), .A3(KEYINPUT116), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n864_), .A2(new_n844_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n850_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n847_), .ZN(new_n867_));
  AOI22_X1  g666(.A1(new_n865_), .A2(new_n867_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n868_));
  OAI21_X1  g667(.A(KEYINPUT57), .B1(new_n868_), .B2(new_n648_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n855_), .A2(new_n843_), .A3(new_n676_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n841_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n662_), .B1(new_n871_), .B2(KEYINPUT122), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n842_), .B(KEYINPUT122), .C1(new_n856_), .C2(new_n857_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n810_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n875_), .A2(new_n862_), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n552_), .B(new_n863_), .C1(new_n876_), .C2(new_n861_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(G113gat), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n876_), .A2(new_n394_), .A3(new_n552_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1340gat));
  OAI211_X1 g679(.A(new_n624_), .B(new_n863_), .C1(new_n876_), .C2(new_n861_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(G120gat), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n392_), .B1(new_n625_), .B2(KEYINPUT60), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n876_), .B(new_n883_), .C1(KEYINPUT60), .C2(new_n392_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n882_), .A2(new_n884_), .ZN(G1341gat));
  OAI211_X1 g684(.A(new_n671_), .B(new_n863_), .C1(new_n876_), .C2(new_n861_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(G127gat), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n876_), .A2(new_n389_), .A3(new_n671_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1342gat));
  OAI211_X1 g688(.A(new_n649_), .B(new_n863_), .C1(new_n876_), .C2(new_n861_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(G134gat), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n876_), .A2(new_n387_), .A3(new_n648_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1343gat));
  NOR2_X1   g692(.A1(new_n381_), .A2(new_n502_), .ZN(new_n894_));
  AND2_X1   g693(.A1(new_n875_), .A2(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n684_), .A2(new_n680_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n895_), .A2(new_n552_), .A3(new_n896_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g697(.A1(new_n895_), .A2(new_n624_), .A3(new_n896_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g699(.A1(new_n895_), .A2(new_n671_), .A3(new_n896_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT61), .B(G155gat), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1346gat));
  NAND2_X1  g702(.A1(new_n895_), .A2(new_n896_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n649_), .ZN(new_n905_));
  OAI21_X1  g704(.A(G162gat), .B1(new_n904_), .B2(new_n905_), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n676_), .A2(G162gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n904_), .B2(new_n907_), .ZN(G1347gat));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n233_), .B1(new_n909_), .B2(KEYINPUT62), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n703_), .B1(new_n810_), .B2(new_n859_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n457_), .A2(new_n487_), .A3(new_n443_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n910_), .B1(new_n913_), .B2(new_n754_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n909_), .A2(KEYINPUT62), .ZN(new_n915_));
  OR2_X1    g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n913_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n917_), .A2(new_n244_), .A3(new_n552_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n914_), .A2(new_n915_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n916_), .A2(new_n918_), .A3(new_n919_), .ZN(G1348gat));
  AOI21_X1  g719(.A(G176gat), .B1(new_n917_), .B2(new_n624_), .ZN(new_n921_));
  AND2_X1   g720(.A1(new_n875_), .A2(new_n381_), .ZN(new_n922_));
  AND3_X1   g721(.A1(new_n624_), .A2(G176gat), .A3(new_n912_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n921_), .B1(new_n922_), .B2(new_n923_), .ZN(G1349gat));
  AND2_X1   g723(.A1(new_n912_), .A2(new_n671_), .ZN(new_n925_));
  AOI21_X1  g724(.A(G183gat), .B1(new_n922_), .B2(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n229_), .ZN(new_n927_));
  AND2_X1   g726(.A1(new_n925_), .A2(new_n927_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n926_), .B1(new_n911_), .B2(new_n928_), .ZN(G1350gat));
  OAI21_X1  g728(.A(G190gat), .B1(new_n913_), .B2(new_n905_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n648_), .A2(new_n230_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n930_), .B1(new_n913_), .B2(new_n931_), .ZN(G1351gat));
  NOR2_X1   g731(.A1(new_n457_), .A2(new_n487_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n895_), .A2(new_n552_), .A3(new_n933_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g734(.A1(new_n895_), .A2(new_n624_), .A3(new_n933_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(KEYINPUT125), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n936_), .B(new_n938_), .ZN(G1353gat));
  NAND4_X1  g738(.A1(new_n875_), .A2(new_n671_), .A3(new_n894_), .A4(new_n933_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(KEYINPUT63), .B(G211gat), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n940_), .A2(new_n941_), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT63), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n940_), .A2(new_n943_), .A3(new_n214_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT126), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(new_n946_));
  NAND4_X1  g745(.A1(new_n940_), .A2(KEYINPUT126), .A3(new_n943_), .A4(new_n214_), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n942_), .B1(new_n946_), .B2(new_n947_), .ZN(G1354gat));
  NAND4_X1  g747(.A1(new_n875_), .A2(new_n649_), .A3(new_n894_), .A4(new_n933_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n949_), .A2(G218gat), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n676_), .A2(G218gat), .ZN(new_n951_));
  NAND4_X1  g750(.A1(new_n875_), .A2(new_n894_), .A3(new_n933_), .A4(new_n951_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n950_), .A2(new_n952_), .ZN(new_n953_));
  INV_X1    g752(.A(KEYINPUT127), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n953_), .A2(new_n954_), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n950_), .A2(KEYINPUT127), .A3(new_n952_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n955_), .A2(new_n956_), .ZN(G1355gat));
endmodule


