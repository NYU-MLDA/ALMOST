//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 1 1 1 1 1 1 0 1 1 1 1 0 1 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n853_, new_n855_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n912_;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT8), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT6), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT66), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n204_), .B(KEYINPUT6), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT66), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  OR2_X1    g010(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n212_));
  NAND2_X1  g011(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n211_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  AND2_X1   g013(.A1(new_n211_), .A2(new_n213_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n208_), .A2(new_n210_), .A3(new_n216_), .ZN(new_n217_));
  XOR2_X1   g016(.A(G85gat), .B(G92gat), .Z(new_n218_));
  AOI21_X1  g017(.A(new_n203_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n203_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n220_), .B1(new_n216_), .B2(new_n209_), .ZN(new_n221_));
  OR2_X1    g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(KEYINPUT10), .B(G99gat), .Z(new_n223_));
  INV_X1    g022(.A(G106gat), .ZN(new_n224_));
  AOI22_X1  g023(.A1(KEYINPUT9), .A2(new_n218_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT64), .B(G85gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT9), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(new_n227_), .A3(G92gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n225_), .A2(new_n209_), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n222_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT67), .B(G71gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(G78gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G57gat), .B(G64gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT11), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n233_), .B(KEYINPUT11), .Z(new_n236_));
  OAI21_X1  g035(.A(new_n235_), .B1(new_n236_), .B2(new_n232_), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n230_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n230_), .A2(new_n237_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(KEYINPUT12), .A3(new_n239_), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n239_), .A2(KEYINPUT12), .ZN(new_n241_));
  AOI22_X1  g040(.A1(new_n240_), .A2(new_n241_), .B1(G230gat), .B2(G233gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G230gat), .A2(G233gat), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n243_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  XOR2_X1   g044(.A(G120gat), .B(G148gat), .Z(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G176gat), .B(G204gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n245_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT13), .ZN(new_n252_));
  INV_X1    g051(.A(new_n250_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n253_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n251_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n252_), .B1(new_n251_), .B2(new_n254_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n202_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n251_), .A2(new_n254_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT13), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n260_), .A2(KEYINPUT69), .A3(new_n255_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G1gat), .B(G8gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT74), .ZN(new_n264_));
  OR2_X1    g063(.A1(G15gat), .A2(G22gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G15gat), .A2(G22gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G1gat), .A2(G8gat), .ZN(new_n267_));
  AOI22_X1  g066(.A1(new_n265_), .A2(new_n266_), .B1(KEYINPUT14), .B2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n264_), .B(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G29gat), .B(G36gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G43gat), .B(G50gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n269_), .B(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G229gat), .A2(G233gat), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  XOR2_X1   g075(.A(new_n276_), .B(KEYINPUT77), .Z(new_n277_));
  XOR2_X1   g076(.A(new_n272_), .B(KEYINPUT15), .Z(new_n278_));
  NOR2_X1   g077(.A1(new_n278_), .A2(new_n269_), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n269_), .A2(new_n272_), .ZN(new_n280_));
  OR3_X1    g079(.A1(new_n279_), .A2(new_n280_), .A3(new_n275_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n277_), .A2(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(G113gat), .B(G141gat), .Z(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT78), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G169gat), .B(G197gat), .ZN(new_n285_));
  XOR2_X1   g084(.A(new_n284_), .B(new_n285_), .Z(new_n286_));
  NAND2_X1  g085(.A1(new_n282_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n286_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n277_), .A2(new_n281_), .A3(new_n288_), .ZN(new_n289_));
  AND3_X1   g088(.A1(new_n287_), .A2(KEYINPUT79), .A3(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(KEYINPUT79), .B1(new_n287_), .B2(new_n289_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n262_), .A2(new_n293_), .ZN(new_n294_));
  OR3_X1    g093(.A1(KEYINPUT89), .A2(G155gat), .A3(G162gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT89), .B1(G155gat), .B2(G162gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297_));
  AND3_X1   g096(.A1(new_n295_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(G141gat), .A2(G148gat), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT90), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT3), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT90), .B1(G141gat), .B2(G148gat), .ZN(new_n303_));
  AND3_X1   g102(.A1(new_n301_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G141gat), .A2(G148gat), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT91), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT2), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n309_));
  AOI21_X1  g108(.A(KEYINPUT91), .B1(G141gat), .B2(G148gat), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n308_), .B(new_n309_), .C1(new_n307_), .C2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n298_), .B1(new_n304_), .B2(new_n311_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n297_), .A2(KEYINPUT1), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n297_), .A2(KEYINPUT1), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n313_), .A2(new_n295_), .A3(new_n296_), .A4(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n305_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n316_), .A2(new_n299_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n312_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G127gat), .B(G134gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G113gat), .B(G120gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n319_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n301_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT2), .B1(new_n316_), .B2(KEYINPUT91), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n325_), .A2(new_n326_), .A3(new_n309_), .A4(new_n308_), .ZN(new_n327_));
  AOI22_X1  g126(.A1(new_n327_), .A2(new_n298_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(new_n322_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G225gat), .A2(G233gat), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n324_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G1gat), .B(G29gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(G85gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT0), .B(G57gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT33), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  AND3_X1   g136(.A1(new_n312_), .A2(new_n322_), .A3(new_n318_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n322_), .B1(new_n312_), .B2(new_n318_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT4), .ZN(new_n340_));
  NOR3_X1   g139(.A1(new_n338_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n319_), .A2(new_n340_), .A3(new_n323_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n330_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n331_), .B(new_n337_), .C1(new_n341_), .C2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT98), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n324_), .A2(new_n329_), .A3(KEYINPUT4), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n348_), .A2(new_n343_), .A3(new_n342_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n349_), .A2(KEYINPUT98), .A3(new_n331_), .A4(new_n337_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n347_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n335_), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n331_), .B(new_n352_), .C1(new_n341_), .C2(new_n344_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n348_), .A2(new_n330_), .A3(new_n342_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n338_), .A2(new_n339_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n352_), .B1(new_n355_), .B2(new_n343_), .ZN(new_n356_));
  AOI22_X1  g155(.A1(new_n353_), .A2(new_n336_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT80), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G169gat), .A2(G176gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT24), .ZN(new_n360_));
  NOR2_X1   g159(.A1(G169gat), .A2(G176gat), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n358_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(G183gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT25), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT25), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(G183gat), .ZN(new_n366_));
  INV_X1    g165(.A(G190gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT26), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT26), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(G190gat), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n364_), .A2(new_n366_), .A3(new_n368_), .A4(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(G169gat), .ZN(new_n372_));
  INV_X1    g171(.A(G176gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n374_), .A2(KEYINPUT80), .A3(KEYINPUT24), .A4(new_n359_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n362_), .A2(new_n371_), .A3(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT81), .ZN(new_n377_));
  AND3_X1   g176(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n378_));
  AOI21_X1  g177(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT24), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n381_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n382_));
  AOI21_X1  g181(.A(KEYINPUT82), .B1(new_n380_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G183gat), .A2(G190gat), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT23), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n387_));
  AND4_X1   g186(.A1(KEYINPUT82), .A2(new_n382_), .A3(new_n386_), .A4(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n383_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT81), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n362_), .A2(new_n371_), .A3(new_n390_), .A4(new_n375_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n377_), .A2(new_n389_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT21), .ZN(new_n393_));
  AND2_X1   g192(.A1(G197gat), .A2(G204gat), .ZN(new_n394_));
  NOR2_X1   g193(.A1(G197gat), .A2(G204gat), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n393_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT93), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  OAI211_X1 g197(.A(KEYINPUT93), .B(new_n393_), .C1(new_n394_), .C2(new_n395_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n394_), .A2(new_n395_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT21), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G211gat), .B(G218gat), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n398_), .A2(new_n399_), .A3(new_n401_), .A4(new_n402_), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n401_), .A2(new_n402_), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n386_), .B(new_n387_), .C1(G183gat), .C2(G190gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(KEYINPUT83), .A2(KEYINPUT22), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(G169gat), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n372_), .A2(KEYINPUT83), .A3(KEYINPUT22), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(new_n409_), .A3(new_n373_), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n410_), .A2(KEYINPUT84), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(KEYINPUT84), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n359_), .B(new_n406_), .C1(new_n411_), .C2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n392_), .A2(new_n405_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT20), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n382_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT97), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n360_), .A2(new_n361_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n382_), .A2(new_n386_), .A3(KEYINPUT97), .A4(new_n387_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n418_), .A2(new_n420_), .A3(new_n371_), .A4(new_n421_), .ZN(new_n422_));
  XOR2_X1   g221(.A(KEYINPUT22), .B(G169gat), .Z(new_n423_));
  OAI211_X1 g222(.A(new_n406_), .B(new_n359_), .C1(G176gat), .C2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n403_), .A2(new_n404_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n415_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n414_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G226gat), .A2(G233gat), .ZN(new_n429_));
  XOR2_X1   g228(.A(new_n429_), .B(KEYINPUT19), .Z(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(KEYINPUT96), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n388_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT82), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n416_), .A2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n391_), .A2(new_n433_), .A3(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT25), .B(G183gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT26), .B(G190gat), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n419_), .A2(KEYINPUT80), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n390_), .B1(new_n439_), .B2(new_n362_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n413_), .B1(new_n436_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n426_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n422_), .A2(new_n403_), .A3(new_n404_), .A4(new_n424_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n443_), .A2(KEYINPUT20), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(new_n444_), .A3(new_n430_), .ZN(new_n445_));
  XOR2_X1   g244(.A(G8gat), .B(G36gat), .Z(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT18), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G64gat), .B(G92gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n432_), .A2(new_n445_), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n449_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n443_), .A2(KEYINPUT20), .A3(new_n430_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n452_), .B1(new_n441_), .B2(new_n426_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n431_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n454_), .B1(new_n414_), .B2(new_n427_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n451_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n351_), .A2(new_n357_), .A3(new_n450_), .A4(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n331_), .B1(new_n341_), .B2(new_n344_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n335_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(new_n353_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n453_), .A2(new_n455_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n449_), .A2(KEYINPUT32), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n443_), .A2(KEYINPUT20), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT99), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT99), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n443_), .A2(new_n466_), .A3(KEYINPUT20), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n467_), .A3(new_n442_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n430_), .ZN(new_n469_));
  AND2_X1   g268(.A1(new_n414_), .A2(new_n427_), .ZN(new_n470_));
  AOI22_X1  g269(.A1(new_n468_), .A2(new_n469_), .B1(new_n470_), .B2(new_n454_), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n460_), .B(new_n463_), .C1(new_n471_), .C2(new_n462_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n457_), .A2(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n474_));
  OAI21_X1  g273(.A(new_n474_), .B1(new_n319_), .B2(KEYINPUT29), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G22gat), .B(G50gat), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT29), .ZN(new_n477_));
  INV_X1    g276(.A(new_n474_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n328_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n475_), .A2(new_n476_), .A3(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n476_), .B1(new_n475_), .B2(new_n479_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT94), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G228gat), .A2(G233gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n426_), .A2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n477_), .B1(new_n312_), .B2(new_n318_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n484_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n319_), .A2(KEYINPUT29), .ZN(new_n489_));
  INV_X1    g288(.A(new_n485_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n490_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n489_), .A2(KEYINPUT94), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n488_), .A2(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(G78gat), .B(G106gat), .Z(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n496_));
  OAI21_X1  g295(.A(new_n426_), .B1(new_n328_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(new_n490_), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n493_), .A2(new_n495_), .A3(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n495_), .B1(new_n493_), .B2(new_n498_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n483_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  NOR3_X1   g300(.A1(new_n486_), .A2(new_n487_), .A3(new_n484_), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT94), .B1(new_n489_), .B2(new_n491_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n498_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n494_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n493_), .A2(new_n495_), .A3(new_n498_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(new_n482_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n501_), .A2(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n352_), .B1(new_n349_), .B2(new_n331_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n353_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  AND3_X1   g310(.A1(new_n501_), .A2(new_n507_), .A3(new_n511_), .ZN(new_n512_));
  AOI22_X1  g311(.A1(new_n464_), .A2(KEYINPUT99), .B1(new_n441_), .B2(new_n426_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n430_), .B1(new_n513_), .B2(new_n467_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n428_), .A2(new_n431_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n451_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT27), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n517_), .B1(new_n461_), .B2(new_n449_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n456_), .A2(new_n450_), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n516_), .A2(new_n518_), .B1(new_n519_), .B2(new_n517_), .ZN(new_n520_));
  AOI22_X1  g319(.A1(new_n473_), .A2(new_n508_), .B1(new_n512_), .B2(new_n520_), .ZN(new_n521_));
  XOR2_X1   g320(.A(G71gat), .B(G99gat), .Z(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT85), .B(G43gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(KEYINPUT86), .B(G15gat), .Z(new_n525_));
  NAND2_X1  g324(.A1(G227gat), .A2(G233gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(new_n524_), .B(new_n527_), .Z(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n392_), .A2(KEYINPUT30), .A3(new_n413_), .ZN(new_n530_));
  AOI21_X1  g329(.A(KEYINPUT30), .B1(new_n392_), .B2(new_n413_), .ZN(new_n531_));
  NOR3_X1   g330(.A1(new_n530_), .A2(new_n531_), .A3(KEYINPUT87), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT87), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT30), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n441_), .A2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n392_), .A2(KEYINPUT30), .A3(new_n413_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n533_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n529_), .B1(new_n532_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT88), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT87), .B1(new_n530_), .B2(new_n531_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n528_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n538_), .A2(new_n539_), .A3(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n535_), .A2(new_n533_), .A3(new_n536_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n528_), .B1(new_n540_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n535_), .A2(new_n536_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n529_), .B1(new_n545_), .B2(KEYINPUT87), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT88), .B1(new_n544_), .B2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n542_), .A2(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n322_), .B(KEYINPUT31), .Z(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n542_), .A2(new_n547_), .A3(new_n549_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT100), .B1(new_n521_), .B2(new_n553_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n542_), .A2(new_n547_), .A3(new_n549_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n549_), .B1(new_n542_), .B2(new_n547_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT100), .ZN(new_n558_));
  AOI22_X1  g357(.A1(new_n457_), .A2(new_n472_), .B1(new_n507_), .B2(new_n501_), .ZN(new_n559_));
  OAI211_X1 g358(.A(KEYINPUT27), .B(new_n450_), .C1(new_n471_), .C2(new_n449_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n519_), .A2(new_n517_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n501_), .A2(new_n511_), .A3(new_n507_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n557_), .B(new_n558_), .C1(new_n559_), .C2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n508_), .A2(new_n561_), .A3(new_n560_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n566_), .B1(new_n552_), .B2(new_n551_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(new_n511_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n554_), .A2(new_n565_), .A3(new_n568_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n294_), .A2(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n278_), .B1(new_n222_), .B2(new_n229_), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n229_), .B(new_n272_), .C1(new_n219_), .C2(new_n221_), .ZN(new_n572_));
  XOR2_X1   g371(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n573_));
  NAND2_X1  g372(.A1(G232gat), .A2(G233gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT35), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n572_), .A2(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n571_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT71), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n572_), .A2(new_n580_), .A3(new_n577_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n575_), .A2(new_n576_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n583_), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n581_), .B(new_n582_), .C1(new_n571_), .C2(new_n578_), .ZN(new_n585_));
  AOI21_X1  g384(.A(KEYINPUT73), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G190gat), .B(G218gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G134gat), .B(G162gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT36), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n586_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n584_), .A2(KEYINPUT73), .A3(new_n585_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT37), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n589_), .A2(KEYINPUT36), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n584_), .A2(new_n585_), .A3(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n593_), .A2(new_n594_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n596_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n590_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n599_));
  OAI21_X1  g398(.A(KEYINPUT37), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT72), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  OAI211_X1 g401(.A(KEYINPUT72), .B(KEYINPUT37), .C1(new_n598_), .C2(new_n599_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n597_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(G231gat), .A2(G233gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n237_), .B(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(new_n269_), .ZN(new_n608_));
  XOR2_X1   g407(.A(G127gat), .B(G155gat), .Z(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT16), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G183gat), .B(G211gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT17), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n608_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT75), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT17), .ZN(new_n616_));
  OR3_X1    g415(.A1(new_n608_), .A2(new_n616_), .A3(new_n612_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n614_), .A2(KEYINPUT75), .ZN(new_n619_));
  OR3_X1    g418(.A1(new_n618_), .A2(KEYINPUT76), .A3(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(KEYINPUT76), .B1(new_n618_), .B2(new_n619_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n605_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n570_), .A2(new_n623_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n624_), .A2(G1gat), .A3(new_n511_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT101), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n626_), .A2(KEYINPUT38), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(KEYINPUT38), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT102), .ZN(new_n629_));
  INV_X1    g428(.A(new_n262_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(new_n292_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n629_), .B1(new_n631_), .B2(new_n622_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n593_), .A2(new_n596_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT103), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n557_), .B1(new_n559_), .B2(new_n564_), .ZN(new_n635_));
  AOI22_X1  g434(.A1(new_n635_), .A2(KEYINPUT100), .B1(new_n511_), .B2(new_n567_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n634_), .B1(new_n565_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n622_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n294_), .A2(KEYINPUT102), .A3(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n632_), .A2(new_n637_), .A3(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G1gat), .B1(new_n640_), .B2(new_n511_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n627_), .A2(new_n628_), .A3(new_n641_), .ZN(G1324gat));
  OR3_X1    g441(.A1(new_n624_), .A2(G8gat), .A3(new_n520_), .ZN(new_n643_));
  OR2_X1    g442(.A1(new_n640_), .A2(new_n520_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT39), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n644_), .A2(new_n645_), .A3(G8gat), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n645_), .B1(new_n644_), .B2(G8gat), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n643_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g449(.A(G15gat), .B1(new_n640_), .B2(new_n557_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT41), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n624_), .A2(G15gat), .A3(new_n557_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1326gat));
  OAI21_X1  g453(.A(G22gat), .B1(new_n640_), .B2(new_n508_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT42), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n508_), .A2(G22gat), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n656_), .B1(new_n624_), .B2(new_n657_), .ZN(G1327gat));
  NOR2_X1   g457(.A1(new_n638_), .A2(new_n633_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n570_), .A2(new_n659_), .ZN(new_n660_));
  OR3_X1    g459(.A1(new_n660_), .A2(G29gat), .A3(new_n511_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT105), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n604_), .B1(new_n636_), .B2(new_n565_), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n662_), .B(KEYINPUT43), .C1(new_n663_), .C2(KEYINPUT104), .ZN(new_n664_));
  AND4_X1   g463(.A1(new_n622_), .A2(new_n258_), .A3(new_n261_), .A4(new_n292_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT43), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n666_), .B1(new_n663_), .B2(new_n662_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n569_), .A2(new_n605_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT104), .ZN(new_n669_));
  AOI21_X1  g468(.A(KEYINPUT105), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  OAI211_X1 g469(.A(new_n664_), .B(new_n665_), .C1(new_n667_), .C2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n672_));
  OR3_X1    g471(.A1(new_n671_), .A2(KEYINPUT109), .A3(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(KEYINPUT109), .B1(new_n671_), .B2(new_n672_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n675_), .A2(new_n511_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n671_), .A2(KEYINPUT106), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n662_), .B1(new_n663_), .B2(KEYINPUT104), .ZN(new_n678_));
  AOI21_X1  g477(.A(KEYINPUT43), .B1(new_n668_), .B2(KEYINPUT105), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT106), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n680_), .A2(new_n681_), .A3(new_n664_), .A4(new_n665_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n677_), .A2(new_n682_), .ZN(new_n683_));
  XOR2_X1   g482(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT108), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n683_), .A2(KEYINPUT108), .A3(new_n684_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n676_), .A2(new_n689_), .A3(KEYINPUT110), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(G29gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(KEYINPUT110), .B1(new_n676_), .B2(new_n689_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n661_), .B1(new_n691_), .B2(new_n692_), .ZN(G1328gat));
  INV_X1    g492(.A(G36gat), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n675_), .A2(new_n520_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n695_), .B2(new_n689_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT46), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n660_), .A2(G36gat), .A3(new_n520_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT45), .ZN(new_n699_));
  OR3_X1    g498(.A1(new_n696_), .A2(new_n697_), .A3(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n697_), .B1(new_n696_), .B2(new_n699_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1329gat));
  INV_X1    g501(.A(G43gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n703_), .B1(new_n660_), .B2(new_n557_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT111), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n553_), .A2(G43gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n705_), .B1(new_n689_), .B2(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(KEYINPUT108), .B1(new_n683_), .B2(new_n684_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n684_), .ZN(new_n710_));
  AOI211_X1 g509(.A(new_n686_), .B(new_n710_), .C1(new_n677_), .C2(new_n682_), .ZN(new_n711_));
  OAI211_X1 g510(.A(new_n707_), .B(new_n705_), .C1(new_n709_), .C2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n704_), .B1(new_n708_), .B2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT47), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT47), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n716_), .B(new_n704_), .C1(new_n708_), .C2(new_n713_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(G1330gat));
  INV_X1    g517(.A(new_n660_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n508_), .ZN(new_n720_));
  AOI21_X1  g519(.A(G50gat), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(G50gat), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n675_), .A2(new_n722_), .A3(new_n508_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n721_), .B1(new_n723_), .B2(new_n689_), .ZN(G1331gat));
  NAND4_X1  g523(.A1(new_n637_), .A2(new_n638_), .A3(new_n293_), .A4(new_n262_), .ZN(new_n725_));
  OAI21_X1  g524(.A(G57gat), .B1(new_n725_), .B2(new_n511_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n262_), .A2(new_n569_), .A3(new_n293_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(new_n623_), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n511_), .A2(G57gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n726_), .B1(new_n728_), .B2(new_n729_), .ZN(G1332gat));
  OAI21_X1  g529(.A(G64gat), .B1(new_n725_), .B2(new_n520_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT48), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n520_), .A2(G64gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n728_), .B2(new_n733_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT112), .Z(G1333gat));
  OAI21_X1  g534(.A(G71gat), .B1(new_n725_), .B2(new_n557_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT49), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n557_), .A2(G71gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n737_), .B1(new_n728_), .B2(new_n738_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT113), .Z(G1334gat));
  OAI21_X1  g539(.A(G78gat), .B1(new_n725_), .B2(new_n508_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT50), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n508_), .A2(G78gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n742_), .B1(new_n728_), .B2(new_n743_), .ZN(G1335gat));
  NAND2_X1  g543(.A1(new_n727_), .A2(new_n659_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(G85gat), .B1(new_n746_), .B2(new_n460_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n630_), .A2(new_n638_), .A3(new_n292_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n748_), .A2(new_n680_), .A3(new_n664_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n460_), .A2(new_n226_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n747_), .B1(new_n749_), .B2(new_n750_), .ZN(G1336gat));
  NOR3_X1   g550(.A1(new_n745_), .A2(G92gat), .A3(new_n520_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n749_), .A2(new_n562_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n753_), .B2(G92gat), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT114), .Z(G1337gat));
  NAND3_X1  g554(.A1(new_n746_), .A2(new_n223_), .A3(new_n553_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n749_), .A2(new_n553_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n757_), .A2(KEYINPUT115), .A3(G99gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT115), .B1(new_n757_), .B2(G99gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n756_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g560(.A(KEYINPUT116), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n749_), .A2(new_n720_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(G106gat), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n746_), .A2(new_n224_), .A3(new_n720_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  AOI211_X1 g567(.A(KEYINPUT116), .B(new_n224_), .C1(new_n749_), .C2(new_n720_), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n764_), .A2(new_n769_), .A3(new_n765_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n768_), .A2(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n771_), .B(new_n772_), .ZN(G1339gat));
  NAND2_X1  g572(.A1(new_n567_), .A2(new_n460_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT122), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n242_), .A2(new_n776_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n240_), .A2(new_n241_), .A3(G230gat), .A4(G233gat), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n250_), .B1(new_n242_), .B2(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT56), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT119), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n779_), .A2(KEYINPUT56), .A3(new_n780_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n783_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n781_), .A2(KEYINPUT119), .A3(new_n782_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n786_), .A2(new_n292_), .A3(new_n251_), .A4(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n289_), .ZN(new_n789_));
  OR3_X1    g588(.A1(new_n279_), .A2(new_n280_), .A3(new_n274_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n288_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n789_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(new_n259_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n788_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n633_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT120), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n796_), .A2(KEYINPUT57), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT121), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n783_), .A2(new_n798_), .A3(new_n785_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n779_), .A2(KEYINPUT121), .A3(KEYINPUT56), .A4(new_n780_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n792_), .A2(new_n251_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n799_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT58), .ZN(new_n803_));
  OR2_X1    g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n604_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n805_));
  AOI22_X1  g604(.A1(new_n795_), .A2(new_n797_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n794_), .B(new_n633_), .C1(new_n796_), .C2(KEYINPUT57), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n638_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n293_), .A2(new_n638_), .A3(KEYINPUT118), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n260_), .A2(new_n255_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT118), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n292_), .B2(new_n622_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n809_), .A2(new_n810_), .A3(new_n812_), .ZN(new_n813_));
  OR3_X1    g612(.A1(new_n813_), .A2(KEYINPUT54), .A3(new_n605_), .ZN(new_n814_));
  OAI21_X1  g613(.A(KEYINPUT54), .B1(new_n813_), .B2(new_n605_), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n775_), .B1(new_n808_), .B2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n795_), .A2(new_n797_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n804_), .A2(new_n805_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n807_), .A3(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n622_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n814_), .A2(new_n815_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n821_), .A2(KEYINPUT122), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n774_), .B1(new_n817_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(G113gat), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n824_), .A2(new_n825_), .A3(new_n292_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n808_), .A2(new_n816_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT59), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n567_), .A2(new_n828_), .A3(new_n460_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n827_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n831_), .B(new_n292_), .C1(new_n824_), .C2(new_n828_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n826_), .B1(new_n833_), .B2(new_n825_), .ZN(G1340gat));
  INV_X1    g633(.A(G120gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n835_), .B1(new_n630_), .B2(KEYINPUT60), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n824_), .B(new_n836_), .C1(KEYINPUT60), .C2(new_n835_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n831_), .B(new_n262_), .C1(new_n824_), .C2(new_n828_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n837_), .B1(new_n839_), .B2(new_n835_), .ZN(G1341gat));
  AOI21_X1  g639(.A(G127gat), .B1(new_n824_), .B2(new_n638_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n824_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n830_), .B1(new_n842_), .B2(KEYINPUT59), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n622_), .A2(KEYINPUT123), .ZN(new_n844_));
  MUX2_X1   g643(.A(KEYINPUT123), .B(new_n844_), .S(G127gat), .Z(new_n845_));
  AOI21_X1  g644(.A(new_n841_), .B1(new_n843_), .B2(new_n845_), .ZN(G1342gat));
  AOI21_X1  g645(.A(G134gat), .B1(new_n824_), .B2(new_n634_), .ZN(new_n847_));
  XOR2_X1   g646(.A(KEYINPUT124), .B(G134gat), .Z(new_n848_));
  NOR2_X1   g647(.A1(new_n604_), .A2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n847_), .B1(new_n843_), .B2(new_n849_), .ZN(G1343gat));
  AOI21_X1  g649(.A(new_n553_), .B1(new_n817_), .B2(new_n823_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n562_), .A2(new_n508_), .A3(new_n511_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n292_), .A3(new_n852_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g653(.A1(new_n851_), .A2(new_n262_), .A3(new_n852_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g655(.A1(new_n851_), .A2(new_n638_), .A3(new_n852_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(KEYINPUT61), .B(G155gat), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(G1346gat));
  NAND2_X1  g658(.A1(new_n851_), .A2(new_n852_), .ZN(new_n860_));
  OAI21_X1  g659(.A(G162gat), .B1(new_n860_), .B2(new_n604_), .ZN(new_n861_));
  INV_X1    g660(.A(G162gat), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n634_), .A2(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n861_), .B1(new_n860_), .B2(new_n863_), .ZN(G1347gat));
  INV_X1    g663(.A(KEYINPUT62), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n557_), .A2(new_n460_), .A3(new_n520_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n508_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n827_), .A2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n292_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n865_), .B1(new_n869_), .B2(G169gat), .ZN(new_n870_));
  AOI211_X1 g669(.A(KEYINPUT62), .B(new_n372_), .C1(new_n868_), .C2(new_n292_), .ZN(new_n871_));
  OAI21_X1  g670(.A(KEYINPUT125), .B1(new_n827_), .B2(new_n867_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT125), .ZN(new_n873_));
  INV_X1    g672(.A(new_n867_), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n873_), .B(new_n874_), .C1(new_n808_), .C2(new_n816_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n872_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n293_), .A2(new_n423_), .ZN(new_n878_));
  OAI22_X1  g677(.A1(new_n870_), .A2(new_n871_), .B1(new_n877_), .B2(new_n878_), .ZN(G1348gat));
  AOI21_X1  g678(.A(G176gat), .B1(new_n876_), .B2(new_n262_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n720_), .B1(new_n817_), .B2(new_n823_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT126), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n866_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  AOI211_X1 g682(.A(KEYINPUT126), .B(new_n720_), .C1(new_n817_), .C2(new_n823_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n630_), .A2(new_n373_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n880_), .B1(new_n885_), .B2(new_n886_), .ZN(G1349gat));
  AOI211_X1 g686(.A(new_n622_), .B(new_n437_), .C1(new_n872_), .C2(new_n875_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n817_), .A2(new_n823_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n508_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT126), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n881_), .A2(new_n882_), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n891_), .A2(new_n638_), .A3(new_n892_), .A4(new_n866_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n888_), .B1(new_n893_), .B2(new_n363_), .ZN(G1350gat));
  OAI21_X1  g693(.A(G190gat), .B1(new_n877_), .B2(new_n604_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n876_), .A2(new_n438_), .A3(new_n634_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(G1351gat));
  NOR2_X1   g696(.A1(new_n520_), .A2(new_n563_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n851_), .A2(new_n292_), .A3(new_n898_), .ZN(new_n899_));
  XOR2_X1   g698(.A(KEYINPUT127), .B(G197gat), .Z(new_n900_));
  XNOR2_X1  g699(.A(new_n899_), .B(new_n900_), .ZN(G1352gat));
  NAND3_X1  g700(.A1(new_n851_), .A2(new_n262_), .A3(new_n898_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g702(.A1(new_n851_), .A2(new_n638_), .A3(new_n898_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(KEYINPUT63), .B(G211gat), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n904_), .B2(new_n907_), .ZN(G1354gat));
  NAND2_X1  g707(.A1(new_n851_), .A2(new_n898_), .ZN(new_n909_));
  OAI21_X1  g708(.A(G218gat), .B1(new_n909_), .B2(new_n604_), .ZN(new_n910_));
  INV_X1    g709(.A(G218gat), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n634_), .A2(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n910_), .B1(new_n909_), .B2(new_n912_), .ZN(G1355gat));
endmodule


