//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n897_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_;
  XNOR2_X1  g000(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT23), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n205_), .A2(G183gat), .A3(G190gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT83), .ZN(new_n207_));
  INV_X1    g006(.A(G183gat), .ZN(new_n208_));
  INV_X1    g007(.A(G190gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT23), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n207_), .B(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n208_), .A2(new_n209_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT22), .B(G169gat), .ZN(new_n216_));
  INV_X1    g015(.A(G176gat), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n215_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n213_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT26), .B(G190gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT25), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n220_), .B1(new_n221_), .B2(G183gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(KEYINPUT80), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT80), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT25), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n208_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n226_), .A2(KEYINPUT81), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(KEYINPUT81), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n222_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  AND3_X1   g028(.A1(new_n210_), .A2(KEYINPUT82), .A3(new_n206_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n206_), .B1(new_n210_), .B2(KEYINPUT82), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n233_), .A2(KEYINPUT24), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(KEYINPUT24), .A3(new_n214_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n232_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n219_), .B1(new_n229_), .B2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G211gat), .B(G218gat), .ZN(new_n238_));
  INV_X1    g037(.A(G197gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(G204gat), .ZN(new_n240_));
  INV_X1    g039(.A(G204gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(G197gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n243_), .A2(KEYINPUT89), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT89), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT21), .B1(new_n240_), .B2(new_n245_), .ZN(new_n246_));
  OAI221_X1 g045(.A(new_n238_), .B1(KEYINPUT21), .B2(new_n243_), .C1(new_n244_), .C2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n243_), .A2(KEYINPUT21), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n248_), .A2(new_n238_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT20), .B1(new_n237_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n250_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n216_), .B(KEYINPUT96), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n215_), .B1(new_n253_), .B2(new_n217_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT97), .ZN(new_n255_));
  AND3_X1   g054(.A1(new_n232_), .A2(new_n255_), .A3(new_n212_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n255_), .B1(new_n232_), .B2(new_n212_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n254_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT25), .B(G183gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n220_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(new_n235_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT95), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n262_), .A2(new_n211_), .A3(new_n234_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n252_), .B1(new_n258_), .B2(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n204_), .B1(new_n251_), .B2(new_n264_), .ZN(new_n265_));
  XOR2_X1   g064(.A(G8gat), .B(G36gat), .Z(new_n266_));
  XNOR2_X1  g065(.A(G64gat), .B(G92gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT20), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n272_), .B1(new_n237_), .B2(new_n250_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n258_), .A2(new_n263_), .A3(new_n252_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n204_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n265_), .A2(new_n271_), .A3(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT27), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n251_), .A2(new_n264_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n275_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n275_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n271_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n283_));
  OR3_X1    g082(.A1(new_n278_), .A2(new_n283_), .A3(KEYINPUT101), .ZN(new_n284_));
  XOR2_X1   g083(.A(G127gat), .B(G134gat), .Z(new_n285_));
  XOR2_X1   g084(.A(G113gat), .B(G120gat), .Z(new_n286_));
  XOR2_X1   g085(.A(new_n285_), .B(new_n286_), .Z(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(G155gat), .A2(G162gat), .ZN(new_n289_));
  INV_X1    g088(.A(G155gat), .ZN(new_n290_));
  INV_X1    g089(.A(G162gat), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT1), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n289_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n294_), .B1(new_n293_), .B2(new_n292_), .ZN(new_n295_));
  INV_X1    g094(.A(G141gat), .ZN(new_n296_));
  INV_X1    g095(.A(G148gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G141gat), .A2(G148gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT84), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n295_), .A2(new_n298_), .A3(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(KEYINPUT85), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT3), .ZN(new_n303_));
  NOR2_X1   g102(.A1(G141gat), .A2(G148gat), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT85), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n302_), .A2(new_n303_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT86), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT2), .ZN(new_n310_));
  OAI22_X1  g109(.A1(new_n304_), .A2(new_n303_), .B1(new_n299_), .B2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n311_), .B1(new_n300_), .B2(new_n310_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n292_), .A2(new_n289_), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n288_), .B(new_n301_), .C1(new_n313_), .C2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT100), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n314_), .B1(new_n309_), .B2(new_n312_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n301_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n316_), .B(new_n287_), .C1(new_n317_), .C2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n315_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT4), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G225gat), .A2(G233gat), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT4), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n319_), .A2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n321_), .A2(new_n323_), .A3(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G1gat), .B(G29gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(G85gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT0), .B(G57gat), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n328_), .B(new_n329_), .Z(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n317_), .A2(new_n318_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(new_n288_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(new_n322_), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n326_), .A2(new_n331_), .A3(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n331_), .B1(new_n326_), .B2(new_n334_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT27), .ZN(new_n338_));
  INV_X1    g137(.A(new_n277_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n271_), .B1(new_n265_), .B2(new_n276_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n338_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT101), .B1(new_n278_), .B2(new_n283_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n284_), .A2(new_n337_), .A3(new_n341_), .A4(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G71gat), .B(G99gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(G43gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n237_), .B(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(new_n287_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G227gat), .A2(G233gat), .ZN(new_n348_));
  INV_X1    g147(.A(G15gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT30), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT31), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n347_), .B(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT29), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n332_), .A2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT88), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  XOR2_X1   g157(.A(G22gat), .B(G50gat), .Z(new_n359_));
  NOR4_X1   g158(.A1(new_n317_), .A2(KEYINPUT29), .A3(new_n318_), .A4(new_n357_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n358_), .A2(new_n359_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n359_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n357_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n364_), .B1(new_n332_), .B2(new_n354_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n363_), .B1(new_n365_), .B2(new_n360_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n362_), .A2(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(KEYINPUT91), .B(KEYINPUT29), .Z(new_n368_));
  OAI21_X1  g167(.A(new_n368_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(new_n250_), .ZN(new_n370_));
  AND2_X1   g169(.A1(G228gat), .A2(G233gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT93), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G78gat), .B(G106gat), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(KEYINPUT29), .B1(new_n317_), .B2(new_n318_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n252_), .A2(new_n371_), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n376_), .A2(KEYINPUT90), .A3(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(KEYINPUT90), .B1(new_n376_), .B2(new_n377_), .ZN(new_n379_));
  OAI221_X1 g178(.A(new_n372_), .B1(new_n373_), .B2(new_n375_), .C1(new_n378_), .C2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n372_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n374_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n367_), .B(new_n380_), .C1(new_n382_), .C2(new_n373_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n372_), .B(new_n375_), .C1(new_n378_), .C2(new_n379_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n367_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT92), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n383_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  AOI211_X1 g186(.A(KEYINPUT92), .B(new_n367_), .C1(new_n382_), .C2(new_n384_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n353_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n367_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n376_), .A2(new_n377_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT90), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n376_), .A2(KEYINPUT90), .A3(new_n377_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n375_), .B1(new_n395_), .B2(new_n372_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n384_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n390_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT92), .ZN(new_n399_));
  INV_X1    g198(.A(new_n352_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n347_), .B(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n385_), .A2(new_n386_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n399_), .A2(new_n401_), .A3(new_n402_), .A4(new_n383_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n343_), .B1(new_n389_), .B2(new_n403_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n399_), .A2(new_n353_), .A3(new_n402_), .A4(new_n383_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n271_), .A2(KEYINPUT32), .ZN(new_n406_));
  INV_X1    g205(.A(new_n280_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n406_), .B1(new_n407_), .B2(new_n281_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n265_), .A2(new_n276_), .ZN(new_n409_));
  OAI221_X1 g208(.A(new_n408_), .B1(new_n409_), .B2(new_n406_), .C1(new_n335_), .C2(new_n336_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT33), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n336_), .B(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n323_), .B1(new_n321_), .B2(new_n325_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n331_), .B1(new_n333_), .B2(new_n322_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT99), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n416_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n340_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n418_), .A2(KEYINPUT99), .A3(new_n277_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n415_), .B1(new_n417_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n412_), .A2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n405_), .B1(new_n410_), .B2(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n404_), .A2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G113gat), .B(G141gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT78), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G169gat), .B(G197gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT76), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G1gat), .B(G8gat), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n429_), .A2(KEYINPUT72), .ZN(new_n430_));
  INV_X1    g229(.A(G22gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n349_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G15gat), .A2(G22gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G1gat), .A2(G8gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT14), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n429_), .A2(KEYINPUT72), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n430_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n437_), .B1(new_n430_), .B2(new_n438_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G29gat), .B(G36gat), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  XOR2_X1   g242(.A(G43gat), .B(G50gat), .Z(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G43gat), .B(G50gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n442_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  NOR3_X1   g247(.A1(new_n440_), .A2(new_n441_), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n448_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n430_), .A2(new_n438_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n437_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n450_), .B1(new_n453_), .B2(new_n439_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n428_), .B1(new_n449_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G229gat), .A2(G233gat), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n448_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n453_), .A2(new_n450_), .A3(new_n439_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(KEYINPUT76), .A3(new_n459_), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n455_), .A2(new_n457_), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT15), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n448_), .A2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n445_), .A2(KEYINPUT15), .A3(new_n447_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n463_), .A2(new_n453_), .A3(new_n439_), .A4(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n465_), .A2(new_n458_), .A3(new_n456_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT77), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT77), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n465_), .A2(new_n458_), .A3(new_n468_), .A4(new_n456_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n427_), .B1(new_n461_), .B2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n455_), .A2(new_n457_), .A3(new_n460_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n427_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n472_), .A2(new_n467_), .A3(new_n469_), .A4(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n471_), .A2(KEYINPUT79), .A3(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT79), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n476_), .B(new_n427_), .C1(new_n461_), .C2(new_n470_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n423_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G99gat), .A2(G106gat), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT6), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  OR2_X1    g283(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n485_));
  INV_X1    g284(.A(G106gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n485_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G85gat), .A2(G92gat), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n489_), .A2(KEYINPUT9), .ZN(new_n490_));
  OR2_X1    g289(.A1(G85gat), .A2(G92gat), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n491_), .A2(KEYINPUT9), .A3(new_n489_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n484_), .A2(new_n488_), .A3(new_n490_), .A4(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT7), .ZN(new_n494_));
  INV_X1    g293(.A(G99gat), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n494_), .A2(new_n495_), .A3(new_n486_), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n496_), .A2(new_n482_), .A3(new_n483_), .A4(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT8), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n491_), .A2(new_n489_), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n498_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n499_), .B1(new_n498_), .B2(new_n500_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n493_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT64), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT64), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n505_), .B(new_n493_), .C1(new_n501_), .C2(new_n502_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n504_), .A2(new_n448_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G232gat), .A2(G233gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT34), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n509_), .A2(KEYINPUT35), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT68), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n507_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT35), .ZN(new_n513_));
  INV_X1    g312(.A(new_n509_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n463_), .A2(new_n464_), .ZN(new_n515_));
  AOI21_X1  g314(.A(KEYINPUT67), .B1(new_n515_), .B2(new_n503_), .ZN(new_n516_));
  AND3_X1   g315(.A1(new_n515_), .A2(KEYINPUT67), .A3(new_n503_), .ZN(new_n517_));
  OAI221_X1 g316(.A(new_n512_), .B1(new_n513_), .B2(new_n514_), .C1(new_n516_), .C2(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n517_), .A2(new_n516_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n507_), .A2(new_n511_), .ZN(new_n520_));
  OAI211_X1 g319(.A(KEYINPUT35), .B(new_n509_), .C1(new_n519_), .C2(new_n520_), .ZN(new_n521_));
  XOR2_X1   g320(.A(G190gat), .B(G218gat), .Z(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT69), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G134gat), .B(G162gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n525_), .A2(KEYINPUT36), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n518_), .A2(new_n521_), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n525_), .B(KEYINPUT36), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n529_), .B1(new_n518_), .B2(new_n521_), .ZN(new_n530_));
  OAI21_X1  g329(.A(KEYINPUT37), .B1(new_n528_), .B2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(KEYINPUT70), .B(KEYINPUT37), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n518_), .A2(new_n521_), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n527_), .B(new_n532_), .C1(new_n533_), .C2(new_n529_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n531_), .A2(new_n534_), .A3(KEYINPUT71), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n528_), .A2(new_n530_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT71), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n536_), .A2(new_n537_), .A3(new_n532_), .ZN(new_n538_));
  XOR2_X1   g337(.A(KEYINPUT73), .B(KEYINPUT16), .Z(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT74), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G127gat), .B(G155gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G183gat), .B(G211gat), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n542_), .B(new_n543_), .Z(new_n544_));
  INV_X1    g343(.A(KEYINPUT17), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(G64gat), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(G57gat), .ZN(new_n548_));
  INV_X1    g347(.A(G57gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(G64gat), .ZN(new_n550_));
  AOI21_X1  g349(.A(KEYINPUT65), .B1(new_n548_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n548_), .A2(new_n550_), .A3(KEYINPUT65), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT11), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n548_), .A2(new_n550_), .A3(KEYINPUT65), .ZN(new_n556_));
  OAI21_X1  g355(.A(KEYINPUT11), .B1(new_n556_), .B2(new_n551_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G71gat), .B(G78gat), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n555_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n560_));
  OAI211_X1 g359(.A(KEYINPUT11), .B(new_n558_), .C1(new_n556_), .C2(new_n551_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G231gat), .A2(G233gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n440_), .A2(new_n441_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n546_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n566_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n568_), .B1(new_n545_), .B2(new_n544_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(G230gat), .ZN(new_n571_));
  INV_X1    g370(.A(G233gat), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n504_), .A2(new_n506_), .A3(new_n562_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n562_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n573_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n504_), .A2(new_n506_), .A3(new_n562_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n560_), .A2(new_n561_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n578_), .A2(KEYINPUT12), .A3(new_n503_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n577_), .B(new_n579_), .C1(new_n575_), .C2(KEYINPUT12), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n576_), .B1(new_n580_), .B2(new_n573_), .ZN(new_n581_));
  XOR2_X1   g380(.A(G120gat), .B(G148gat), .Z(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT66), .B(KEYINPUT5), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G176gat), .B(G204gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n581_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n586_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n576_), .B(new_n588_), .C1(new_n580_), .C2(new_n573_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT13), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n535_), .A2(new_n538_), .A3(new_n570_), .A4(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n593_), .A2(KEYINPUT75), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(KEYINPUT75), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n479_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  NOR3_X1   g395(.A1(new_n596_), .A2(G1gat), .A3(new_n337_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n600_), .B(KEYINPUT103), .Z(new_n601_));
  NOR2_X1   g400(.A1(new_n423_), .A2(new_n536_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n337_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n478_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n591_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n570_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n602_), .A2(new_n603_), .A3(new_n607_), .ZN(new_n608_));
  AOI22_X1  g407(.A1(new_n598_), .A2(new_n599_), .B1(G1gat), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n601_), .A2(new_n609_), .ZN(G1324gat));
  NAND2_X1  g409(.A1(new_n602_), .A2(new_n607_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n342_), .A2(new_n341_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(new_n284_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(G8gat), .B1(new_n611_), .B2(new_n614_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n615_), .A2(KEYINPUT104), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(KEYINPUT104), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n616_), .A2(KEYINPUT39), .A3(new_n617_), .ZN(new_n618_));
  OR3_X1    g417(.A1(new_n596_), .A2(G8gat), .A3(new_n614_), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n618_), .B(new_n619_), .C1(KEYINPUT39), .C2(new_n617_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT40), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(G1325gat));
  OAI21_X1  g421(.A(G15gat), .B1(new_n611_), .B2(new_n353_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n624_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n401_), .A2(new_n349_), .ZN(new_n627_));
  OAI211_X1 g426(.A(new_n625_), .B(new_n626_), .C1(new_n596_), .C2(new_n627_), .ZN(G1326gat));
  NOR2_X1   g427(.A1(new_n387_), .A2(new_n388_), .ZN(new_n629_));
  OAI21_X1  g428(.A(G22gat), .B1(new_n611_), .B2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT42), .ZN(new_n631_));
  INV_X1    g430(.A(new_n629_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(new_n431_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n631_), .B1(new_n596_), .B2(new_n633_), .ZN(G1327gat));
  INV_X1    g433(.A(new_n591_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n536_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n635_), .A2(new_n636_), .A3(new_n570_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n479_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(G29gat), .B1(new_n639_), .B2(new_n603_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n605_), .A2(new_n570_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT43), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n389_), .A2(new_n403_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n343_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n421_), .A2(new_n410_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n405_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n645_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n535_), .A2(new_n538_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n642_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n642_), .B(new_n650_), .C1(new_n404_), .C2(new_n422_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  OAI211_X1 g452(.A(KEYINPUT44), .B(new_n641_), .C1(new_n651_), .C2(new_n653_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n654_), .A2(G29gat), .A3(new_n603_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n650_), .ZN(new_n656_));
  OAI21_X1  g455(.A(KEYINPUT43), .B1(new_n423_), .B2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(new_n652_), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT44), .B1(new_n658_), .B2(new_n641_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n640_), .B1(new_n655_), .B2(new_n660_), .ZN(G1328gat));
  INV_X1    g460(.A(KEYINPUT107), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT46), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT45), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n614_), .A2(G36gat), .ZN(new_n665_));
  OR3_X1    g464(.A1(new_n638_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n664_), .B1(new_n638_), .B2(new_n665_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n654_), .A2(new_n613_), .ZN(new_n669_));
  OAI21_X1  g468(.A(G36gat), .B1(new_n669_), .B2(new_n659_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n668_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  OAI211_X1 g471(.A(KEYINPUT106), .B(G36gat), .C1(new_n669_), .C2(new_n659_), .ZN(new_n673_));
  AOI211_X1 g472(.A(new_n662_), .B(new_n663_), .C1(new_n672_), .C2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n670_), .A2(new_n671_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n668_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n675_), .A2(new_n673_), .A3(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT46), .B1(new_n677_), .B2(KEYINPUT107), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n674_), .A2(new_n678_), .ZN(G1329gat));
  NAND3_X1  g478(.A1(new_n654_), .A2(G43gat), .A3(new_n401_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n638_), .A2(new_n353_), .ZN(new_n681_));
  OAI22_X1  g480(.A1(new_n680_), .A2(new_n659_), .B1(G43gat), .B2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g482(.A(G50gat), .B1(new_n639_), .B2(new_n632_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n654_), .A2(G50gat), .A3(new_n632_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n685_), .B2(new_n660_), .ZN(G1331gat));
  NOR2_X1   g485(.A1(new_n591_), .A2(new_n604_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n649_), .A2(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n688_), .A2(new_n656_), .A3(new_n570_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n337_), .B1(new_n690_), .B2(KEYINPUT108), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n691_), .B1(KEYINPUT108), .B2(new_n690_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n602_), .A2(new_n570_), .A3(new_n687_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT109), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n337_), .A2(new_n549_), .ZN(new_n696_));
  AOI22_X1  g495(.A1(new_n692_), .A2(new_n549_), .B1(new_n695_), .B2(new_n696_), .ZN(G1332gat));
  AOI21_X1  g496(.A(new_n547_), .B1(new_n695_), .B2(new_n613_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT48), .Z(new_n699_));
  NAND3_X1  g498(.A1(new_n690_), .A2(new_n547_), .A3(new_n613_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1333gat));
  INV_X1    g500(.A(G71gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n702_), .B1(new_n695_), .B2(new_n401_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT49), .Z(new_n704_));
  NAND3_X1  g503(.A1(new_n690_), .A2(new_n702_), .A3(new_n401_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1334gat));
  INV_X1    g505(.A(G78gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n707_), .B1(new_n695_), .B2(new_n632_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT50), .Z(new_n709_));
  NAND3_X1  g508(.A1(new_n690_), .A2(new_n707_), .A3(new_n632_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1335gat));
  NAND3_X1  g510(.A1(new_n688_), .A2(new_n536_), .A3(new_n606_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(G85gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n713_), .A2(new_n714_), .A3(new_n603_), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n658_), .A2(new_n606_), .A3(new_n687_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n716_), .A2(new_n603_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n715_), .B1(new_n717_), .B2(new_n714_), .ZN(G1336gat));
  AOI21_X1  g517(.A(G92gat), .B1(new_n713_), .B2(new_n613_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n613_), .A2(G92gat), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT110), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n719_), .B1(new_n716_), .B2(new_n721_), .ZN(G1337gat));
  AND4_X1   g521(.A1(new_n401_), .A2(new_n713_), .A3(new_n485_), .A4(new_n487_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n495_), .B1(new_n716_), .B2(new_n401_), .ZN(new_n724_));
  OAI22_X1  g523(.A1(new_n723_), .A2(new_n724_), .B1(KEYINPUT111), .B2(KEYINPUT51), .ZN(new_n725_));
  NAND2_X1  g524(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT112), .Z(new_n727_));
  XNOR2_X1  g526(.A(new_n725_), .B(new_n727_), .ZN(G1338gat));
  NAND3_X1  g527(.A1(new_n713_), .A2(new_n486_), .A3(new_n632_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT52), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n716_), .A2(new_n632_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n731_), .B2(G106gat), .ZN(new_n732_));
  AOI211_X1 g531(.A(KEYINPUT52), .B(new_n486_), .C1(new_n716_), .C2(new_n632_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n729_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT53), .ZN(G1339gat));
  OAI21_X1  g534(.A(KEYINPUT54), .B1(new_n592_), .B2(new_n604_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT113), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  OAI211_X1 g537(.A(KEYINPUT113), .B(KEYINPUT54), .C1(new_n592_), .C2(new_n604_), .ZN(new_n739_));
  OR3_X1    g538(.A1(new_n592_), .A2(KEYINPUT54), .A3(new_n604_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n738_), .A2(new_n739_), .A3(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n455_), .A2(new_n456_), .A3(new_n460_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n465_), .A2(new_n458_), .A3(new_n457_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n742_), .A2(new_n427_), .A3(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n474_), .A2(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT116), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n746_), .B(new_n747_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n475_), .A2(new_n477_), .A3(new_n589_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT55), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n750_), .B1(new_n580_), .B2(new_n573_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n573_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n752_), .A2(KEYINPUT114), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n753_), .B1(new_n580_), .B2(new_n750_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n579_), .A2(new_n577_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n498_), .A2(new_n500_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT8), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n498_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n505_), .B1(new_n759_), .B2(new_n493_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n506_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n578_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT12), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n753_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n755_), .A2(new_n764_), .A3(KEYINPUT55), .A4(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n751_), .A2(new_n754_), .A3(new_n766_), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n767_), .A2(KEYINPUT56), .A3(new_n586_), .ZN(new_n768_));
  XOR2_X1   g567(.A(KEYINPUT115), .B(KEYINPUT56), .Z(new_n769_));
  AOI21_X1  g568(.A(new_n769_), .B1(new_n767_), .B2(new_n586_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n749_), .B1(new_n768_), .B2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n748_), .A2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT57), .B1(new_n772_), .B2(new_n636_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT57), .ZN(new_n774_));
  AOI211_X1 g573(.A(new_n774_), .B(new_n536_), .C1(new_n748_), .C2(new_n771_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n589_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n777_), .A2(new_n745_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n767_), .A2(new_n586_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT56), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n767_), .A2(KEYINPUT56), .A3(new_n586_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n779_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(KEYINPUT58), .B1(new_n784_), .B2(KEYINPUT117), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT56), .B1(new_n767_), .B2(new_n586_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n778_), .B1(new_n768_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT117), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT58), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n787_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n785_), .A2(new_n650_), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT118), .B1(new_n776_), .B2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n475_), .A2(new_n477_), .A3(new_n589_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n769_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n780_), .A2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n793_), .B1(new_n795_), .B2(new_n783_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n474_), .A2(new_n744_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n755_), .A2(new_n764_), .A3(new_n752_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n588_), .B1(new_n798_), .B2(new_n576_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n797_), .B1(new_n777_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n747_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n746_), .A2(KEYINPUT116), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n636_), .B1(new_n796_), .B2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n774_), .ZN(new_n805_));
  OAI211_X1 g604(.A(KEYINPUT57), .B(new_n636_), .C1(new_n796_), .C2(new_n803_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n791_), .A2(new_n805_), .A3(KEYINPUT118), .A4(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n606_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n741_), .B1(new_n792_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT119), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  OAI211_X1 g610(.A(KEYINPUT119), .B(new_n741_), .C1(new_n792_), .C2(new_n808_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n613_), .A2(new_n337_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n814_), .A2(new_n403_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n811_), .A2(new_n812_), .A3(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT59), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n791_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n606_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n741_), .A2(new_n819_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n815_), .A3(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(G113gat), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n478_), .A2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n817_), .A2(new_n822_), .A3(new_n824_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n811_), .A2(new_n604_), .A3(new_n812_), .A4(new_n815_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT120), .ZN(new_n827_));
  AND3_X1   g626(.A1(new_n826_), .A2(new_n827_), .A3(new_n823_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n827_), .B1(new_n826_), .B2(new_n823_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n825_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT122), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT122), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n825_), .B(new_n832_), .C1(new_n828_), .C2(new_n829_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(G1340gat));
  INV_X1    g633(.A(new_n816_), .ZN(new_n835_));
  INV_X1    g634(.A(G120gat), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n836_), .A2(KEYINPUT60), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n591_), .B2(KEYINPUT60), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT123), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n837_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n835_), .B(new_n840_), .C1(new_n839_), .C2(new_n838_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n822_), .ZN(new_n842_));
  AOI211_X1 g641(.A(new_n591_), .B(new_n842_), .C1(new_n816_), .C2(KEYINPUT59), .ZN(new_n843_));
  OAI21_X1  g642(.A(G120gat), .B1(new_n843_), .B2(KEYINPUT124), .ZN(new_n844_));
  AND4_X1   g643(.A1(KEYINPUT124), .A2(new_n817_), .A3(new_n635_), .A4(new_n822_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n841_), .B1(new_n844_), .B2(new_n845_), .ZN(G1341gat));
  INV_X1    g645(.A(G127gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n835_), .A2(new_n847_), .A3(new_n570_), .ZN(new_n848_));
  AOI211_X1 g647(.A(new_n606_), .B(new_n842_), .C1(new_n816_), .C2(KEYINPUT59), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(new_n847_), .ZN(G1342gat));
  INV_X1    g649(.A(G134gat), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n835_), .A2(new_n851_), .A3(new_n536_), .ZN(new_n852_));
  AOI211_X1 g651(.A(new_n656_), .B(new_n842_), .C1(new_n816_), .C2(KEYINPUT59), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n851_), .ZN(G1343gat));
  INV_X1    g653(.A(new_n389_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n811_), .A2(new_n855_), .A3(new_n812_), .A4(new_n813_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n856_), .A2(new_n478_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(new_n296_), .ZN(G1344gat));
  NOR2_X1   g657(.A1(new_n856_), .A2(new_n591_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(new_n297_), .ZN(G1345gat));
  XNOR2_X1  g659(.A(KEYINPUT61), .B(G155gat), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT125), .B1(new_n856_), .B2(new_n606_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n856_), .A2(KEYINPUT125), .A3(new_n606_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n862_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n865_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(new_n863_), .A3(new_n861_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n868_), .ZN(G1346gat));
  OAI21_X1  g668(.A(G162gat), .B1(new_n856_), .B2(new_n656_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n536_), .A2(new_n291_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n856_), .B2(new_n871_), .ZN(G1347gat));
  NOR2_X1   g671(.A1(new_n614_), .A2(new_n603_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n401_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n874_), .A2(new_n632_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n820_), .A2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n604_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(G169gat), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(KEYINPUT126), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n876_), .A2(new_n604_), .A3(new_n253_), .ZN(new_n882_));
  OR2_X1    g681(.A1(new_n878_), .A2(KEYINPUT126), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n878_), .A2(KEYINPUT126), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n883_), .A2(KEYINPUT62), .A3(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n881_), .A2(new_n882_), .A3(new_n885_), .ZN(G1348gat));
  AOI21_X1  g685(.A(G176gat), .B1(new_n876_), .B2(new_n635_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n811_), .A2(new_n812_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n888_), .A2(new_n632_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n874_), .A2(new_n217_), .A3(new_n591_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n887_), .B1(new_n889_), .B2(new_n890_), .ZN(G1349gat));
  INV_X1    g690(.A(new_n876_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n892_), .A2(new_n259_), .A3(new_n606_), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n889_), .A2(new_n401_), .A3(new_n570_), .A4(new_n873_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n893_), .B1(new_n894_), .B2(new_n208_), .ZN(G1350gat));
  OAI21_X1  g694(.A(G190gat), .B1(new_n892_), .B2(new_n656_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n876_), .A2(new_n220_), .A3(new_n536_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1351gat));
  NOR2_X1   g697(.A1(new_n888_), .A2(new_n389_), .ZN(new_n899_));
  AND2_X1   g698(.A1(new_n899_), .A2(new_n873_), .ZN(new_n900_));
  AOI21_X1  g699(.A(G197gat), .B1(new_n900_), .B2(new_n604_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n873_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n902_), .A2(new_n239_), .A3(new_n478_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n901_), .A2(new_n903_), .ZN(G1352gat));
  NAND3_X1  g703(.A1(new_n900_), .A2(new_n241_), .A3(new_n635_), .ZN(new_n905_));
  OAI21_X1  g704(.A(G204gat), .B1(new_n902_), .B2(new_n591_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1353gat));
  XOR2_X1   g706(.A(KEYINPUT63), .B(G211gat), .Z(new_n908_));
  NAND3_X1  g707(.A1(new_n900_), .A2(new_n570_), .A3(new_n908_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n910_), .B1(new_n902_), .B2(new_n606_), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n909_), .A2(new_n911_), .ZN(G1354gat));
  NAND3_X1  g711(.A1(new_n900_), .A2(KEYINPUT127), .A3(new_n536_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n899_), .A2(new_n536_), .A3(new_n873_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT127), .ZN(new_n915_));
  AOI21_X1  g714(.A(G218gat), .B1(new_n914_), .B2(new_n915_), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n650_), .A2(G218gat), .ZN(new_n917_));
  AOI22_X1  g716(.A1(new_n913_), .A2(new_n916_), .B1(new_n900_), .B2(new_n917_), .ZN(G1355gat));
endmodule


