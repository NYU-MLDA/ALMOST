//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 1 1 1 0 1 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 0 0 0 0 0 0 1 0 0 1 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n863_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n899_, new_n900_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(KEYINPUT36), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G29gat), .B(G36gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT70), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G43gat), .B(G50gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT15), .ZN(new_n210_));
  XOR2_X1   g009(.A(G85gat), .B(G92gat), .Z(new_n211_));
  NOR2_X1   g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT7), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT6), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n215_), .B(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n211_), .B1(new_n214_), .B2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n218_), .B(KEYINPUT8), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n217_), .B1(KEYINPUT9), .B2(new_n211_), .ZN(new_n220_));
  XOR2_X1   g019(.A(KEYINPUT10), .B(G99gat), .Z(new_n221_));
  INV_X1    g020(.A(G106gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT65), .B(G92gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT9), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(new_n225_), .A3(G85gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n220_), .A2(new_n223_), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n219_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n210_), .A2(new_n228_), .ZN(new_n229_));
  XOR2_X1   g028(.A(new_n207_), .B(new_n208_), .Z(new_n230_));
  OAI21_X1  g029(.A(new_n229_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT71), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G232gat), .A2(G233gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n231_), .A2(new_n232_), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n204_), .A2(KEYINPUT36), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n236_), .B(new_n237_), .C1(KEYINPUT35), .C2(new_n231_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n235_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n205_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n231_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT35), .ZN(new_n242_));
  AOI22_X1  g041(.A1(new_n241_), .A2(new_n242_), .B1(KEYINPUT36), .B2(new_n204_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n239_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n205_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .A4(new_n236_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n240_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT37), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n240_), .A2(KEYINPUT37), .A3(new_n246_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(G71gat), .B(G78gat), .Z(new_n252_));
  XNOR2_X1  g051(.A(G57gat), .B(G64gat), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n252_), .B1(KEYINPUT11), .B2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT66), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(KEYINPUT11), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n254_), .A2(KEYINPUT66), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n254_), .A2(KEYINPUT66), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n258_), .A2(KEYINPUT11), .A3(new_n253_), .A4(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT73), .ZN(new_n262_));
  XOR2_X1   g061(.A(KEYINPUT72), .B(G1gat), .Z(new_n263_));
  INV_X1    g062(.A(G8gat), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT14), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G15gat), .B(G22gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G1gat), .B(G8gat), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n265_), .A2(new_n266_), .A3(new_n268_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G231gat), .A2(G233gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n262_), .B(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT17), .ZN(new_n276_));
  XOR2_X1   g075(.A(G127gat), .B(G155gat), .Z(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G183gat), .B(G211gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  OR3_X1    g080(.A1(new_n275_), .A2(new_n276_), .A3(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(KEYINPUT17), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n275_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n251_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT75), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  OR3_X1    g087(.A1(KEYINPUT80), .A2(G169gat), .A3(G176gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT80), .B1(G169gat), .B2(G176gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n289_), .A2(KEYINPUT24), .A3(new_n290_), .A4(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT24), .ZN(new_n293_));
  INV_X1    g092(.A(new_n290_), .ZN(new_n294_));
  NOR3_X1   g093(.A1(KEYINPUT80), .A2(G169gat), .A3(G176gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n293_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT23), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT23), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n299_), .A2(G183gat), .A3(G190gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  AND3_X1   g100(.A1(new_n292_), .A2(new_n296_), .A3(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT25), .B(G183gat), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT26), .ZN(new_n304_));
  INV_X1    g103(.A(G190gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT78), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT78), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(G190gat), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n304_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n310_));
  OAI211_X1 g109(.A(KEYINPUT79), .B(new_n303_), .C1(new_n309_), .C2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n310_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT78), .B(G190gat), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n313_), .B1(new_n314_), .B2(new_n304_), .ZN(new_n315_));
  AOI21_X1  g114(.A(KEYINPUT79), .B1(new_n315_), .B2(new_n303_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n302_), .B1(new_n312_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(G183gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n314_), .A2(new_n318_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n299_), .A2(KEYINPUT82), .A3(G183gat), .A4(G190gat), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT82), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n298_), .A2(new_n300_), .A3(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n319_), .A2(new_n320_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT83), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n319_), .A2(KEYINPUT83), .A3(new_n320_), .A4(new_n322_), .ZN(new_n326_));
  INV_X1    g125(.A(G169gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT22), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT22), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(G169gat), .ZN(new_n330_));
  AOI21_X1  g129(.A(KEYINPUT81), .B1(new_n328_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(G176gat), .B1(new_n328_), .B2(KEYINPUT81), .ZN(new_n333_));
  AOI22_X1  g132(.A1(new_n332_), .A2(new_n333_), .B1(G169gat), .B2(G176gat), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n325_), .A2(new_n326_), .A3(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n317_), .A2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT85), .B(G43gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT31), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G71gat), .B(G99gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT86), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(G15gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G227gat), .A2(G233gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT84), .B(KEYINPUT30), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n346_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G127gat), .B(G134gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G113gat), .B(G120gat), .Z(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT87), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G113gat), .B(G120gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n349_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n352_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n349_), .A2(new_n354_), .A3(KEYINPUT87), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n347_), .A2(new_n348_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n358_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n340_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n361_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(new_n339_), .A3(new_n359_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G155gat), .A2(G162gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT1), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT88), .ZN(new_n368_));
  NOR2_X1   g167(.A1(G155gat), .A2(G162gat), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT88), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n366_), .A2(new_n371_), .A3(KEYINPUT1), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n366_), .A2(KEYINPUT1), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n368_), .A2(new_n370_), .A3(new_n372_), .A4(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G141gat), .A2(G148gat), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(G141gat), .A2(G148gat), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n374_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n352_), .A2(new_n355_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT3), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n377_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT2), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n375_), .A2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n382_), .A2(new_n384_), .A3(new_n385_), .A4(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n387_), .A2(new_n370_), .A3(new_n366_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n379_), .A2(new_n380_), .A3(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT99), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n379_), .A2(new_n388_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n358_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT99), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n379_), .A2(new_n380_), .A3(new_n393_), .A4(new_n388_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n390_), .A2(new_n392_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G225gat), .A2(G233gat), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(KEYINPUT4), .B1(new_n358_), .B2(new_n391_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n399_), .B1(new_n395_), .B2(KEYINPUT4), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n398_), .B1(new_n400_), .B2(new_n396_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G1gat), .B(G29gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(G85gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT0), .B(G57gat), .ZN(new_n404_));
  XOR2_X1   g203(.A(new_n403_), .B(new_n404_), .Z(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n401_), .A2(new_n406_), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n398_), .B(new_n405_), .C1(new_n400_), .C2(new_n396_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n365_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT102), .B(KEYINPUT27), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G226gat), .A2(G233gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT19), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT20), .ZN(new_n418_));
  NOR2_X1   g217(.A1(G197gat), .A2(G204gat), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT90), .B(G197gat), .ZN(new_n421_));
  INV_X1    g220(.A(G204gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n420_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G211gat), .B(G218gat), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT21), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n424_), .A2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT91), .B1(new_n422_), .B2(G197gat), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n430_), .B1(new_n421_), .B2(G204gat), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT91), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT90), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n433_), .A2(G197gat), .ZN(new_n434_));
  INV_X1    g233(.A(G197gat), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n435_), .A2(KEYINPUT90), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n432_), .B(new_n422_), .C1(new_n434_), .C2(new_n436_), .ZN(new_n437_));
  AND3_X1   g236(.A1(new_n431_), .A2(KEYINPUT21), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n435_), .A2(KEYINPUT90), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n433_), .A2(G197gat), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n422_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n426_), .B1(new_n441_), .B2(new_n419_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(new_n425_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n428_), .B1(new_n438_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT92), .ZN(new_n445_));
  INV_X1    g244(.A(new_n425_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n446_), .B1(new_n423_), .B2(new_n426_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n431_), .A2(KEYINPUT21), .A3(new_n437_), .ZN(new_n448_));
  AOI22_X1  g247(.A1(new_n447_), .A2(new_n448_), .B1(new_n424_), .B2(new_n427_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT92), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n445_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n336_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n418_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n322_), .A2(new_n320_), .ZN(new_n455_));
  AOI21_X1  g254(.A(KEYINPUT24), .B1(new_n289_), .B2(new_n290_), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT95), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT95), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n296_), .A2(new_n458_), .A3(new_n320_), .A4(new_n322_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT26), .B(G190gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n303_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n292_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n460_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n328_), .A2(new_n330_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(G176gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n301_), .B1(G183gat), .B2(G190gat), .ZN(new_n470_));
  XOR2_X1   g269(.A(new_n291_), .B(KEYINPUT96), .Z(new_n471_));
  NAND3_X1  g270(.A1(new_n469_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n465_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(new_n444_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n417_), .B1(new_n454_), .B2(new_n474_), .ZN(new_n475_));
  OAI211_X1 g274(.A(KEYINPUT20), .B(new_n417_), .C1(new_n473_), .C2(new_n444_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n445_), .A2(new_n336_), .A3(new_n451_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT97), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n445_), .A2(new_n336_), .A3(new_n451_), .A4(KEYINPUT97), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n476_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(G8gat), .B(G36gat), .Z(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G64gat), .B(G92gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NOR3_X1   g286(.A1(new_n475_), .A2(new_n481_), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n476_), .ZN(new_n489_));
  AOI221_X4 g288(.A(KEYINPUT92), .B1(new_n424_), .B2(new_n427_), .C1(new_n447_), .C2(new_n448_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n447_), .A2(new_n448_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n450_), .B1(new_n491_), .B2(new_n428_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(KEYINPUT97), .B1(new_n493_), .B2(new_n336_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n480_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n489_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n474_), .B(KEYINPUT20), .C1(new_n493_), .C2(new_n336_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(new_n416_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n486_), .B1(new_n496_), .B2(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n414_), .B1(new_n488_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT103), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n487_), .B1(new_n475_), .B2(new_n481_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n496_), .A2(new_n498_), .A3(new_n486_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n505_), .A2(KEYINPUT103), .A3(new_n414_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n465_), .A2(KEYINPUT100), .A3(new_n472_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT100), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n463_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n472_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n508_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT94), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n444_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n449_), .A2(KEYINPUT94), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n507_), .A2(new_n511_), .A3(new_n513_), .A4(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT20), .ZN(new_n516_));
  AOI22_X1  g315(.A1(new_n516_), .A2(KEYINPUT101), .B1(new_n479_), .B2(new_n480_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT101), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n515_), .A2(new_n518_), .A3(KEYINPUT20), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n417_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n497_), .A2(new_n416_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n487_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n504_), .A2(KEYINPUT27), .ZN(new_n523_));
  AOI22_X1  g322(.A1(new_n502_), .A2(new_n506_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G78gat), .B(G106gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G22gat), .B(G50gat), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n525_), .B(new_n526_), .Z(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n513_), .A2(new_n514_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT93), .B(KEYINPUT29), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n530_), .B1(new_n379_), .B2(new_n388_), .ZN(new_n531_));
  OAI211_X1 g330(.A(G228gat), .B(G233gat), .C1(new_n529_), .C2(new_n531_), .ZN(new_n532_));
  OR2_X1    g331(.A1(new_n391_), .A2(KEYINPUT29), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT28), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G228gat), .A2(G233gat), .ZN(new_n535_));
  AOI21_X1  g334(.A(KEYINPUT89), .B1(new_n391_), .B2(KEYINPUT29), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n391_), .A2(KEYINPUT89), .A3(KEYINPUT29), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n493_), .B(new_n535_), .C1(new_n536_), .C2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n532_), .A2(new_n534_), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n534_), .B1(new_n532_), .B2(new_n538_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n528_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n532_), .A2(new_n538_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n534_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n545_), .A2(new_n539_), .A3(new_n527_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n542_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n412_), .A2(new_n524_), .A3(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n475_), .A2(new_n481_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n486_), .A2(KEYINPUT32), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n550_), .A2(new_n551_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n516_), .A2(KEYINPUT101), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n479_), .A2(new_n480_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n553_), .A2(new_n519_), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n521_), .B1(new_n555_), .B2(new_n416_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n552_), .B1(new_n556_), .B2(new_n551_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n408_), .B(KEYINPUT33), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n395_), .A2(new_n396_), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n559_), .B(new_n406_), .C1(new_n400_), .C2(new_n397_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n558_), .A2(new_n504_), .A3(new_n503_), .A4(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n547_), .B1(new_n557_), .B2(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n409_), .B1(new_n542_), .B2(new_n546_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n562_), .B1(new_n524_), .B2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n549_), .B1(new_n564_), .B2(new_n365_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n261_), .A2(new_n228_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n261_), .A2(new_n228_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n567_), .B1(new_n568_), .B2(KEYINPUT12), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G230gat), .A2(G233gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT64), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n261_), .A2(new_n228_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT12), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n573_), .A2(KEYINPUT68), .A3(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(KEYINPUT68), .B1(new_n573_), .B2(new_n574_), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n569_), .B(new_n572_), .C1(new_n575_), .C2(new_n576_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n261_), .A2(new_n228_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT67), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n578_), .A2(new_n579_), .A3(new_n573_), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n580_), .B(new_n571_), .C1(new_n579_), .C2(new_n578_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n577_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G120gat), .B(G148gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT5), .ZN(new_n584_));
  XOR2_X1   g383(.A(G176gat), .B(G204gat), .Z(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n582_), .A2(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n586_), .B(KEYINPUT69), .Z(new_n588_));
  AOI21_X1  g387(.A(new_n588_), .B1(new_n577_), .B2(new_n581_), .ZN(new_n589_));
  OR3_X1    g388(.A1(new_n587_), .A2(KEYINPUT13), .A3(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(KEYINPUT13), .B1(new_n587_), .B2(new_n589_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G229gat), .A2(G233gat), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT76), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n230_), .A2(new_n594_), .A3(new_n272_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n594_), .B1(new_n230_), .B2(new_n272_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n210_), .A2(new_n272_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n593_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n596_), .A2(new_n597_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n209_), .A2(new_n271_), .A3(new_n270_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n600_), .B1(new_n603_), .B2(new_n593_), .ZN(new_n604_));
  XOR2_X1   g403(.A(G113gat), .B(G141gat), .Z(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT77), .ZN(new_n606_));
  XOR2_X1   g405(.A(G169gat), .B(G197gat), .Z(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n604_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n604_), .A2(new_n609_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n592_), .A2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n566_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n288_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT104), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n409_), .A2(new_n263_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT105), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT38), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT105), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n618_), .B(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(KEYINPUT38), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT106), .ZN(new_n625_));
  INV_X1    g424(.A(new_n247_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n625_), .B1(new_n566_), .B2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n565_), .A2(KEYINPUT106), .A3(new_n247_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n613_), .A2(new_n285_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G1gat), .B1(new_n632_), .B2(new_n410_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n621_), .A2(new_n624_), .A3(new_n633_), .ZN(G1324gat));
  INV_X1    g433(.A(new_n524_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n616_), .A2(new_n264_), .A3(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n629_), .A2(new_n635_), .A3(new_n630_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT39), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n637_), .A2(new_n638_), .A3(G8gat), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n638_), .B1(new_n637_), .B2(G8gat), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n636_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT40), .Z(G1325gat));
  AND2_X1   g441(.A1(new_n362_), .A2(new_n364_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n615_), .A2(G15gat), .A3(new_n643_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT107), .Z(new_n645_));
  INV_X1    g444(.A(G15gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n646_), .B1(new_n631_), .B2(new_n365_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT41), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n648_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n645_), .A2(new_n649_), .A3(new_n650_), .ZN(G1326gat));
  OR3_X1    g450(.A1(new_n615_), .A2(G22gat), .A3(new_n548_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n631_), .A2(new_n547_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(KEYINPUT108), .B(KEYINPUT42), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n653_), .A2(G22gat), .A3(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n654_), .B1(new_n653_), .B2(G22gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n652_), .B1(new_n655_), .B2(new_n656_), .ZN(G1327gat));
  INV_X1    g456(.A(new_n285_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n658_), .A2(new_n247_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n614_), .A2(new_n659_), .ZN(new_n660_));
  OR3_X1    g459(.A1(new_n660_), .A2(G29gat), .A3(new_n410_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n613_), .A2(new_n658_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT43), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n663_), .B1(new_n565_), .B2(new_n251_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n557_), .A2(new_n561_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(new_n548_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n523_), .B1(new_n556_), .B2(new_n486_), .ZN(new_n667_));
  AOI21_X1  g466(.A(KEYINPUT103), .B1(new_n505_), .B2(new_n414_), .ZN(new_n668_));
  AOI211_X1 g467(.A(new_n501_), .B(new_n413_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n669_));
  OAI211_X1 g468(.A(new_n563_), .B(new_n667_), .C1(new_n668_), .C2(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n365_), .B1(new_n666_), .B2(new_n670_), .ZN(new_n671_));
  OAI211_X1 g470(.A(new_n548_), .B(new_n667_), .C1(new_n668_), .C2(new_n669_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n672_), .A2(new_n411_), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n663_), .B(new_n251_), .C1(new_n671_), .C2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n662_), .B1(new_n664_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT109), .ZN(new_n679_));
  OAI211_X1 g478(.A(KEYINPUT44), .B(new_n662_), .C1(new_n664_), .C2(new_n675_), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n678_), .A2(new_n679_), .A3(new_n409_), .A4(new_n680_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n681_), .A2(G29gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n678_), .A2(new_n409_), .A3(new_n680_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT109), .ZN(new_n684_));
  AOI21_X1  g483(.A(KEYINPUT110), .B1(new_n682_), .B2(new_n684_), .ZN(new_n685_));
  AND4_X1   g484(.A1(KEYINPUT110), .A2(new_n684_), .A3(G29gat), .A4(new_n681_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n661_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT111), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT111), .ZN(new_n689_));
  OAI211_X1 g488(.A(new_n689_), .B(new_n661_), .C1(new_n685_), .C2(new_n686_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(G1328gat));
  NOR3_X1   g490(.A1(new_n660_), .A2(G36gat), .A3(new_n524_), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT45), .Z(new_n693_));
  NAND2_X1  g492(.A1(new_n678_), .A2(new_n680_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G36gat), .B1(new_n694_), .B2(new_n524_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT46), .Z(G1329gat));
  NAND2_X1  g496(.A1(new_n365_), .A2(G43gat), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n660_), .A2(new_n643_), .ZN(new_n699_));
  OAI22_X1  g498(.A1(new_n694_), .A2(new_n698_), .B1(G43gat), .B2(new_n699_), .ZN(new_n700_));
  XOR2_X1   g499(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n701_));
  XNOR2_X1  g500(.A(new_n700_), .B(new_n701_), .ZN(G1330gat));
  OAI21_X1  g501(.A(G50gat), .B1(new_n694_), .B2(new_n548_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n548_), .A2(G50gat), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT113), .Z(new_n705_));
  OAI21_X1  g504(.A(new_n703_), .B1(new_n660_), .B2(new_n705_), .ZN(G1331gat));
  NOR3_X1   g505(.A1(new_n592_), .A2(new_n285_), .A3(new_n612_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n629_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n709_), .A2(G57gat), .A3(new_n409_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n710_), .A2(KEYINPUT114), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(KEYINPUT114), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n566_), .A2(new_n612_), .A3(new_n592_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n288_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(G57gat), .B1(new_n715_), .B2(new_n409_), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n711_), .A2(new_n712_), .A3(new_n716_), .ZN(G1332gat));
  OR3_X1    g516(.A1(new_n714_), .A2(G64gat), .A3(new_n524_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n709_), .A2(new_n635_), .ZN(new_n719_));
  XOR2_X1   g518(.A(KEYINPUT115), .B(KEYINPUT48), .Z(new_n720_));
  AND3_X1   g519(.A1(new_n719_), .A2(G64gat), .A3(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n719_), .B2(G64gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n718_), .B1(new_n721_), .B2(new_n722_), .ZN(G1333gat));
  OR3_X1    g522(.A1(new_n714_), .A2(G71gat), .A3(new_n643_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n709_), .A2(new_n365_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT49), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n725_), .A2(new_n726_), .A3(G71gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n725_), .B2(G71gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n724_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT116), .ZN(G1334gat));
  INV_X1    g529(.A(G78gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n715_), .A2(new_n731_), .A3(new_n547_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT50), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n709_), .A2(new_n547_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n734_), .B2(G78gat), .ZN(new_n735_));
  AOI211_X1 g534(.A(KEYINPUT50), .B(new_n731_), .C1(new_n709_), .C2(new_n547_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n732_), .B1(new_n735_), .B2(new_n736_), .ZN(G1335gat));
  NAND2_X1  g536(.A1(new_n713_), .A2(new_n659_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(G85gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(new_n740_), .A3(new_n409_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n664_), .A2(new_n675_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n592_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n612_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(new_n285_), .A3(new_n744_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n742_), .A2(new_n745_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT117), .Z(new_n747_));
  AND2_X1   g546(.A1(new_n747_), .A2(new_n409_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n741_), .B1(new_n748_), .B2(new_n740_), .ZN(G1336gat));
  AOI21_X1  g548(.A(G92gat), .B1(new_n739_), .B2(new_n635_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n635_), .A2(new_n224_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n747_), .B2(new_n751_), .ZN(G1337gat));
  NAND2_X1  g551(.A1(new_n746_), .A2(new_n365_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(G99gat), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT118), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n753_), .A2(KEYINPUT118), .A3(G99gat), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n365_), .A2(new_n221_), .ZN(new_n758_));
  AOI22_X1  g557(.A1(new_n756_), .A2(new_n757_), .B1(new_n739_), .B2(new_n758_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(KEYINPUT119), .B(KEYINPUT51), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n759_), .B(new_n760_), .Z(G1338gat));
  NAND3_X1  g560(.A1(new_n739_), .A2(new_n222_), .A3(new_n547_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n746_), .A2(new_n547_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n764_), .B2(G106gat), .ZN(new_n765_));
  AOI211_X1 g564(.A(KEYINPUT52), .B(new_n222_), .C1(new_n746_), .C2(new_n547_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n762_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g567(.A1(new_n365_), .A2(new_n409_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n672_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n598_), .A2(new_n599_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n593_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n609_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n603_), .A2(new_n593_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n611_), .A2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(KEYINPUT120), .B1(new_n777_), .B2(new_n587_), .ZN(new_n778_));
  OR2_X1    g577(.A1(new_n582_), .A2(new_n586_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT120), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n779_), .A2(new_n780_), .A3(new_n611_), .A4(new_n776_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n778_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n569_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n784_), .B2(new_n571_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n577_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n785_), .B(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n588_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT56), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n785_), .A2(new_n786_), .ZN(new_n790_));
  NOR3_X1   g589(.A1(new_n784_), .A2(new_n783_), .A3(new_n571_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n788_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT56), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n782_), .B1(new_n789_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT58), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n251_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT121), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n787_), .A2(KEYINPUT56), .A3(new_n788_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n792_), .A2(new_n793_), .ZN(new_n801_));
  AOI22_X1  g600(.A1(new_n800_), .A2(new_n801_), .B1(new_n778_), .B2(new_n781_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT58), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT121), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n804_), .B(new_n251_), .C1(new_n802_), .C2(KEYINPUT58), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n799_), .A2(new_n803_), .A3(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n612_), .A2(new_n779_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n587_), .A2(new_n589_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n809_), .A2(new_n777_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n247_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(KEYINPUT57), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n658_), .B1(new_n806_), .B2(new_n812_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n249_), .A2(new_n250_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n612_), .A2(new_n285_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n814_), .A2(new_n592_), .A3(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n816_), .B(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(KEYINPUT122), .B1(new_n813_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT57), .ZN(new_n820_));
  OR2_X1    g619(.A1(new_n811_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n811_), .A2(new_n820_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n804_), .B1(new_n797_), .B2(new_n251_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n805_), .A2(new_n803_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n821_), .B(new_n822_), .C1(new_n823_), .C2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n285_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT122), .ZN(new_n827_));
  INV_X1    g626(.A(new_n818_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n826_), .A2(new_n827_), .A3(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n771_), .B1(new_n819_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(G113gat), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n830_), .A2(new_n831_), .A3(new_n612_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n826_), .A2(new_n828_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n771_), .A2(KEYINPUT59), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT59), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n612_), .B(new_n835_), .C1(new_n830_), .C2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n832_), .B1(new_n838_), .B2(new_n831_), .ZN(G1340gat));
  INV_X1    g638(.A(G120gat), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n592_), .B2(KEYINPUT60), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n830_), .B(new_n841_), .C1(KEYINPUT60), .C2(new_n840_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n743_), .B(new_n835_), .C1(new_n830_), .C2(new_n836_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n842_), .B1(new_n844_), .B2(new_n840_), .ZN(G1341gat));
  INV_X1    g644(.A(G127gat), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n830_), .A2(new_n846_), .A3(new_n658_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n658_), .B(new_n835_), .C1(new_n830_), .C2(new_n836_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n847_), .B1(new_n849_), .B2(new_n846_), .ZN(G1342gat));
  AOI21_X1  g649(.A(G134gat), .B1(new_n830_), .B2(new_n626_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n830_), .ZN(new_n852_));
  AOI22_X1  g651(.A1(new_n852_), .A2(KEYINPUT59), .B1(new_n833_), .B2(new_n834_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n251_), .A2(G134gat), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(KEYINPUT123), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n851_), .B1(new_n853_), .B2(new_n855_), .ZN(G1343gat));
  NAND2_X1  g655(.A1(new_n819_), .A2(new_n829_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n548_), .A2(new_n365_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n524_), .A2(new_n858_), .A3(new_n409_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n857_), .A2(new_n612_), .A3(new_n860_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g661(.A1(new_n857_), .A2(new_n743_), .A3(new_n860_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G148gat), .ZN(G1345gat));
  AOI21_X1  g663(.A(new_n827_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n865_));
  AOI211_X1 g664(.A(KEYINPUT122), .B(new_n818_), .C1(new_n825_), .C2(new_n285_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n658_), .B(new_n860_), .C1(new_n865_), .C2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(KEYINPUT124), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT124), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n857_), .A2(new_n869_), .A3(new_n658_), .A4(new_n860_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(KEYINPUT61), .B(G155gat), .ZN(new_n871_));
  AND3_X1   g670(.A1(new_n868_), .A2(new_n870_), .A3(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n871_), .B1(new_n868_), .B2(new_n870_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n872_), .A2(new_n873_), .ZN(G1346gat));
  INV_X1    g673(.A(G162gat), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n857_), .A2(new_n875_), .A3(new_n626_), .A4(new_n860_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n857_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n877_), .A2(new_n814_), .A3(new_n859_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n876_), .B1(new_n878_), .B2(new_n875_), .ZN(G1347gat));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n635_), .A2(new_n412_), .ZN(new_n881_));
  XOR2_X1   g680(.A(new_n881_), .B(KEYINPUT125), .Z(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n833_), .A2(new_n548_), .A3(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n744_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n880_), .B1(new_n885_), .B2(new_n327_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n467_), .ZN(new_n887_));
  OAI211_X1 g686(.A(KEYINPUT62), .B(G169gat), .C1(new_n884_), .C2(new_n744_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n886_), .A2(new_n887_), .A3(new_n888_), .ZN(G1348gat));
  OAI21_X1  g688(.A(new_n468_), .B1(new_n884_), .B2(new_n592_), .ZN(new_n890_));
  OR2_X1    g689(.A1(new_n890_), .A2(KEYINPUT126), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(KEYINPUT126), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n877_), .A2(new_n547_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n882_), .A2(new_n468_), .A3(new_n592_), .ZN(new_n894_));
  AOI22_X1  g693(.A1(new_n891_), .A2(new_n892_), .B1(new_n893_), .B2(new_n894_), .ZN(G1349gat));
  NOR3_X1   g694(.A1(new_n884_), .A2(new_n285_), .A3(new_n303_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n893_), .A2(new_n658_), .A3(new_n883_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n896_), .B1(new_n897_), .B2(new_n318_), .ZN(G1350gat));
  OAI21_X1  g697(.A(G190gat), .B1(new_n884_), .B2(new_n814_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n626_), .A2(new_n461_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n884_), .B2(new_n900_), .ZN(G1351gat));
  NAND2_X1  g700(.A1(new_n858_), .A2(new_n410_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(KEYINPUT127), .ZN(new_n903_));
  AOI211_X1 g702(.A(new_n524_), .B(new_n903_), .C1(new_n819_), .C2(new_n829_), .ZN(new_n904_));
  AND3_X1   g703(.A1(new_n904_), .A2(G197gat), .A3(new_n612_), .ZN(new_n905_));
  AOI21_X1  g704(.A(G197gat), .B1(new_n904_), .B2(new_n612_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1352gat));
  NAND2_X1  g706(.A1(new_n904_), .A2(new_n743_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(G204gat), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n904_), .A2(new_n422_), .A3(new_n743_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1353gat));
  OR2_X1    g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  NAND2_X1  g711(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n913_));
  AND4_X1   g712(.A1(new_n658_), .A2(new_n904_), .A3(new_n912_), .A4(new_n913_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n912_), .B1(new_n904_), .B2(new_n658_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1354gat));
  INV_X1    g715(.A(G218gat), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n904_), .A2(new_n917_), .A3(new_n626_), .ZN(new_n918_));
  AND2_X1   g717(.A1(new_n904_), .A2(new_n251_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n919_), .B2(new_n917_), .ZN(G1355gat));
endmodule


