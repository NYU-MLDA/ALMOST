//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 0 1 1 0 1 1 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 1 0 0 0 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n643_, new_n644_, new_n645_, new_n647_, new_n648_, new_n649_,
    new_n651_, new_n652_, new_n653_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n833_,
    new_n834_, new_n835_, new_n837_, new_n838_, new_n840_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_;
  XOR2_X1   g000(.A(G197gat), .B(G204gat), .Z(new_n202_));
  NOR2_X1   g001(.A1(new_n202_), .A2(KEYINPUT21), .ZN(new_n203_));
  XOR2_X1   g002(.A(G211gat), .B(G218gat), .Z(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT91), .ZN(new_n206_));
  INV_X1    g005(.A(G204gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n206_), .A2(new_n207_), .A3(G197gat), .ZN(new_n208_));
  OAI211_X1 g007(.A(KEYINPUT21), .B(new_n208_), .C1(new_n202_), .C2(new_n206_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n205_), .A2(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n202_), .A2(new_n204_), .A3(KEYINPUT21), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  AND2_X1   g012(.A1(KEYINPUT89), .A2(G228gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(KEYINPUT89), .A2(G228gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(G233gat), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  XOR2_X1   g015(.A(new_n216_), .B(KEYINPUT90), .Z(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G141gat), .A2(G148gat), .ZN(new_n219_));
  INV_X1    g018(.A(G141gat), .ZN(new_n220_));
  INV_X1    g019(.A(G148gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT1), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT85), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226_));
  XOR2_X1   g025(.A(new_n226_), .B(KEYINPUT84), .Z(new_n227_));
  INV_X1    g026(.A(KEYINPUT86), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n225_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n229_), .B1(KEYINPUT1), .B2(new_n223_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n228_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n219_), .B(new_n222_), .C1(new_n230_), .C2(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(new_n219_), .B(KEYINPUT2), .Z(new_n233_));
  NAND3_X1  g032(.A1(new_n220_), .A2(new_n221_), .A3(KEYINPUT87), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n233_), .B1(KEYINPUT3), .B2(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n235_), .B1(KEYINPUT3), .B2(new_n234_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n236_), .A2(new_n227_), .A3(new_n223_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n232_), .A2(new_n237_), .ZN(new_n238_));
  AOI211_X1 g037(.A(new_n213_), .B(new_n218_), .C1(new_n238_), .C2(KEYINPUT29), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT92), .ZN(new_n240_));
  XOR2_X1   g039(.A(G78gat), .B(G106gat), .Z(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n238_), .A2(KEYINPUT29), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT93), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  XOR2_X1   g044(.A(new_n212_), .B(KEYINPUT94), .Z(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n243_), .A2(new_n244_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n218_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  AND3_X1   g048(.A1(new_n240_), .A2(new_n242_), .A3(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n242_), .B1(new_n240_), .B2(new_n249_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n238_), .A2(KEYINPUT29), .ZN(new_n252_));
  XOR2_X1   g051(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n253_), .B1(new_n238_), .B2(KEYINPUT29), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  XOR2_X1   g056(.A(G22gat), .B(G50gat), .Z(new_n258_));
  AND2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n257_), .A2(new_n258_), .ZN(new_n260_));
  OAI22_X1  g059(.A1(new_n250_), .A2(new_n251_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n240_), .A2(new_n249_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(new_n241_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n259_), .A2(new_n260_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n240_), .A2(new_n242_), .A3(new_n249_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n263_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n261_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G226gat), .A2(G233gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT19), .ZN(new_n269_));
  XOR2_X1   g068(.A(KEYINPUT80), .B(KEYINPUT23), .Z(new_n270_));
  INV_X1    g069(.A(KEYINPUT23), .ZN(new_n271_));
  AND2_X1   g070(.A1(G183gat), .A2(G190gat), .ZN(new_n272_));
  MUX2_X1   g071(.A(new_n270_), .B(new_n271_), .S(new_n272_), .Z(new_n273_));
  OAI21_X1  g072(.A(new_n273_), .B1(G183gat), .B2(G190gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT22), .B(G169gat), .ZN(new_n276_));
  XOR2_X1   g075(.A(new_n276_), .B(KEYINPUT97), .Z(new_n277_));
  OAI211_X1 g076(.A(new_n274_), .B(new_n275_), .C1(G176gat), .C2(new_n277_), .ZN(new_n278_));
  XOR2_X1   g077(.A(KEYINPUT95), .B(KEYINPUT24), .Z(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n275_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT96), .ZN(new_n281_));
  NOR2_X1   g080(.A1(G169gat), .A2(G176gat), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT96), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n279_), .A2(new_n284_), .A3(new_n275_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n281_), .A2(new_n283_), .A3(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n272_), .A2(KEYINPUT23), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n287_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT25), .B(G183gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT26), .B(G190gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n279_), .A2(new_n283_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n286_), .A2(new_n288_), .A3(new_n291_), .A4(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n278_), .A2(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n246_), .A2(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n288_), .B1(G183gat), .B2(G190gat), .ZN(new_n296_));
  INV_X1    g095(.A(G176gat), .ZN(new_n297_));
  INV_X1    g096(.A(G169gat), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT81), .B1(new_n298_), .B2(KEYINPUT22), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n297_), .B(new_n299_), .C1(new_n276_), .C2(KEYINPUT81), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n296_), .A2(new_n275_), .A3(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n283_), .A2(KEYINPUT24), .A3(new_n275_), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n283_), .A2(KEYINPUT24), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n273_), .A2(new_n291_), .A3(new_n302_), .A4(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n301_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n212_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT20), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n269_), .B1(new_n295_), .B2(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n213_), .B1(new_n278_), .B2(new_n293_), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT20), .B1(new_n305_), .B2(new_n212_), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n308_), .B1(new_n269_), .B2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G8gat), .B(G36gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT18), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G64gat), .B(G92gat), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n314_), .B(new_n315_), .Z(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n312_), .A2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n269_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n278_), .A2(new_n213_), .A3(new_n293_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n269_), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n320_), .A2(KEYINPUT20), .A3(new_n321_), .A4(new_n306_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n319_), .A2(new_n316_), .A3(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n318_), .A2(KEYINPUT27), .A3(new_n323_), .ZN(new_n324_));
  OR2_X1    g123(.A1(new_n323_), .A2(KEYINPUT98), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(KEYINPUT98), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n319_), .A2(new_n322_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(new_n317_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n325_), .A2(new_n326_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT27), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n324_), .A2(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n267_), .A2(new_n332_), .ZN(new_n333_));
  XOR2_X1   g132(.A(G1gat), .B(G29gat), .Z(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G57gat), .B(G85gat), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n336_), .B(new_n337_), .Z(new_n338_));
  NAND2_X1  g137(.A1(G225gat), .A2(G233gat), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G127gat), .B(G134gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G113gat), .B(G120gat), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n341_), .B(new_n342_), .Z(new_n343_));
  NAND2_X1  g142(.A1(new_n238_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n343_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n232_), .A2(new_n237_), .A3(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n340_), .B1(new_n344_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n344_), .A2(KEYINPUT4), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n344_), .A2(KEYINPUT4), .A3(new_n346_), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n338_), .B(new_n348_), .C1(new_n351_), .C2(new_n339_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n338_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n339_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n353_), .B1(new_n354_), .B2(new_n347_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n352_), .A2(new_n355_), .A3(KEYINPUT100), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT100), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n357_), .B(new_n353_), .C1(new_n354_), .C2(new_n347_), .ZN(new_n358_));
  AND3_X1   g157(.A1(new_n356_), .A2(KEYINPUT101), .A3(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(KEYINPUT101), .B1(new_n356_), .B2(new_n358_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G71gat), .B(G99gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT83), .ZN(new_n363_));
  XOR2_X1   g162(.A(G15gat), .B(G43gat), .Z(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n305_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(new_n345_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G227gat), .A2(G233gat), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n368_), .B(KEYINPUT82), .Z(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT30), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT31), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n367_), .B(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n333_), .A2(new_n361_), .A3(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n332_), .B1(new_n261_), .B2(new_n266_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n267_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n344_), .A2(new_n340_), .A3(new_n346_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(new_n338_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n378_), .B1(new_n351_), .B2(new_n339_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n329_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT33), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n355_), .A2(new_n381_), .ZN(new_n382_));
  OAI211_X1 g181(.A(KEYINPUT33), .B(new_n353_), .C1(new_n354_), .C2(new_n347_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n380_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n356_), .A2(new_n358_), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n316_), .A2(KEYINPUT32), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n312_), .A2(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n387_), .B1(new_n386_), .B2(new_n327_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n384_), .B1(new_n385_), .B2(new_n388_), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n361_), .A2(new_n375_), .B1(new_n376_), .B2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n374_), .B1(new_n390_), .B2(new_n373_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT79), .B(G15gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(G22gat), .ZN(new_n393_));
  INV_X1    g192(.A(G1gat), .ZN(new_n394_));
  INV_X1    g193(.A(G8gat), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT14), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n393_), .A2(new_n396_), .ZN(new_n397_));
  XOR2_X1   g196(.A(G1gat), .B(G8gat), .Z(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G29gat), .B(G36gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G43gat), .B(G50gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n399_), .B(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G229gat), .A2(G233gat), .ZN(new_n405_));
  OR2_X1    g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(new_n402_), .B(KEYINPUT15), .Z(new_n407_));
  OR2_X1    g206(.A1(new_n399_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n399_), .A2(new_n402_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(new_n409_), .A3(new_n405_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n406_), .A2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G113gat), .B(G141gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G169gat), .B(G197gat), .ZN(new_n413_));
  XOR2_X1   g212(.A(new_n412_), .B(new_n413_), .Z(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n411_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n406_), .A2(new_n410_), .A3(new_n414_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(G85gat), .A2(G92gat), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  AND2_X1   g219(.A1(G85gat), .A2(G92gat), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n421_), .A2(new_n419_), .ZN(new_n422_));
  AOI21_X1  g221(.A(KEYINPUT9), .B1(new_n422_), .B2(KEYINPUT67), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT67), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT9), .ZN(new_n425_));
  NOR4_X1   g224(.A1(new_n421_), .A2(new_n419_), .A3(new_n424_), .A4(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n420_), .B1(new_n423_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT68), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT68), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n429_), .B(new_n420_), .C1(new_n423_), .C2(new_n426_), .ZN(new_n430_));
  OR2_X1    g229(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(G106gat), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n434_), .A2(KEYINPUT66), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT66), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n437_), .B1(new_n433_), .B2(G106gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G99gat), .A2(G106gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT6), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT6), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n441_), .A2(G99gat), .A3(G106gat), .ZN(new_n442_));
  AOI22_X1  g241(.A1(new_n436_), .A2(new_n438_), .B1(new_n440_), .B2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n428_), .A2(new_n430_), .A3(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G57gat), .B(G64gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT11), .ZN(new_n446_));
  XOR2_X1   g245(.A(G71gat), .B(G78gat), .Z(new_n447_));
  NOR2_X1   g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n446_), .A2(new_n447_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n445_), .A2(KEYINPUT11), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n448_), .B1(new_n449_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(G99gat), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n454_), .A2(new_n435_), .A3(KEYINPUT69), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT7), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n440_), .A2(new_n442_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT7), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n458_), .A2(new_n454_), .A3(new_n435_), .A4(KEYINPUT69), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n456_), .A2(new_n457_), .A3(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(new_n422_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT70), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT70), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n460_), .A2(new_n463_), .A3(new_n422_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n462_), .A2(KEYINPUT8), .A3(new_n464_), .ZN(new_n465_));
  AOI211_X1 g264(.A(new_n463_), .B(KEYINPUT8), .C1(new_n460_), .C2(new_n422_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n444_), .A2(new_n453_), .A3(new_n465_), .A4(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G230gat), .A2(G233gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n468_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT8), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n474_), .B1(new_n461_), .B2(KEYINPUT70), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n466_), .B1(new_n475_), .B2(new_n464_), .ZN(new_n476_));
  AOI211_X1 g275(.A(KEYINPUT12), .B(new_n453_), .C1(new_n476_), .C2(new_n444_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT12), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n444_), .A2(new_n467_), .A3(new_n465_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n478_), .B1(new_n479_), .B2(new_n452_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n473_), .B1(new_n477_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n479_), .A2(new_n452_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n472_), .B1(new_n483_), .B2(new_n468_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G120gat), .B(G148gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT5), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G176gat), .B(G204gat), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n486_), .B(new_n487_), .Z(new_n488_));
  OR3_X1    g287(.A1(new_n482_), .A2(new_n484_), .A3(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n488_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n491_), .A2(KEYINPUT13), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT71), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(KEYINPUT13), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT72), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G232gat), .A2(G233gat), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n498_), .B(KEYINPUT34), .Z(new_n499_));
  XOR2_X1   g298(.A(KEYINPUT73), .B(KEYINPUT35), .Z(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n476_), .A2(new_n402_), .A3(new_n444_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n479_), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n501_), .B(new_n502_), .C1(new_n503_), .C2(new_n407_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n499_), .A2(new_n500_), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n505_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G190gat), .B(G218gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT74), .ZN(new_n509_));
  XOR2_X1   g308(.A(G134gat), .B(G162gat), .Z(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n511_), .A2(KEYINPUT36), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT75), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n506_), .A2(new_n507_), .A3(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n506_), .A2(new_n507_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n511_), .B(KEYINPUT36), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT77), .ZN(new_n517_));
  OAI211_X1 g316(.A(KEYINPUT76), .B(new_n514_), .C1(new_n515_), .C2(new_n517_), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n514_), .A2(KEYINPUT76), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT37), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT78), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n518_), .A2(new_n519_), .A3(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n520_), .A2(KEYINPUT78), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n523_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n399_), .B(new_n453_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G231gat), .A2(G233gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT17), .ZN(new_n531_));
  XOR2_X1   g330(.A(G127gat), .B(G155gat), .Z(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT16), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G183gat), .B(G211gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  OR3_X1    g334(.A1(new_n530_), .A2(new_n531_), .A3(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(KEYINPUT17), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n530_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n526_), .A2(new_n539_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n391_), .A2(new_n418_), .A3(new_n497_), .A4(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT102), .ZN(new_n542_));
  INV_X1    g341(.A(new_n360_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n356_), .A2(KEYINPUT101), .A3(new_n358_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n542_), .A2(new_n394_), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT38), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n375_), .A2(new_n544_), .A3(new_n543_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n376_), .A2(new_n389_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n373_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n333_), .A2(new_n361_), .A3(new_n373_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n518_), .A2(new_n519_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT103), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n497_), .A2(new_n418_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n557_), .A2(new_n539_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(G1gat), .B1(new_n559_), .B2(new_n361_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n546_), .A2(new_n547_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n548_), .A2(new_n560_), .A3(new_n561_), .ZN(G1324gat));
  NAND3_X1  g361(.A1(new_n542_), .A2(new_n395_), .A3(new_n332_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT39), .ZN(new_n564_));
  INV_X1    g363(.A(new_n559_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(new_n332_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n564_), .B1(new_n566_), .B2(G8gat), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n324_), .A2(new_n331_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n564_), .B(G8gat), .C1(new_n559_), .C2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n563_), .B1(new_n567_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT40), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n563_), .B(KEYINPUT40), .C1(new_n567_), .C2(new_n570_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(G1325gat));
  INV_X1    g374(.A(G15gat), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n542_), .A2(new_n576_), .A3(new_n373_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n565_), .A2(new_n373_), .ZN(new_n578_));
  AOI21_X1  g377(.A(KEYINPUT41), .B1(new_n578_), .B2(G15gat), .ZN(new_n579_));
  OAI211_X1 g378(.A(KEYINPUT41), .B(G15gat), .C1(new_n559_), .C2(new_n372_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n577_), .B1(new_n579_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT104), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n577_), .B(KEYINPUT104), .C1(new_n579_), .C2(new_n581_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(G1326gat));
  OAI21_X1  g385(.A(G22gat), .B1(new_n559_), .B2(new_n376_), .ZN(new_n587_));
  XOR2_X1   g386(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(G22gat), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n542_), .A2(new_n590_), .A3(new_n267_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n591_), .ZN(G1327gat));
  INV_X1    g391(.A(new_n497_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n539_), .A2(new_n554_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n391_), .A2(new_n418_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(G29gat), .B1(new_n597_), .B2(new_n545_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n539_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n557_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT43), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n601_), .B(new_n526_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n601_), .B1(new_n391_), .B2(new_n526_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n600_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT44), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  OAI211_X1 g406(.A(KEYINPUT44), .B(new_n600_), .C1(new_n603_), .C2(new_n604_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n545_), .A2(G29gat), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n598_), .B1(new_n609_), .B2(new_n610_), .ZN(G1328gat));
  NAND3_X1  g410(.A1(new_n607_), .A2(new_n332_), .A3(new_n608_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(G36gat), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT46), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT106), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT107), .Z(new_n616_));
  OR2_X1    g415(.A1(new_n568_), .A2(G36gat), .ZN(new_n617_));
  OR3_X1    g416(.A1(new_n596_), .A2(KEYINPUT45), .A3(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(KEYINPUT45), .B1(new_n596_), .B2(new_n617_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n613_), .A2(new_n616_), .A3(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n616_), .B1(new_n613_), .B2(new_n620_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(G1329gat));
  NAND4_X1  g422(.A1(new_n607_), .A2(G43gat), .A3(new_n373_), .A4(new_n608_), .ZN(new_n624_));
  AOI21_X1  g423(.A(G43gat), .B1(new_n597_), .B2(new_n373_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g427(.A1(new_n596_), .A2(G50gat), .A3(new_n376_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n607_), .A2(new_n267_), .A3(new_n608_), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n630_), .A2(KEYINPUT108), .A3(G50gat), .ZN(new_n631_));
  AOI21_X1  g430(.A(KEYINPUT108), .B1(new_n630_), .B2(G50gat), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n629_), .B1(new_n631_), .B2(new_n632_), .ZN(G1331gat));
  INV_X1    g432(.A(new_n418_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n556_), .A2(new_n634_), .A3(new_n593_), .A4(new_n599_), .ZN(new_n635_));
  INV_X1    g434(.A(G57gat), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n635_), .A2(new_n636_), .A3(new_n361_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n553_), .A2(new_n418_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n638_), .A2(new_n593_), .A3(new_n540_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n361_), .B1(new_n639_), .B2(KEYINPUT109), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n640_), .B1(KEYINPUT109), .B2(new_n639_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n637_), .B1(new_n641_), .B2(new_n636_), .ZN(G1332gat));
  OAI21_X1  g441(.A(G64gat), .B1(new_n635_), .B2(new_n568_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT48), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n568_), .A2(G64gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n644_), .B1(new_n639_), .B2(new_n645_), .ZN(G1333gat));
  OAI21_X1  g445(.A(G71gat), .B1(new_n635_), .B2(new_n372_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT49), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n372_), .A2(G71gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n648_), .B1(new_n639_), .B2(new_n649_), .ZN(G1334gat));
  OAI21_X1  g449(.A(G78gat), .B1(new_n635_), .B2(new_n376_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT50), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n376_), .A2(G78gat), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n652_), .B1(new_n639_), .B2(new_n653_), .ZN(G1335gat));
  NOR2_X1   g453(.A1(new_n497_), .A2(new_n594_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n638_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(G85gat), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n657_), .A2(new_n658_), .A3(new_n545_), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n603_), .A2(new_n604_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n497_), .A2(new_n418_), .A3(new_n599_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n662_), .A2(new_n545_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n659_), .B1(new_n663_), .B2(new_n658_), .ZN(G1336gat));
  INV_X1    g463(.A(G92gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n657_), .A2(new_n665_), .A3(new_n332_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n662_), .A2(new_n332_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n666_), .B1(new_n667_), .B2(new_n665_), .ZN(G1337gat));
  INV_X1    g467(.A(KEYINPUT110), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT51), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n656_), .A2(new_n372_), .A3(new_n433_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n662_), .A2(new_n373_), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n670_), .B(new_n672_), .C1(new_n673_), .C2(new_n454_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n454_), .B1(new_n662_), .B2(new_n373_), .ZN(new_n675_));
  OAI211_X1 g474(.A(new_n669_), .B(KEYINPUT51), .C1(new_n675_), .C2(new_n671_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(G1338gat));
  NAND3_X1  g476(.A1(new_n657_), .A2(new_n435_), .A3(new_n267_), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n267_), .B(new_n661_), .C1(new_n603_), .C2(new_n604_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT52), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n679_), .A2(new_n680_), .A3(G106gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n679_), .B2(G106gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n678_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT53), .ZN(G1339gat));
  OAI21_X1  g483(.A(new_n468_), .B1(new_n477_), .B2(new_n480_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n481_), .A2(KEYINPUT55), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT55), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n687_), .B(new_n473_), .C1(new_n477_), .C2(new_n480_), .ZN(new_n688_));
  AOI221_X4 g487(.A(KEYINPUT112), .B1(new_n685_), .B2(new_n471_), .C1(new_n686_), .C2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT112), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n686_), .A2(new_n688_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n685_), .A2(new_n471_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n690_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n488_), .B1(new_n689_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT56), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n488_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n697_), .A2(new_n695_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n698_), .B1(new_n689_), .B2(new_n693_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT114), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n483_), .A2(KEYINPUT12), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n479_), .A2(new_n478_), .A3(new_n452_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n687_), .B1(new_n704_), .B2(new_n473_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n688_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n692_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT112), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n691_), .A2(new_n690_), .A3(new_n692_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n710_), .A2(KEYINPUT114), .A3(new_n698_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n696_), .A2(new_n701_), .A3(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n405_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n408_), .A2(new_n409_), .A3(new_n713_), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n714_), .B(new_n415_), .C1(new_n404_), .C2(new_n713_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n417_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(new_n489_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT113), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n712_), .A2(KEYINPUT58), .A3(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT115), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n712_), .A2(new_n718_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT58), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT115), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n712_), .A2(new_n724_), .A3(KEYINPUT58), .A4(new_n718_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n720_), .A2(new_n723_), .A3(new_n526_), .A4(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n491_), .A2(new_n716_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n697_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n699_), .B1(new_n729_), .B2(KEYINPUT56), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n418_), .A2(new_n489_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n728_), .B1(new_n730_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT57), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n733_), .A2(new_n734_), .A3(new_n554_), .ZN(new_n735_));
  AOI22_X1  g534(.A1(new_n694_), .A2(new_n695_), .B1(new_n710_), .B2(new_n698_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n727_), .B1(new_n736_), .B2(new_n731_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n554_), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT57), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n735_), .A2(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n599_), .B1(new_n726_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n526_), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n742_), .A2(new_n497_), .A3(new_n634_), .A4(new_n599_), .ZN(new_n743_));
  XOR2_X1   g542(.A(KEYINPUT111), .B(KEYINPUT54), .Z(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n540_), .A2(new_n497_), .A3(new_n634_), .A4(new_n744_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n741_), .A2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n333_), .A2(new_n545_), .A3(new_n373_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(G113gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(new_n752_), .A3(new_n418_), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n751_), .A2(KEYINPUT59), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n751_), .A2(KEYINPUT59), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n634_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n753_), .B1(new_n756_), .B2(new_n752_), .ZN(G1340gat));
  INV_X1    g556(.A(G120gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n758_), .B1(new_n497_), .B2(KEYINPUT60), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n751_), .B(new_n759_), .C1(KEYINPUT60), .C2(new_n758_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n497_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(new_n758_), .ZN(G1341gat));
  INV_X1    g561(.A(G127gat), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n751_), .A2(new_n763_), .A3(new_n599_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n539_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(new_n763_), .ZN(G1342gat));
  INV_X1    g565(.A(G134gat), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n751_), .A2(new_n767_), .A3(new_n555_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n742_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n768_), .B1(new_n769_), .B2(new_n767_), .ZN(G1343gat));
  NAND2_X1  g569(.A1(new_n726_), .A2(new_n740_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n539_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n746_), .A2(new_n747_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n545_), .A2(new_n375_), .A3(new_n372_), .ZN(new_n775_));
  XOR2_X1   g574(.A(new_n775_), .B(KEYINPUT116), .Z(new_n776_));
  AND2_X1   g575(.A1(new_n774_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n418_), .ZN(new_n778_));
  XOR2_X1   g577(.A(KEYINPUT117), .B(G141gat), .Z(new_n779_));
  XNOR2_X1  g578(.A(new_n778_), .B(new_n779_), .ZN(G1344gat));
  NAND2_X1  g579(.A1(new_n777_), .A2(new_n593_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g581(.A(KEYINPUT118), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n774_), .A2(new_n783_), .A3(new_n599_), .A4(new_n776_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT119), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n599_), .B(new_n776_), .C1(new_n741_), .C2(new_n748_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT118), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n784_), .A2(new_n785_), .A3(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n785_), .B1(new_n784_), .B2(new_n787_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(KEYINPUT61), .B(G155gat), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n788_), .A2(new_n789_), .A3(new_n791_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n786_), .A2(KEYINPUT118), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n786_), .A2(KEYINPUT118), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT119), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n784_), .A2(new_n787_), .A3(new_n785_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n790_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n792_), .A2(new_n797_), .ZN(G1346gat));
  INV_X1    g597(.A(G162gat), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n777_), .A2(new_n799_), .A3(new_n555_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n777_), .A2(new_n526_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n800_), .B1(new_n802_), .B2(new_n799_), .ZN(G1347gat));
  NAND4_X1  g602(.A1(new_n543_), .A2(new_n544_), .A3(new_n332_), .A4(new_n373_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT120), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n805_), .A2(KEYINPUT121), .A3(new_n418_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT121), .B1(new_n805_), .B2(new_n418_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n376_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(G169gat), .B1(new_n808_), .B2(new_n749_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT123), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n809_), .A2(new_n810_), .A3(KEYINPUT62), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n810_), .B1(new_n809_), .B2(KEYINPUT62), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT62), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n814_), .B(G169gat), .C1(new_n808_), .C2(new_n749_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(KEYINPUT122), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT124), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n805_), .A2(new_n376_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n817_), .B1(new_n749_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n818_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n774_), .A2(KEYINPUT124), .A3(new_n820_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n819_), .A2(new_n821_), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n634_), .A2(new_n277_), .ZN(new_n823_));
  OAI22_X1  g622(.A1(new_n813_), .A2(new_n816_), .B1(new_n822_), .B2(new_n823_), .ZN(G1348gat));
  NOR2_X1   g623(.A1(new_n749_), .A2(new_n818_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(G176gat), .A3(new_n593_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT125), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n828_), .B(new_n297_), .C1(new_n822_), .C2(new_n497_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n497_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n830_));
  OAI21_X1  g629(.A(KEYINPUT125), .B1(new_n830_), .B2(G176gat), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n827_), .B1(new_n829_), .B2(new_n831_), .ZN(G1349gat));
  AOI21_X1  g631(.A(G183gat), .B1(new_n825_), .B2(new_n599_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n822_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n539_), .A2(new_n289_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n833_), .B1(new_n834_), .B2(new_n835_), .ZN(G1350gat));
  OAI21_X1  g635(.A(G190gat), .B1(new_n822_), .B2(new_n742_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n555_), .A2(new_n290_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(new_n822_), .B2(new_n838_), .ZN(G1351gat));
  NAND4_X1  g638(.A1(new_n361_), .A2(new_n267_), .A3(new_n332_), .A4(new_n372_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n749_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n418_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n593_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n845_));
  XOR2_X1   g644(.A(new_n844_), .B(new_n845_), .Z(G1353gat));
  NAND2_X1  g645(.A1(new_n841_), .A2(new_n599_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n848_));
  AND2_X1   g647(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n847_), .A2(new_n848_), .A3(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n850_), .B1(new_n847_), .B2(new_n848_), .ZN(G1354gat));
  NAND2_X1  g650(.A1(new_n841_), .A2(new_n526_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(G218gat), .ZN(new_n853_));
  INV_X1    g652(.A(G218gat), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n841_), .A2(new_n854_), .A3(new_n555_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n853_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT127), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n853_), .A2(KEYINPUT127), .A3(new_n855_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(G1355gat));
endmodule


