//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 1 1 0 1 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_;
  INV_X1    g000(.A(G85gat), .ZN(new_n202_));
  INV_X1    g001(.A(G92gat), .ZN(new_n203_));
  NOR3_X1   g002(.A1(new_n202_), .A2(new_n203_), .A3(KEYINPUT9), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT10), .B(G99gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n205_), .A2(G106gat), .ZN(new_n206_));
  XOR2_X1   g005(.A(G85gat), .B(G92gat), .Z(new_n207_));
  AOI211_X1 g006(.A(new_n204_), .B(new_n206_), .C1(KEYINPUT9), .C2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT65), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT6), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT64), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  AND3_X1   g013(.A1(new_n211_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n214_), .B1(new_n211_), .B2(new_n213_), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n209_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n214_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n210_), .A2(KEYINPUT64), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n218_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n211_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(KEYINPUT65), .A3(new_n222_), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n217_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n208_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT7), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G99gat), .A2(G106gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n228_), .A2(KEYINPUT67), .A3(new_n229_), .A4(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n233_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n217_), .A2(new_n223_), .A3(new_n231_), .A4(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT8), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n207_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n221_), .A2(new_n222_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n241_), .A2(new_n236_), .A3(new_n231_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n238_), .B1(new_n242_), .B2(new_n207_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n240_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  AOI211_X1 g044(.A(KEYINPUT68), .B(new_n238_), .C1(new_n242_), .C2(new_n207_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n225_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G71gat), .B(G78gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G57gat), .B(G64gat), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n248_), .B1(KEYINPUT11), .B2(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n250_), .B1(KEYINPUT11), .B2(new_n249_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n249_), .A2(new_n248_), .A3(KEYINPUT11), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n247_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT12), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n247_), .A2(KEYINPUT12), .A3(new_n254_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n253_), .B(new_n225_), .C1(new_n245_), .C2(new_n246_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT70), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G230gat), .A2(G233gat), .ZN(new_n261_));
  AND3_X1   g060(.A1(new_n259_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n260_), .B1(new_n259_), .B2(new_n261_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n257_), .B(new_n258_), .C1(new_n262_), .C2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n255_), .A2(KEYINPUT69), .A3(new_n259_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n261_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n247_), .A2(new_n267_), .A3(new_n254_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n265_), .A2(new_n266_), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n264_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G120gat), .B(G148gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT72), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT71), .ZN(new_n273_));
  XOR2_X1   g072(.A(G176gat), .B(G204gat), .Z(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT5), .ZN(new_n275_));
  XOR2_X1   g074(.A(new_n273_), .B(new_n275_), .Z(new_n276_));
  NAND2_X1  g075(.A1(new_n270_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n276_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n264_), .A2(new_n269_), .A3(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n277_), .A2(KEYINPUT73), .A3(new_n279_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT74), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT13), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n285_), .A2(new_n286_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n284_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n282_), .A2(KEYINPUT74), .A3(KEYINPUT13), .A4(new_n283_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G226gat), .A2(G233gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT19), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT20), .ZN(new_n296_));
  INV_X1    g095(.A(G183gat), .ZN(new_n297_));
  INV_X1    g096(.A(G190gat), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT23), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT87), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT23), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(G183gat), .A3(G190gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT88), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n300_), .A2(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT86), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT24), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(G169gat), .ZN(new_n310_));
  INV_X1    g109(.A(G176gat), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT24), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n307_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT26), .B(G190gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT25), .B(G183gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n305_), .A2(new_n309_), .A3(new_n313_), .A4(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n299_), .A2(new_n302_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n318_), .B1(G183gat), .B2(G190gat), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n310_), .A2(new_n311_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT22), .B(G169gat), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n320_), .B1(new_n321_), .B2(new_n311_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n319_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n317_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT96), .ZN(new_n326_));
  NOR2_X1   g125(.A1(G211gat), .A2(G218gat), .ZN(new_n327_));
  AND2_X1   g126(.A1(G211gat), .A2(G218gat), .ZN(new_n328_));
  XOR2_X1   g127(.A(G197gat), .B(G204gat), .Z(new_n329_));
  OAI221_X1 g128(.A(new_n326_), .B1(new_n327_), .B2(new_n328_), .C1(new_n329_), .C2(KEYINPUT21), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(KEYINPUT21), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n296_), .B1(new_n325_), .B2(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n305_), .B1(G183gat), .B2(G190gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n322_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n315_), .B(KEYINPUT98), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n314_), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n337_), .A2(new_n318_), .A3(new_n309_), .A4(new_n313_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n335_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n332_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n295_), .B1(new_n333_), .B2(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT20), .B1(new_n339_), .B2(new_n340_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT99), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n344_), .B1(new_n340_), .B2(new_n324_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n340_), .A2(new_n344_), .A3(new_n324_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n343_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n342_), .B1(new_n348_), .B2(new_n295_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G8gat), .B(G36gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(new_n203_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT18), .B(G64gat), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n351_), .B(new_n352_), .Z(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n349_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n349_), .A2(new_n354_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  AND2_X1   g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(G155gat), .A2(G162gat), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(G141gat), .A2(G148gat), .ZN(new_n362_));
  XOR2_X1   g161(.A(new_n362_), .B(KEYINPUT3), .Z(new_n363_));
  NAND2_X1  g162(.A1(G141gat), .A2(G148gat), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n364_), .B(KEYINPUT2), .Z(new_n365_));
  OAI21_X1  g164(.A(new_n361_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT1), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n360_), .B1(new_n359_), .B2(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n368_), .B1(new_n367_), .B2(new_n359_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n362_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n369_), .A2(new_n370_), .A3(new_n364_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n366_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G127gat), .B(G134gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G113gat), .B(G120gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n373_), .A2(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n374_), .A2(new_n375_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT89), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n380_), .B1(new_n376_), .B2(new_n379_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n372_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n377_), .A2(KEYINPUT4), .A3(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT100), .B1(new_n382_), .B2(KEYINPUT4), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT100), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT4), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n381_), .A2(new_n372_), .A3(new_n385_), .A4(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n383_), .A2(new_n384_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G225gat), .A2(G233gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  OR2_X1    g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G1gat), .B(G29gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(new_n202_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT0), .B(G57gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n377_), .A2(new_n382_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n395_), .B1(new_n396_), .B2(new_n390_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n383_), .A2(new_n384_), .A3(new_n390_), .A4(new_n387_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(new_n389_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(new_n399_), .A3(new_n395_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT33), .ZN(new_n401_));
  AOI22_X1  g200(.A1(new_n391_), .A2(new_n397_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n400_), .A2(new_n401_), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n354_), .A2(KEYINPUT32), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n398_), .A2(new_n399_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n395_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  AOI22_X1  g207(.A1(new_n349_), .A2(new_n405_), .B1(new_n408_), .B2(new_n400_), .ZN(new_n409_));
  OR3_X1    g208(.A1(new_n348_), .A2(KEYINPUT101), .A3(new_n295_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n333_), .A2(new_n341_), .A3(new_n295_), .ZN(new_n411_));
  OAI211_X1 g210(.A(KEYINPUT101), .B(new_n411_), .C1(new_n348_), .C2(new_n295_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n410_), .A2(KEYINPUT32), .A3(new_n354_), .A4(new_n412_), .ZN(new_n413_));
  AOI22_X1  g212(.A1(new_n358_), .A2(new_n404_), .B1(new_n409_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT29), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n340_), .B1(new_n415_), .B2(new_n373_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT95), .B(G233gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT94), .B(G228gat), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n416_), .A2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n332_), .B1(KEYINPUT29), .B2(new_n372_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n419_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  XOR2_X1   g222(.A(G78gat), .B(G106gat), .Z(new_n424_));
  AND3_X1   g223(.A1(new_n420_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n424_), .B1(new_n420_), .B2(new_n423_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n420_), .A2(new_n423_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n424_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT97), .ZN(new_n431_));
  XOR2_X1   g230(.A(KEYINPUT91), .B(KEYINPUT93), .Z(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n372_), .A2(KEYINPUT29), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G22gat), .B(G50gat), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n434_), .A2(new_n436_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n433_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n439_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n433_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n441_), .A2(new_n442_), .A3(new_n437_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n432_), .B1(new_n440_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n440_), .A2(new_n443_), .A3(new_n432_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n427_), .A2(new_n431_), .A3(new_n445_), .A4(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT97), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n446_), .B1(new_n426_), .B2(new_n448_), .ZN(new_n449_));
  OAI22_X1  g248(.A1(new_n449_), .A2(new_n444_), .B1(new_n426_), .B2(new_n425_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n447_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT102), .B1(new_n414_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT103), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n410_), .A2(new_n412_), .A3(new_n353_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n355_), .A2(KEYINPUT27), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n454_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n408_), .A2(new_n400_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n451_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT27), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n461_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n455_), .A2(KEYINPUT103), .A3(KEYINPUT27), .A4(new_n355_), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n458_), .A2(new_n460_), .A3(new_n462_), .A4(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n357_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n465_), .A2(new_n402_), .A3(new_n355_), .A4(new_n403_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n413_), .A2(new_n409_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT102), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n468_), .A2(new_n469_), .A3(new_n451_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n453_), .A2(new_n464_), .A3(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G227gat), .A2(G233gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n324_), .B(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G71gat), .B(G99gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(G43gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(KEYINPUT30), .B(G15gat), .Z(new_n476_));
  XOR2_X1   g275(.A(new_n475_), .B(new_n476_), .Z(new_n477_));
  XNOR2_X1  g276(.A(new_n473_), .B(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n381_), .B(KEYINPUT31), .ZN(new_n480_));
  OR3_X1    g279(.A1(new_n479_), .A2(KEYINPUT90), .A3(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n480_), .B(KEYINPUT90), .Z(new_n482_));
  NAND2_X1  g281(.A1(new_n479_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n471_), .A2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n458_), .A2(new_n463_), .A3(new_n462_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n486_), .A2(new_n452_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n484_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n459_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n485_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G169gat), .B(G197gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT85), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G113gat), .B(G141gat), .ZN(new_n494_));
  XOR2_X1   g293(.A(new_n493_), .B(new_n494_), .Z(new_n495_));
  XNOR2_X1  g294(.A(G29gat), .B(G36gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G43gat), .B(G50gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n498_), .B(KEYINPUT15), .Z(new_n499_));
  XOR2_X1   g298(.A(G15gat), .B(G22gat), .Z(new_n500_));
  NAND2_X1  g299(.A1(G1gat), .A2(G8gat), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n500_), .B1(KEYINPUT14), .B2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT81), .ZN(new_n503_));
  XOR2_X1   g302(.A(G1gat), .B(G8gat), .Z(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT81), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n502_), .B(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n504_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n499_), .B1(new_n505_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n505_), .A2(new_n509_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n498_), .ZN(new_n512_));
  OR3_X1    g311(.A1(new_n511_), .A2(KEYINPUT84), .A3(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT84), .B1(new_n511_), .B2(new_n512_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n510_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G229gat), .A2(G233gat), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  AOI22_X1  g316(.A1(new_n513_), .A2(new_n514_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n518_), .A2(new_n516_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n495_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n515_), .A2(new_n516_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n495_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n521_), .B(new_n522_), .C1(new_n516_), .C2(new_n518_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n520_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n491_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT104), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n292_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n524_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n528_), .B1(new_n485_), .B2(new_n490_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT104), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G231gat), .A2(G233gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n511_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(new_n253_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G127gat), .B(G155gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(G211gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT16), .B(G183gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT17), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n539_), .B(KEYINPUT82), .Z(new_n540_));
  NOR2_X1   g339(.A1(new_n534_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT83), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n538_), .A2(KEYINPUT17), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n534_), .A2(new_n539_), .A3(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT75), .ZN(new_n547_));
  INV_X1    g346(.A(G99gat), .ZN(new_n548_));
  INV_X1    g347(.A(G106gat), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n230_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n235_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n552_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n215_), .A2(new_n216_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n207_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT8), .ZN(new_n556_));
  AOI22_X1  g355(.A1(new_n556_), .A2(KEYINPUT68), .B1(new_n237_), .B2(new_n239_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n243_), .A2(new_n244_), .ZN(new_n558_));
  AOI22_X1  g357(.A1(new_n557_), .A2(new_n558_), .B1(new_n224_), .B2(new_n208_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n547_), .B1(new_n559_), .B2(new_n499_), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n225_), .B(new_n498_), .C1(new_n245_), .C2(new_n246_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n499_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n247_), .A2(KEYINPUT75), .A3(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n560_), .A2(new_n561_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G232gat), .A2(G233gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT34), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n567_), .A2(KEYINPUT35), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n567_), .A2(KEYINPUT35), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n565_), .A2(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(G190gat), .B(G218gat), .Z(new_n572_));
  XNOR2_X1  g371(.A(G134gat), .B(G162gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT77), .B(KEYINPUT36), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT76), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n563_), .A2(new_n561_), .ZN(new_n578_));
  AOI21_X1  g377(.A(KEYINPUT75), .B1(new_n247_), .B2(new_n562_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n577_), .B(new_n568_), .C1(new_n578_), .C2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n577_), .B1(new_n564_), .B2(new_n568_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n571_), .B(new_n576_), .C1(new_n581_), .C2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT78), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n568_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(KEYINPUT76), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(new_n580_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT78), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n587_), .A2(new_n588_), .A3(new_n571_), .A4(new_n576_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n584_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT79), .ZN(new_n591_));
  AOI22_X1  g390(.A1(new_n586_), .A2(new_n580_), .B1(new_n565_), .B2(new_n570_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n574_), .B(KEYINPUT36), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n591_), .B1(new_n592_), .B2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n571_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n596_), .A2(KEYINPUT79), .A3(new_n593_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(KEYINPUT37), .B1(new_n590_), .B2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n584_), .A2(new_n589_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n596_), .A2(new_n593_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(KEYINPUT80), .B(KEYINPUT37), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n600_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n546_), .B1(new_n599_), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n531_), .A2(new_n604_), .ZN(new_n605_));
  OR3_X1    g404(.A1(new_n605_), .A2(G1gat), .A3(new_n489_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT38), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n292_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n600_), .A2(new_n601_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n611_), .A2(new_n546_), .ZN(new_n612_));
  AND3_X1   g411(.A1(new_n529_), .A2(new_n609_), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(G1gat), .B1(new_n614_), .B2(new_n489_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n606_), .A2(new_n607_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n608_), .A2(new_n615_), .A3(new_n616_), .ZN(G1324gat));
  INV_X1    g416(.A(G8gat), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n618_), .B1(new_n613_), .B2(new_n486_), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n619_), .B(KEYINPUT39), .Z(new_n620_));
  INV_X1    g419(.A(new_n605_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT105), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n486_), .A2(new_n618_), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n621_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n622_), .B1(new_n621_), .B2(new_n623_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n620_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT40), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  OAI211_X1 g427(.A(KEYINPUT40), .B(new_n620_), .C1(new_n624_), .C2(new_n625_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(G1325gat));
  OAI21_X1  g429(.A(G15gat), .B1(new_n614_), .B2(new_n484_), .ZN(new_n631_));
  XOR2_X1   g430(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n484_), .A2(G15gat), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n633_), .B1(new_n605_), .B2(new_n634_), .ZN(G1326gat));
  INV_X1    g434(.A(G22gat), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n621_), .A2(new_n636_), .A3(new_n452_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n636_), .B1(new_n613_), .B2(new_n452_), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n638_), .B(KEYINPUT42), .Z(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(G1327gat));
  NOR2_X1   g439(.A1(new_n610_), .A2(new_n545_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n527_), .A2(new_n530_), .A3(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(G29gat), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n642_), .A2(new_n643_), .A3(new_n459_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT44), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n645_), .A2(KEYINPUT107), .ZN(new_n646_));
  NOR4_X1   g445(.A1(new_n292_), .A2(new_n545_), .A3(new_n528_), .A4(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT37), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n592_), .A2(new_n591_), .A3(new_n594_), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT79), .B1(new_n596_), .B2(new_n593_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n648_), .B1(new_n651_), .B2(new_n600_), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n600_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n491_), .A2(new_n654_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n655_), .A2(KEYINPUT43), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(KEYINPUT43), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n647_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n645_), .A2(KEYINPUT107), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n655_), .B(KEYINPUT43), .ZN(new_n661_));
  INV_X1    g460(.A(new_n659_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n661_), .A2(new_n662_), .A3(new_n647_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n489_), .B1(new_n660_), .B2(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n644_), .B1(new_n664_), .B2(new_n643_), .ZN(G1328gat));
  INV_X1    g464(.A(KEYINPUT46), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n666_), .A2(KEYINPUT110), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(KEYINPUT110), .ZN(new_n668_));
  INV_X1    g467(.A(G36gat), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n660_), .A2(new_n663_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n669_), .B1(new_n670_), .B2(new_n486_), .ZN(new_n671_));
  XOR2_X1   g470(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n672_));
  INV_X1    g471(.A(KEYINPUT108), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n486_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n486_), .A2(new_n673_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n676_), .A2(G36gat), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n672_), .B1(new_n642_), .B2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n527_), .A2(new_n530_), .A3(new_n641_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n677_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n672_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n679_), .A2(new_n680_), .A3(new_n681_), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n678_), .A2(new_n682_), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n667_), .B(new_n668_), .C1(new_n671_), .C2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n670_), .A2(new_n486_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(G36gat), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n678_), .A2(new_n682_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n686_), .A2(KEYINPUT110), .A3(new_n666_), .A4(new_n687_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n684_), .A2(new_n688_), .ZN(G1329gat));
  INV_X1    g488(.A(G43gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n690_), .B1(new_n679_), .B2(new_n484_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT112), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n691_), .B(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n484_), .A2(new_n690_), .ZN(new_n694_));
  AOI21_X1  g493(.A(KEYINPUT111), .B1(new_n670_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT111), .ZN(new_n696_));
  INV_X1    g495(.A(new_n694_), .ZN(new_n697_));
  AOI211_X1 g496(.A(new_n696_), .B(new_n697_), .C1(new_n660_), .C2(new_n663_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n693_), .B1(new_n695_), .B2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(KEYINPUT47), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT47), .ZN(new_n701_));
  OAI211_X1 g500(.A(new_n693_), .B(new_n701_), .C1(new_n695_), .C2(new_n698_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(G1330gat));
  OR3_X1    g502(.A1(new_n679_), .A2(G50gat), .A3(new_n451_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n451_), .B1(new_n660_), .B2(new_n663_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n705_), .A2(KEYINPUT113), .ZN(new_n706_));
  OAI21_X1  g505(.A(G50gat), .B1(new_n705_), .B2(KEYINPUT113), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n704_), .B1(new_n706_), .B2(new_n707_), .ZN(G1331gat));
  NOR2_X1   g507(.A1(new_n609_), .A2(new_n524_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n709_), .A2(new_n491_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(new_n612_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n712_), .A2(G57gat), .A3(new_n459_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n710_), .A2(new_n604_), .ZN(new_n714_));
  AOI21_X1  g513(.A(G57gat), .B1(new_n714_), .B2(new_n459_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1332gat));
  INV_X1    g515(.A(G64gat), .ZN(new_n717_));
  INV_X1    g516(.A(new_n676_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n714_), .A2(new_n717_), .A3(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G64gat), .B1(new_n711_), .B2(new_n676_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(KEYINPUT114), .B(KEYINPUT48), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n721_), .A2(new_n722_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n719_), .B1(new_n723_), .B2(new_n724_), .ZN(G1333gat));
  INV_X1    g524(.A(G71gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n714_), .A2(new_n726_), .A3(new_n488_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT49), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n712_), .A2(new_n488_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(G71gat), .ZN(new_n730_));
  AOI211_X1 g529(.A(KEYINPUT49), .B(new_n726_), .C1(new_n712_), .C2(new_n488_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT115), .Z(G1334gat));
  INV_X1    g532(.A(G78gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n714_), .A2(new_n734_), .A3(new_n452_), .ZN(new_n735_));
  OAI21_X1  g534(.A(G78gat), .B1(new_n711_), .B2(new_n451_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n736_), .A2(KEYINPUT50), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n736_), .A2(KEYINPUT50), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n735_), .B1(new_n737_), .B2(new_n738_), .ZN(G1335gat));
  AND2_X1   g538(.A1(new_n710_), .A2(new_n641_), .ZN(new_n740_));
  AOI21_X1  g539(.A(G85gat), .B1(new_n740_), .B2(new_n459_), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n661_), .A2(new_n546_), .A3(new_n709_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n489_), .A2(new_n202_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n741_), .B1(new_n742_), .B2(new_n743_), .ZN(G1336gat));
  AOI21_X1  g543(.A(G92gat), .B1(new_n740_), .B2(new_n486_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n676_), .A2(new_n203_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n742_), .B2(new_n746_), .ZN(G1337gat));
  AOI21_X1  g546(.A(new_n548_), .B1(new_n742_), .B2(new_n488_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n484_), .A2(new_n205_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n740_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n750_), .B(new_n751_), .ZN(G1338gat));
  NAND3_X1  g551(.A1(new_n740_), .A2(new_n549_), .A3(new_n452_), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n661_), .A2(new_n546_), .A3(new_n452_), .A4(new_n709_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT52), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n754_), .A2(new_n755_), .A3(G106gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n754_), .B2(G106gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n753_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g558(.A(KEYINPUT121), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT59), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n264_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT117), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n264_), .A2(KEYINPUT117), .A3(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n259_), .A2(new_n261_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT70), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n259_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n247_), .A2(KEYINPUT12), .A3(new_n254_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT12), .B1(new_n247_), .B2(new_n254_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n770_), .A2(new_n773_), .A3(KEYINPUT55), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n257_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n266_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n765_), .A2(new_n766_), .A3(new_n774_), .A4(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT118), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n777_), .A2(new_n778_), .A3(KEYINPUT56), .A4(new_n276_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n524_), .A2(new_n279_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(KEYINPUT55), .B1(new_n770_), .B2(new_n773_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n774_), .B(new_n776_), .C1(new_n782_), .C2(KEYINPUT117), .ZN(new_n783_));
  INV_X1    g582(.A(new_n766_), .ZN(new_n784_));
  OAI211_X1 g583(.A(KEYINPUT56), .B(new_n276_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT56), .B1(new_n777_), .B2(new_n276_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n781_), .B1(new_n788_), .B2(KEYINPUT118), .ZN(new_n789_));
  INV_X1    g588(.A(new_n516_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n515_), .A2(new_n790_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n791_), .B(new_n495_), .C1(new_n790_), .C2(new_n518_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n792_), .A2(new_n523_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n284_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  OAI211_X1 g594(.A(KEYINPUT57), .B(new_n610_), .C1(new_n789_), .C2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT119), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n777_), .A2(new_n276_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT56), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n801_), .A2(KEYINPUT118), .A3(new_n785_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n781_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n794_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n805_), .A2(KEYINPUT119), .A3(KEYINPUT57), .A4(new_n610_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n795_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n807_), .B1(new_n808_), .B2(new_n611_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n279_), .B(new_n793_), .C1(new_n786_), .C2(new_n787_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT58), .ZN(new_n811_));
  OR2_X1    g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n811_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n812_), .A2(new_n654_), .A3(new_n813_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n798_), .A2(new_n806_), .A3(new_n809_), .A4(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n546_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n545_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n290_), .A2(new_n528_), .A3(new_n291_), .ZN(new_n818_));
  OAI21_X1  g617(.A(KEYINPUT54), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n290_), .A2(new_n528_), .A3(new_n291_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n604_), .A2(new_n820_), .A3(new_n821_), .A4(new_n822_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n819_), .A2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n604_), .A2(new_n822_), .A3(new_n821_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT116), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n489_), .B1(new_n816_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n487_), .A2(new_n488_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n761_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n831_));
  AOI22_X1  g630(.A1(new_n815_), .A2(new_n546_), .B1(new_n826_), .B2(new_n824_), .ZN(new_n832_));
  NOR4_X1   g631(.A1(new_n832_), .A2(KEYINPUT59), .A3(new_n489_), .A4(new_n829_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n524_), .A2(G113gat), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(KEYINPUT120), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NOR3_X1   g635(.A1(new_n831_), .A2(new_n833_), .A3(new_n836_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n832_), .A2(new_n489_), .A3(new_n829_), .ZN(new_n838_));
  AOI21_X1  g637(.A(G113gat), .B1(new_n838_), .B2(new_n524_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n760_), .B1(new_n837_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n828_), .A2(new_n830_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT59), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n838_), .A2(new_n761_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n843_), .A3(new_n835_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n839_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(new_n845_), .A3(KEYINPUT121), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n840_), .A2(new_n846_), .ZN(G1340gat));
  INV_X1    g646(.A(G120gat), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n609_), .B2(KEYINPUT60), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n838_), .B(new_n849_), .C1(KEYINPUT60), .C2(new_n848_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n831_), .A2(new_n833_), .A3(new_n609_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n848_), .ZN(G1341gat));
  AOI21_X1  g651(.A(G127gat), .B1(new_n838_), .B2(new_n545_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n831_), .A2(new_n833_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n545_), .A2(G127gat), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n853_), .B1(new_n854_), .B2(new_n855_), .ZN(G1342gat));
  AOI21_X1  g655(.A(G134gat), .B1(new_n838_), .B2(new_n611_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n654_), .A2(G134gat), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n857_), .B1(new_n854_), .B2(new_n858_), .ZN(G1343gat));
  NOR3_X1   g658(.A1(new_n718_), .A2(new_n488_), .A3(new_n451_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n828_), .A2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n524_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n292_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g664(.A1(new_n828_), .A2(new_n545_), .A3(new_n860_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(KEYINPUT122), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n828_), .A2(new_n868_), .A3(new_n545_), .A4(new_n860_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(KEYINPUT61), .B(G155gat), .ZN(new_n870_));
  AND3_X1   g669(.A1(new_n867_), .A2(new_n869_), .A3(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n870_), .B1(new_n867_), .B2(new_n869_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n871_), .A2(new_n872_), .ZN(G1346gat));
  AOI21_X1  g672(.A(G162gat), .B1(new_n861_), .B2(new_n611_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n654_), .A2(G162gat), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n861_), .B2(new_n875_), .ZN(G1347gat));
  NOR2_X1   g675(.A1(new_n832_), .A2(new_n676_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n452_), .A2(new_n484_), .A3(new_n459_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(G169gat), .B1(new_n879_), .B2(new_n528_), .ZN(new_n880_));
  XOR2_X1   g679(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n879_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n884_), .A2(new_n524_), .A3(new_n321_), .ZN(new_n885_));
  OAI211_X1 g684(.A(G169gat), .B(new_n881_), .C1(new_n879_), .C2(new_n528_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n883_), .A2(new_n885_), .A3(new_n886_), .ZN(G1348gat));
  NOR2_X1   g686(.A1(new_n879_), .A2(new_n609_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(new_n311_), .ZN(G1349gat));
  NOR2_X1   g688(.A1(new_n879_), .A2(new_n546_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n336_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n891_), .B1(new_n297_), .B2(new_n890_), .ZN(G1350gat));
  INV_X1    g691(.A(new_n654_), .ZN(new_n893_));
  OAI21_X1  g692(.A(G190gat), .B1(new_n879_), .B2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n611_), .A2(new_n314_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n879_), .B2(new_n895_), .ZN(G1351gat));
  NAND2_X1  g695(.A1(new_n460_), .A2(new_n484_), .ZN(new_n897_));
  XOR2_X1   g696(.A(new_n897_), .B(KEYINPUT124), .Z(new_n898_));
  NAND2_X1  g697(.A1(new_n877_), .A2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(G197gat), .ZN(new_n900_));
  OAI22_X1  g699(.A1(new_n899_), .A2(new_n528_), .B1(KEYINPUT125), .B2(new_n900_), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n900_), .A2(KEYINPUT125), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1352gat));
  INV_X1    g702(.A(new_n899_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n292_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g705(.A(new_n546_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n904_), .A2(new_n907_), .ZN(new_n908_));
  XOR2_X1   g707(.A(KEYINPUT126), .B(KEYINPUT127), .Z(new_n909_));
  NOR2_X1   g708(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n909_), .B(new_n910_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n908_), .B(new_n911_), .ZN(G1354gat));
  AND3_X1   g711(.A1(new_n904_), .A2(G218gat), .A3(new_n654_), .ZN(new_n913_));
  AOI21_X1  g712(.A(G218gat), .B1(new_n904_), .B2(new_n611_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1355gat));
endmodule


