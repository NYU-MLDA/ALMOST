//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 1 0 1 1 1 1 1 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n797_, new_n798_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n953_, new_n954_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n962_,
    new_n963_, new_n965_, new_n966_, new_n967_, new_n969_, new_n970_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT6), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT7), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n204_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G85gat), .ZN(new_n211_));
  INV_X1    g010(.A(G92gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G85gat), .A2(G92gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NOR3_X1   g014(.A1(new_n210_), .A2(KEYINPUT8), .A3(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n204_), .B1(KEYINPUT66), .B2(new_n209_), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n209_), .A2(KEYINPUT66), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n215_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT8), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n217_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  XOR2_X1   g021(.A(G71gat), .B(G78gat), .Z(new_n223_));
  XNOR2_X1  g022(.A(G57gat), .B(G64gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n223_), .B1(KEYINPUT11), .B2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(KEYINPUT11), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n225_), .B(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT9), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n213_), .B1(new_n229_), .B2(new_n214_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT64), .B(G85gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n229_), .B1(new_n231_), .B2(new_n212_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n230_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n234_), .B1(new_n233_), .B2(new_n232_), .ZN(new_n235_));
  INV_X1    g034(.A(G106gat), .ZN(new_n236_));
  XOR2_X1   g035(.A(KEYINPUT10), .B(G99gat), .Z(new_n237_));
  AOI21_X1  g036(.A(new_n204_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n235_), .A2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n222_), .A2(new_n228_), .A3(new_n239_), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n240_), .A2(KEYINPUT67), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(KEYINPUT67), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT68), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n241_), .A2(new_n245_), .A3(new_n242_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n220_), .A2(new_n221_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n247_), .A2(new_n216_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n239_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n227_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n244_), .A2(new_n246_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G230gat), .A2(G233gat), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n222_), .A2(new_n255_), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n217_), .B(KEYINPUT69), .C1(new_n221_), .C2(new_n220_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(new_n239_), .A3(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT12), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n228_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n250_), .A2(new_n259_), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n240_), .A2(new_n252_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n261_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G120gat), .B(G148gat), .ZN(new_n265_));
  INV_X1    g064(.A(G204gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT5), .B(G176gat), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n267_), .B(new_n268_), .Z(new_n269_));
  NAND3_X1  g068(.A1(new_n254_), .A2(new_n264_), .A3(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n269_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n250_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n272_), .B1(new_n243_), .B2(KEYINPUT68), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n252_), .B1(new_n273_), .B2(new_n246_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n264_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n271_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n270_), .A2(new_n276_), .A3(KEYINPUT70), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(KEYINPUT70), .B1(new_n270_), .B2(new_n276_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT13), .ZN(new_n280_));
  NOR3_X1   g079(.A1(new_n278_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n270_), .A2(new_n276_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(KEYINPUT13), .B1(new_n284_), .B2(new_n277_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n281_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G29gat), .B(G36gat), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(G43gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(G50gat), .ZN(new_n291_));
  INV_X1    g090(.A(G43gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n289_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(G50gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n291_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT15), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n291_), .A2(new_n295_), .A3(KEYINPUT15), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G15gat), .B(G22gat), .ZN(new_n301_));
  INV_X1    g100(.A(G1gat), .ZN(new_n302_));
  INV_X1    g101(.A(G8gat), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT14), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n301_), .A2(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(G1gat), .B(G8gat), .Z(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n300_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G229gat), .A2(G233gat), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n309_), .B(new_n310_), .C1(new_n308_), .C2(new_n296_), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n296_), .B(new_n307_), .Z(new_n312_));
  INV_X1    g111(.A(new_n310_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n311_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G113gat), .B(G141gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(G169gat), .ZN(new_n318_));
  INV_X1    g117(.A(G197gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n316_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n320_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n315_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n286_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G8gat), .B(G36gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT18), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(G64gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(G92gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G226gat), .A2(G233gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT19), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT25), .B(G183gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT26), .B(G190gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G183gat), .A2(G190gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT23), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT23), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n339_), .A2(G183gat), .A3(G190gat), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT24), .ZN(new_n341_));
  NOR2_X1   g140(.A1(G169gat), .A2(G176gat), .ZN(new_n342_));
  AOI22_X1  g141(.A1(new_n338_), .A2(new_n340_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n336_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G169gat), .A2(G176gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT76), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT76), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n347_), .A2(G169gat), .A3(G176gat), .ZN(new_n348_));
  INV_X1    g147(.A(new_n342_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n346_), .A2(new_n348_), .A3(new_n349_), .A4(KEYINPUT24), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n346_), .A2(new_n348_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT22), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n352_), .A2(G169gat), .ZN(new_n353_));
  INV_X1    g152(.A(G169gat), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n354_), .A2(KEYINPUT22), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT77), .B1(new_n353_), .B2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(KEYINPUT22), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT77), .ZN(new_n358_));
  AOI21_X1  g157(.A(G176gat), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n351_), .B1(new_n356_), .B2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n338_), .A2(new_n340_), .A3(KEYINPUT78), .ZN(new_n361_));
  OR3_X1    g160(.A1(new_n337_), .A2(KEYINPUT78), .A3(KEYINPUT23), .ZN(new_n362_));
  OR2_X1    g161(.A1(G183gat), .A2(G190gat), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n361_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  AOI22_X1  g163(.A1(new_n344_), .A2(new_n350_), .B1(new_n360_), .B2(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(G197gat), .A2(G204gat), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G197gat), .A2(G204gat), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n367_), .A2(KEYINPUT21), .A3(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT21), .ZN(new_n370_));
  INV_X1    g169(.A(new_n368_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n370_), .B1(new_n371_), .B2(new_n366_), .ZN(new_n372_));
  INV_X1    g171(.A(G218gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(G211gat), .ZN(new_n374_));
  INV_X1    g173(.A(G211gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(G218gat), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT85), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n374_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n377_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n369_), .B(new_n372_), .C1(new_n378_), .C2(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n375_), .A2(G218gat), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n373_), .A2(G211gat), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT85), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NOR3_X1   g182(.A1(new_n371_), .A2(new_n366_), .A3(new_n370_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n374_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n383_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n380_), .A2(KEYINPUT86), .A3(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(KEYINPUT86), .B1(new_n380_), .B2(new_n386_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n365_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT20), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n338_), .A2(new_n340_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n363_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT22), .B(G169gat), .ZN(new_n393_));
  INV_X1    g192(.A(G176gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT90), .ZN(new_n396_));
  AND3_X1   g195(.A1(new_n346_), .A2(new_n348_), .A3(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n396_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n392_), .B(new_n395_), .C1(new_n397_), .C2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT91), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  AND2_X1   g200(.A1(new_n361_), .A2(new_n362_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n341_), .A2(KEYINPUT89), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n341_), .A2(KEYINPUT89), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n345_), .B(new_n349_), .C1(new_n403_), .C2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n342_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n402_), .A2(new_n336_), .A3(new_n405_), .A4(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n351_), .A2(KEYINPUT90), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n346_), .A2(new_n348_), .A3(new_n396_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  AOI22_X1  g210(.A1(new_n391_), .A2(new_n363_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(new_n412_), .A3(KEYINPUT91), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n401_), .A2(new_n408_), .A3(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n378_), .A2(new_n379_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n369_), .A2(new_n372_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n386_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(KEYINPUT92), .B1(new_n414_), .B2(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n390_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n414_), .A2(KEYINPUT92), .A3(new_n417_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n333_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT86), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n417_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n360_), .A2(new_n364_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n350_), .A2(new_n336_), .A3(new_n343_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n380_), .A2(KEYINPUT86), .A3(new_n386_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n423_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n417_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n429_), .A2(new_n401_), .A3(new_n413_), .A4(new_n408_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT20), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n332_), .A2(new_n431_), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n428_), .A2(new_n430_), .A3(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n330_), .B1(new_n421_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n414_), .A2(new_n417_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT92), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n423_), .A2(new_n427_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n431_), .B1(new_n438_), .B2(new_n365_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n437_), .A2(new_n439_), .A3(new_n420_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n433_), .B1(new_n440_), .B2(new_n332_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n330_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n434_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT27), .ZN(new_n445_));
  INV_X1    g244(.A(new_n428_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n405_), .A2(new_n336_), .A3(new_n407_), .ZN(new_n447_));
  AOI22_X1  g246(.A1(new_n447_), .A2(new_n402_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT87), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n417_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n380_), .A2(KEYINPUT87), .A3(new_n386_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n448_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT20), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n446_), .B1(new_n453_), .B2(KEYINPUT95), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT95), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n452_), .A2(new_n455_), .A3(KEYINPUT20), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n333_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n440_), .A2(new_n332_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n330_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n445_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n460_));
  AOI22_X1  g259(.A1(new_n444_), .A2(new_n445_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G1gat), .B(G29gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT0), .ZN(new_n463_));
  INV_X1    g262(.A(G57gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(new_n211_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G225gat), .A2(G233gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G127gat), .B(G134gat), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(G113gat), .B(G120gat), .Z(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT81), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G113gat), .B(G120gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n469_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n472_), .A2(new_n473_), .A3(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n470_), .A2(new_n471_), .A3(KEYINPUT81), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  AND2_X1   g277(.A1(G155gat), .A2(G162gat), .ZN(new_n479_));
  NOR2_X1   g278(.A1(G155gat), .A2(G162gat), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G141gat), .A2(G148gat), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT82), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(KEYINPUT82), .A2(G141gat), .A3(G148gat), .ZN(new_n486_));
  OR2_X1    g285(.A1(KEYINPUT83), .A2(KEYINPUT2), .ZN(new_n487_));
  NAND2_X1  g286(.A1(KEYINPUT83), .A2(KEYINPUT2), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n485_), .A2(new_n486_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT3), .ZN(new_n490_));
  INV_X1    g289(.A(G141gat), .ZN(new_n491_));
  INV_X1    g290(.A(G148gat), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT2), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n493_), .B(new_n494_), .C1(new_n495_), .C2(new_n483_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n482_), .B1(new_n489_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n485_), .A2(new_n486_), .ZN(new_n498_));
  AOI22_X1  g297(.A1(new_n479_), .A2(KEYINPUT1), .B1(new_n491_), .B2(new_n492_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n498_), .B(new_n499_), .C1(new_n481_), .C2(KEYINPUT1), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(KEYINPUT4), .B1(new_n478_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n478_), .A2(new_n501_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n472_), .A2(new_n475_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n503_), .B1(new_n504_), .B2(new_n501_), .ZN(new_n505_));
  AOI211_X1 g304(.A(new_n468_), .B(new_n502_), .C1(new_n505_), .C2(KEYINPUT4), .ZN(new_n506_));
  INV_X1    g305(.A(new_n468_), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n501_), .A2(new_n504_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n507_), .B1(new_n508_), .B2(new_n503_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n467_), .B1(new_n506_), .B2(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n502_), .B1(new_n505_), .B2(KEYINPUT4), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(new_n507_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n509_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(new_n466_), .A3(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n510_), .A2(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n426_), .A2(KEYINPUT79), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT79), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n517_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT30), .ZN(new_n519_));
  NOR3_X1   g318(.A1(new_n516_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n518_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n365_), .A2(new_n517_), .ZN(new_n522_));
  AOI21_X1  g321(.A(KEYINPUT30), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT80), .B1(new_n520_), .B2(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n519_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n521_), .A2(new_n522_), .A3(KEYINPUT30), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT80), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n525_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(G15gat), .B(G43gat), .Z(new_n529_));
  NAND2_X1  g328(.A1(G227gat), .A2(G233gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G71gat), .B(G99gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n524_), .A2(new_n528_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n533_), .ZN(new_n535_));
  OAI211_X1 g334(.A(KEYINPUT80), .B(new_n535_), .C1(new_n520_), .C2(new_n523_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(new_n478_), .B(KEYINPUT31), .Z(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n534_), .A2(new_n538_), .A3(new_n536_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n515_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(G22gat), .B(G50gat), .Z(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT28), .ZN(new_n544_));
  INV_X1    g343(.A(new_n501_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT29), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n544_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  AND4_X1   g346(.A1(new_n546_), .A2(new_n544_), .A3(new_n497_), .A4(new_n500_), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n501_), .A2(KEYINPUT29), .ZN(new_n550_));
  INV_X1    g349(.A(G233gat), .ZN(new_n551_));
  NOR2_X1   g350(.A1(KEYINPUT84), .A2(G228gat), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(KEYINPUT84), .A2(G228gat), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n551_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n550_), .A2(new_n423_), .A3(new_n556_), .A4(new_n427_), .ZN(new_n557_));
  AOI22_X1  g356(.A1(new_n450_), .A2(new_n451_), .B1(KEYINPUT29), .B2(new_n501_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n557_), .B1(new_n558_), .B2(new_n556_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n549_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(KEYINPUT88), .B1(new_n549_), .B2(new_n559_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G78gat), .B(G106gat), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  AOI211_X1 g364(.A(KEYINPUT88), .B(new_n563_), .C1(new_n549_), .C2(new_n559_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n561_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n547_), .A2(new_n548_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n450_), .A2(new_n451_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(new_n550_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(new_n555_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n568_), .B1(new_n571_), .B2(new_n557_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n563_), .B1(new_n572_), .B2(KEYINPUT88), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n562_), .A2(new_n564_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n573_), .A2(new_n574_), .A3(new_n560_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n567_), .A2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n461_), .A2(new_n542_), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT98), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n461_), .A2(new_n542_), .A3(KEYINPUT98), .A4(new_n576_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n440_), .A2(new_n332_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n433_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n442_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  AOI211_X1 g383(.A(new_n330_), .B(new_n433_), .C1(new_n440_), .C2(new_n332_), .ZN(new_n585_));
  OAI21_X1  g384(.A(KEYINPUT93), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT93), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n434_), .A2(new_n443_), .A3(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n466_), .B1(new_n468_), .B2(new_n505_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n511_), .A2(new_n507_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n509_), .B1(new_n511_), .B2(new_n507_), .ZN(new_n592_));
  OAI22_X1  g391(.A1(new_n592_), .A2(new_n466_), .B1(KEYINPUT94), .B2(KEYINPUT33), .ZN(new_n593_));
  NOR2_X1   g392(.A1(KEYINPUT94), .A2(KEYINPUT33), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n467_), .B(new_n594_), .C1(new_n506_), .C2(new_n509_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n591_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n586_), .A2(new_n588_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT32), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n330_), .A2(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n599_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n441_), .B1(new_n598_), .B2(new_n330_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n600_), .A2(new_n601_), .A3(new_n515_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT96), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n600_), .A2(new_n601_), .A3(new_n515_), .A4(KEYINPUT96), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n597_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(new_n576_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n459_), .A2(new_n460_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n445_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n515_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n567_), .A2(new_n611_), .A3(new_n575_), .ZN(new_n612_));
  OAI21_X1  g411(.A(KEYINPUT97), .B1(new_n610_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n612_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT97), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n614_), .A2(new_n461_), .A3(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n607_), .A2(new_n613_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n540_), .A2(new_n541_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n581_), .B1(new_n617_), .B2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n300_), .A2(new_n258_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n296_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n248_), .A2(new_n249_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G232gat), .A2(G233gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT34), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT35), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT72), .B1(new_n626_), .B2(KEYINPUT35), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n621_), .A2(new_n624_), .A3(new_n630_), .A4(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n624_), .A2(new_n632_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n249_), .B1(new_n222_), .B2(new_n255_), .ZN(new_n635_));
  AOI22_X1  g434(.A1(new_n298_), .A2(new_n299_), .B1(new_n635_), .B2(new_n257_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n629_), .B1(new_n634_), .B2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n633_), .A2(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G190gat), .B(G218gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(G134gat), .B(G162gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT36), .Z(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT74), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n638_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT75), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n638_), .A2(KEYINPUT75), .A3(new_n643_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n641_), .A2(KEYINPUT36), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n633_), .A2(new_n637_), .A3(new_n648_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n649_), .A2(KEYINPUT73), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(KEYINPUT73), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n646_), .B(new_n647_), .C1(new_n650_), .C2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT37), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n649_), .B(KEYINPUT73), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n653_), .B1(new_n638_), .B2(new_n643_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n654_), .A2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(G127gat), .B(G155gat), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT16), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(G183gat), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(new_n375_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT17), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n662_), .A2(new_n663_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(G231gat), .A2(G233gat), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n307_), .B(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(new_n228_), .ZN(new_n668_));
  OR3_X1    g467(.A1(new_n664_), .A2(new_n665_), .A3(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n665_), .A2(new_n668_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n620_), .A2(new_n658_), .A3(new_n671_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n326_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n674_), .A2(G1gat), .A3(new_n611_), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n675_), .A2(KEYINPUT38), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(KEYINPUT38), .ZN(new_n677_));
  INV_X1    g476(.A(new_n671_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n652_), .A2(KEYINPUT99), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT99), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n655_), .A2(new_n680_), .A3(new_n646_), .A4(new_n647_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n683_), .A2(new_n620_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n326_), .A2(new_n678_), .A3(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G1gat), .B1(new_n685_), .B2(new_n611_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n676_), .A2(new_n677_), .A3(new_n686_), .ZN(G1324gat));
  NAND3_X1  g486(.A1(new_n673_), .A2(new_n303_), .A3(new_n610_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n326_), .A2(new_n684_), .A3(new_n610_), .A4(new_n678_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT39), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n689_), .A2(new_n690_), .A3(G8gat), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n690_), .B1(new_n689_), .B2(G8gat), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n688_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n694_), .A2(KEYINPUT100), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(KEYINPUT100), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n695_), .A2(KEYINPUT40), .A3(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT40), .B1(new_n695_), .B2(new_n696_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n697_), .A2(new_n698_), .ZN(G1325gat));
  OAI21_X1  g498(.A(G15gat), .B1(new_n685_), .B2(new_n619_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT41), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n674_), .A2(G15gat), .A3(new_n619_), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1326gat));
  XNOR2_X1  g502(.A(new_n576_), .B(KEYINPUT101), .ZN(new_n704_));
  OAI21_X1  g503(.A(G22gat), .B1(new_n685_), .B2(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT42), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n704_), .A2(G22gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n706_), .B1(new_n674_), .B2(new_n707_), .ZN(G1327gat));
  OAI211_X1 g507(.A(new_n324_), .B(new_n671_), .C1(new_n281_), .C2(new_n285_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n620_), .A2(new_n682_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  OR3_X1    g511(.A1(new_n712_), .A2(G29gat), .A3(new_n611_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(KEYINPUT102), .B(KEYINPUT43), .ZN(new_n714_));
  AOI22_X1  g513(.A1(new_n652_), .A2(new_n653_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n714_), .B1(new_n620_), .B2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n616_), .A2(new_n613_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n618_), .B1(new_n718_), .B2(new_n607_), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n658_), .B(new_n717_), .C1(new_n719_), .C2(new_n581_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n709_), .B1(new_n716_), .B2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT44), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n723_), .B1(new_n721_), .B2(KEYINPUT103), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT103), .ZN(new_n725_));
  AOI211_X1 g524(.A(new_n725_), .B(new_n709_), .C1(new_n716_), .C2(new_n720_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n515_), .B(new_n722_), .C1(new_n724_), .C2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT104), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n727_), .A2(new_n728_), .A3(G29gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n727_), .B2(G29gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n713_), .B1(new_n729_), .B2(new_n730_), .ZN(G1328gat));
  NOR2_X1   g530(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT108), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n461_), .B1(new_n721_), .B2(KEYINPUT44), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n734_), .B1(new_n724_), .B2(new_n726_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT105), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT105), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n737_), .B(new_n734_), .C1(new_n724_), .C2(new_n726_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n736_), .A2(G36gat), .A3(new_n738_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n461_), .A2(G36gat), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(KEYINPUT106), .B1(new_n712_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT106), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n710_), .A2(new_n743_), .A3(new_n711_), .A4(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT45), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n739_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n733_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n748_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n733_), .ZN(new_n751_));
  AOI211_X1 g550(.A(new_n750_), .B(new_n751_), .C1(new_n739_), .C2(new_n746_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n749_), .A2(new_n752_), .ZN(G1329gat));
  OAI21_X1  g552(.A(new_n292_), .B1(new_n712_), .B2(new_n619_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n722_), .B1(new_n724_), .B2(new_n726_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n618_), .A2(G43gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n754_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g557(.A(G50gat), .B1(new_n755_), .B2(new_n576_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n704_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n294_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT109), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n759_), .B1(new_n712_), .B2(new_n762_), .ZN(G1331gat));
  NAND4_X1  g562(.A1(new_n684_), .A2(new_n325_), .A3(new_n286_), .A4(new_n678_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(KEYINPUT110), .B(G57gat), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n764_), .A2(new_n611_), .A3(new_n765_), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT111), .Z(new_n767_));
  AND3_X1   g566(.A1(new_n672_), .A2(new_n325_), .A3(new_n286_), .ZN(new_n768_));
  AOI21_X1  g567(.A(G57gat), .B1(new_n768_), .B2(new_n515_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1332gat));
  OAI21_X1  g569(.A(G64gat), .B1(new_n764_), .B2(new_n461_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT48), .ZN(new_n772_));
  INV_X1    g571(.A(G64gat), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n768_), .A2(new_n773_), .A3(new_n610_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(G1333gat));
  OAI21_X1  g574(.A(G71gat), .B1(new_n764_), .B2(new_n619_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT49), .ZN(new_n777_));
  INV_X1    g576(.A(G71gat), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n768_), .A2(new_n778_), .A3(new_n618_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(G1334gat));
  OAI21_X1  g579(.A(G78gat), .B1(new_n764_), .B2(new_n704_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n781_), .B(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(G78gat), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n768_), .A2(new_n784_), .A3(new_n760_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(G1335gat));
  NAND2_X1  g585(.A1(new_n716_), .A2(new_n720_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n280_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n284_), .A2(KEYINPUT13), .A3(new_n277_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NOR3_X1   g589(.A1(new_n790_), .A2(new_n324_), .A3(new_n678_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n787_), .A2(new_n791_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n792_), .A2(new_n231_), .A3(new_n611_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n791_), .A2(new_n711_), .ZN(new_n794_));
  AOI21_X1  g593(.A(G85gat), .B1(new_n794_), .B2(new_n515_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n793_), .A2(new_n795_), .ZN(G1336gat));
  OAI21_X1  g595(.A(G92gat), .B1(new_n792_), .B2(new_n461_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n794_), .A2(new_n212_), .A3(new_n610_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(G1337gat));
  INV_X1    g598(.A(KEYINPUT113), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n800_), .A2(KEYINPUT51), .ZN(new_n801_));
  OAI21_X1  g600(.A(G99gat), .B1(new_n792_), .B2(new_n619_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n794_), .A2(new_n237_), .A3(new_n618_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n801_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n800_), .A2(KEYINPUT51), .ZN(new_n805_));
  XOR2_X1   g604(.A(new_n804_), .B(new_n805_), .Z(G1338gat));
  INV_X1    g605(.A(new_n576_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n794_), .A2(new_n236_), .A3(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n787_), .A2(new_n807_), .A3(new_n791_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n809_), .A2(new_n810_), .A3(G106gat), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n810_), .B1(new_n809_), .B2(G106gat), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n808_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g613(.A(KEYINPUT121), .ZN(new_n815_));
  XOR2_X1   g614(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n324_), .B1(new_n818_), .B2(new_n817_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n715_), .A2(new_n820_), .A3(new_n678_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n819_), .B1(new_n286_), .B2(new_n821_), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n654_), .A2(new_n678_), .A3(new_n657_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n819_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n823_), .A2(new_n790_), .A3(new_n824_), .A4(new_n820_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n822_), .A2(new_n825_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n274_), .A2(new_n275_), .A3(new_n271_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n261_), .A2(new_n262_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(new_n243_), .ZN(new_n830_));
  AOI22_X1  g629(.A1(new_n258_), .A2(new_n260_), .B1(new_n250_), .B2(new_n259_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n831_), .A2(KEYINPUT117), .A3(new_n242_), .A4(new_n241_), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n830_), .A2(new_n832_), .A3(new_n253_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n264_), .A2(KEYINPUT116), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(KEYINPUT55), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n264_), .A2(KEYINPUT116), .A3(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n271_), .B1(new_n833_), .B2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n827_), .B1(new_n839_), .B2(KEYINPUT56), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT56), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n841_), .B(new_n271_), .C1(new_n833_), .C2(new_n838_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n840_), .A2(new_n324_), .A3(new_n842_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n309_), .B(new_n313_), .C1(new_n308_), .C2(new_n296_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n320_), .B1(new_n312_), .B2(new_n310_), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n316_), .A2(new_n320_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n284_), .A2(new_n277_), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n843_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n682_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT57), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  AOI22_X1  g650(.A1(new_n843_), .A2(new_n847_), .B1(new_n681_), .B2(new_n679_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT57), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n840_), .A2(new_n846_), .A3(new_n842_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n840_), .A2(KEYINPUT58), .A3(new_n846_), .A4(new_n842_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n856_), .A2(new_n658_), .A3(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n851_), .A2(new_n853_), .A3(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n826_), .B1(new_n859_), .B2(new_n671_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n461_), .A2(new_n618_), .A3(new_n576_), .A4(new_n515_), .ZN(new_n861_));
  OR2_X1    g660(.A1(new_n861_), .A2(KEYINPUT119), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(KEYINPUT119), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n862_), .A2(new_n863_), .A3(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n860_), .A2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n324_), .A2(G113gat), .ZN(new_n867_));
  XOR2_X1   g666(.A(new_n867_), .B(KEYINPUT120), .Z(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n858_), .B1(KEYINPUT57), .B2(new_n852_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n849_), .A2(new_n850_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n671_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n826_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n861_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(KEYINPUT118), .B1(new_n874_), .B2(new_n863_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n876_), .B(KEYINPUT59), .C1(new_n860_), .C2(new_n861_), .ZN(new_n877_));
  AOI211_X1 g676(.A(new_n866_), .B(new_n869_), .C1(new_n875_), .C2(new_n877_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n860_), .A2(new_n325_), .A3(new_n861_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(G113gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n815_), .B1(new_n878_), .B2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n875_), .A2(new_n877_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n866_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n882_), .A2(new_n883_), .A3(new_n868_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n880_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n884_), .A2(KEYINPUT121), .A3(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n881_), .A2(new_n886_), .ZN(G1340gat));
  INV_X1    g686(.A(G120gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n888_), .B1(new_n790_), .B2(KEYINPUT60), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n874_), .B(new_n889_), .C1(KEYINPUT60), .C2(new_n888_), .ZN(new_n890_));
  AOI211_X1 g689(.A(new_n790_), .B(new_n866_), .C1(new_n875_), .C2(new_n877_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n891_), .B2(new_n888_), .ZN(G1341gat));
  INV_X1    g691(.A(G127gat), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n874_), .A2(new_n893_), .A3(new_n678_), .ZN(new_n894_));
  AOI211_X1 g693(.A(new_n671_), .B(new_n866_), .C1(new_n875_), .C2(new_n877_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(new_n893_), .ZN(G1342gat));
  INV_X1    g695(.A(G134gat), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n874_), .A2(new_n897_), .A3(new_n683_), .ZN(new_n898_));
  AOI211_X1 g697(.A(new_n715_), .B(new_n866_), .C1(new_n875_), .C2(new_n877_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(new_n897_), .ZN(G1343gat));
  NOR2_X1   g699(.A1(new_n618_), .A2(new_n576_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n860_), .A2(new_n902_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n610_), .A2(new_n611_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n903_), .A2(KEYINPUT122), .A3(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  AOI21_X1  g705(.A(KEYINPUT122), .B1(new_n903_), .B2(new_n904_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n324_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(G141gat), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n903_), .A2(new_n904_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n905_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n913_), .A2(new_n491_), .A3(new_n324_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n909_), .A2(new_n914_), .ZN(G1344gat));
  OAI21_X1  g714(.A(new_n286_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(G148gat), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n913_), .A2(new_n492_), .A3(new_n286_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1345gat));
  XNOR2_X1  g718(.A(KEYINPUT61), .B(G155gat), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(KEYINPUT123), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n921_), .B1(new_n913_), .B2(new_n678_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n921_), .ZN(new_n923_));
  AOI211_X1 g722(.A(new_n671_), .B(new_n923_), .C1(new_n912_), .C2(new_n905_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n922_), .A2(new_n924_), .ZN(G1346gat));
  INV_X1    g724(.A(G162gat), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n913_), .A2(new_n926_), .A3(new_n683_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n715_), .B1(new_n912_), .B2(new_n905_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n927_), .B1(new_n926_), .B2(new_n928_), .ZN(G1347gat));
  NOR2_X1   g728(.A1(new_n461_), .A2(new_n515_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(new_n618_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n860_), .A2(new_n760_), .A3(new_n931_), .ZN(new_n932_));
  INV_X1    g731(.A(new_n932_), .ZN(new_n933_));
  OAI21_X1  g732(.A(G169gat), .B1(new_n933_), .B2(new_n325_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT62), .ZN(new_n935_));
  OR2_X1    g734(.A1(new_n934_), .A2(new_n935_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n932_), .A2(new_n324_), .A3(new_n393_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n934_), .A2(new_n935_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n936_), .A2(new_n937_), .A3(new_n938_), .ZN(G1348gat));
  AOI21_X1  g738(.A(G176gat), .B1(new_n932_), .B2(new_n286_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n872_), .A2(new_n873_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(new_n576_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(KEYINPUT124), .ZN(new_n943_));
  NOR3_X1   g742(.A1(new_n790_), .A2(new_n394_), .A3(new_n931_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n940_), .B1(new_n943_), .B2(new_n944_), .ZN(G1349gat));
  NOR2_X1   g744(.A1(new_n671_), .A2(new_n334_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n932_), .A2(new_n946_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT125), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n947_), .B(new_n948_), .ZN(new_n949_));
  NAND4_X1  g748(.A1(new_n943_), .A2(new_n618_), .A3(new_n678_), .A4(new_n930_), .ZN(new_n950_));
  INV_X1    g749(.A(G183gat), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n949_), .B1(new_n950_), .B2(new_n951_), .ZN(G1350gat));
  OAI21_X1  g751(.A(G190gat), .B1(new_n933_), .B2(new_n715_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n932_), .A2(new_n335_), .A3(new_n683_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n953_), .A2(new_n954_), .ZN(G1351gat));
  NAND3_X1  g754(.A1(new_n903_), .A2(new_n324_), .A3(new_n930_), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n956_), .A2(KEYINPUT126), .A3(new_n319_), .ZN(new_n957_));
  INV_X1    g756(.A(new_n957_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n956_), .A2(new_n319_), .ZN(new_n959_));
  AOI21_X1  g758(.A(KEYINPUT126), .B1(new_n956_), .B2(new_n319_), .ZN(new_n960_));
  NOR3_X1   g759(.A1(new_n958_), .A2(new_n959_), .A3(new_n960_), .ZN(G1352gat));
  NAND2_X1  g760(.A1(new_n903_), .A2(new_n930_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n962_), .A2(new_n790_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(new_n963_), .B(new_n266_), .ZN(G1353gat));
  NOR2_X1   g763(.A1(new_n962_), .A2(new_n671_), .ZN(new_n965_));
  NOR3_X1   g764(.A1(new_n965_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n966_));
  XOR2_X1   g765(.A(KEYINPUT63), .B(G211gat), .Z(new_n967_));
  AOI21_X1  g766(.A(new_n966_), .B1(new_n965_), .B2(new_n967_), .ZN(G1354gat));
  OAI21_X1  g767(.A(G218gat), .B1(new_n962_), .B2(new_n715_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n683_), .A2(new_n373_), .ZN(new_n970_));
  OAI21_X1  g769(.A(new_n969_), .B1(new_n962_), .B2(new_n970_), .ZN(G1355gat));
endmodule


