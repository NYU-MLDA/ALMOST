//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 0 1 1 0 0 0 0 1 1 1 0 1 0 0 1 0 0 0 0 1 1 0 1 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n859_, new_n861_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n912_;
  INV_X1    g000(.A(G50gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(G29gat), .A2(G36gat), .ZN(new_n203_));
  INV_X1    g002(.A(G43gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G29gat), .A2(G36gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n204_), .B1(new_n203_), .B2(new_n205_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n202_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n208_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(G50gat), .A3(new_n206_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G15gat), .B(G22gat), .ZN(new_n213_));
  INV_X1    g012(.A(G1gat), .ZN(new_n214_));
  INV_X1    g013(.A(G8gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT14), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G1gat), .B(G8gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n212_), .B(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G229gat), .A2(G233gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(KEYINPUT76), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n212_), .A2(new_n219_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT15), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n212_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n209_), .A2(new_n211_), .A3(KEYINPUT15), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n225_), .B1(new_n229_), .B2(new_n219_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(KEYINPUT77), .A3(new_n221_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n221_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT77), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n224_), .A2(new_n231_), .A3(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G113gat), .B(G141gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT78), .ZN(new_n237_));
  INV_X1    g036(.A(G169gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G197gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n235_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n241_), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n224_), .A2(new_n231_), .A3(new_n234_), .A4(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT93), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G1gat), .B(G29gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(G85gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT0), .ZN(new_n249_));
  INV_X1    g048(.A(G57gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G225gat), .A2(G233gat), .ZN(new_n252_));
  INV_X1    g051(.A(G141gat), .ZN(new_n253_));
  INV_X1    g052(.A(G148gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(KEYINPUT3), .B1(new_n255_), .B2(KEYINPUT83), .ZN(new_n256_));
  NAND3_X1  g055(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT83), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT3), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n258_), .A2(new_n259_), .A3(new_n253_), .A4(new_n254_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G141gat), .A2(G148gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT2), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n256_), .A2(new_n257_), .A3(new_n260_), .A4(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT84), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G155gat), .A2(G162gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n265_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n268_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n270_), .A2(KEYINPUT84), .A3(new_n266_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n264_), .A2(new_n269_), .A3(new_n271_), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n266_), .A2(KEYINPUT1), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n266_), .A2(KEYINPUT1), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(new_n270_), .A3(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n275_), .A2(new_n261_), .A3(new_n255_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n272_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(G120gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G127gat), .B(G134gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(G113gat), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n279_), .A2(G113gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n278_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n279_), .A2(G113gat), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n284_), .A2(G120gat), .A3(new_n280_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n277_), .A2(new_n286_), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n272_), .A2(new_n283_), .A3(new_n276_), .A4(new_n285_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n287_), .A2(KEYINPUT4), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT4), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n277_), .A2(new_n286_), .A3(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n252_), .B1(new_n289_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n252_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n293_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n251_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT33), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n246_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n289_), .A2(new_n291_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(new_n293_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n294_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n301_), .A2(KEYINPUT93), .A3(KEYINPUT33), .A4(new_n251_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G8gat), .B(G36gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT18), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(G64gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(G92gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G226gat), .A2(G233gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT19), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT20), .ZN(new_n311_));
  OR2_X1    g110(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT91), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT91), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n312_), .A2(new_n316_), .A3(new_n313_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT26), .B(G190gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G169gat), .A2(G176gat), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT24), .ZN(new_n321_));
  INV_X1    g120(.A(G176gat), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n238_), .A2(new_n322_), .A3(KEYINPUT80), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT80), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n324_), .B1(G169gat), .B2(G176gat), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n321_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  AOI22_X1  g125(.A1(new_n318_), .A2(new_n319_), .B1(new_n320_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G183gat), .A2(G190gat), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n328_), .A2(KEYINPUT82), .A3(KEYINPUT23), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT23), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n330_), .A2(G183gat), .A3(G190gat), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(KEYINPUT82), .B1(new_n328_), .B2(KEYINPUT23), .ZN(new_n333_));
  NOR3_X1   g132(.A1(new_n329_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  NOR3_X1   g133(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n328_), .A2(KEYINPUT23), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT81), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n328_), .A2(KEYINPUT81), .A3(KEYINPUT23), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(new_n331_), .A3(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n341_), .B1(G183gat), .B2(G190gat), .ZN(new_n342_));
  NOR2_X1   g141(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(G169gat), .ZN(new_n344_));
  AOI22_X1  g143(.A1(new_n327_), .A2(new_n336_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G197gat), .B(G204gat), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT88), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT21), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n346_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G211gat), .B(G218gat), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n346_), .A2(new_n348_), .ZN(new_n352_));
  INV_X1    g151(.A(G204gat), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n347_), .B1(new_n353_), .B2(G197gat), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n351_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT89), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n350_), .B(new_n356_), .ZN(new_n357_));
  AOI22_X1  g156(.A1(new_n349_), .A2(new_n355_), .B1(new_n357_), .B2(new_n352_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n311_), .B1(new_n345_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n352_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n352_), .A2(new_n354_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n361_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(G183gat), .A2(G190gat), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n344_), .B1(new_n334_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n326_), .A2(new_n320_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT79), .ZN(new_n367_));
  INV_X1    g166(.A(G190gat), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT26), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n368_), .A2(KEYINPUT26), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n314_), .B(new_n369_), .C1(new_n367_), .C2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n323_), .A2(new_n325_), .A3(new_n321_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n366_), .A2(new_n371_), .A3(new_n372_), .A4(new_n341_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n365_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n363_), .A2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n310_), .B1(new_n359_), .B2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT20), .B1(new_n363_), .B2(new_n374_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n318_), .A2(new_n319_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n336_), .A2(new_n378_), .A3(new_n366_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n342_), .A2(new_n344_), .ZN(new_n380_));
  AOI22_X1  g179(.A1(new_n379_), .A2(new_n380_), .B1(new_n362_), .B2(new_n360_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n310_), .ZN(new_n382_));
  NOR3_X1   g181(.A1(new_n377_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n308_), .B1(new_n376_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n379_), .A2(new_n380_), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n375_), .B(KEYINPUT20), .C1(new_n385_), .C2(new_n363_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(new_n382_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n377_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n381_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(new_n389_), .A3(new_n310_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n387_), .A2(new_n390_), .A3(new_n307_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT92), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n384_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n387_), .A2(new_n390_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n394_), .A2(KEYINPUT92), .A3(new_n308_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT94), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n295_), .A2(new_n397_), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n296_), .A2(KEYINPUT95), .ZN(new_n399_));
  OAI211_X1 g198(.A(KEYINPUT94), .B(new_n251_), .C1(new_n292_), .C2(new_n294_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n296_), .A2(KEYINPUT95), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n398_), .A2(new_n399_), .A3(new_n400_), .A4(new_n401_), .ZN(new_n402_));
  OR3_X1    g201(.A1(new_n298_), .A2(KEYINPUT97), .A3(new_n293_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n251_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n287_), .A2(new_n288_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT96), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n287_), .A2(KEYINPUT96), .A3(new_n288_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n293_), .A3(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT97), .B1(new_n298_), .B2(new_n293_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n403_), .A2(new_n404_), .A3(new_n409_), .A4(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n303_), .A2(new_n396_), .A3(new_n402_), .A4(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n301_), .B(new_n251_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT98), .ZN(new_n414_));
  AOI22_X1  g213(.A1(new_n394_), .A2(new_n414_), .B1(KEYINPUT32), .B2(new_n308_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n414_), .B1(new_n387_), .B2(new_n390_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n386_), .A2(new_n310_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n388_), .A2(new_n389_), .A3(new_n382_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n308_), .A2(KEYINPUT32), .ZN(new_n420_));
  NOR3_X1   g219(.A1(new_n416_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n413_), .B1(new_n415_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n412_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(G228gat), .ZN(new_n424_));
  OR2_X1    g223(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n424_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n358_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n277_), .A2(KEYINPUT29), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(KEYINPUT90), .B(KEYINPUT29), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n431_), .B1(new_n272_), .B2(new_n276_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n427_), .B1(new_n432_), .B2(new_n358_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n430_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n277_), .A2(KEYINPUT29), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT85), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT85), .B1(new_n277_), .B2(KEYINPUT29), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G22gat), .B(G50gat), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n438_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n440_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n435_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n438_), .A2(new_n439_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n440_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n438_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n446_), .A2(new_n447_), .A3(new_n434_), .ZN(new_n448_));
  XOR2_X1   g247(.A(G78gat), .B(G106gat), .Z(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(KEYINPUT86), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT28), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n443_), .A2(new_n448_), .A3(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n451_), .B1(new_n443_), .B2(new_n448_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  XOR2_X1   g253(.A(G71gat), .B(G99gat), .Z(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT30), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G227gat), .A2(G233gat), .ZN(new_n457_));
  XOR2_X1   g256(.A(new_n456_), .B(new_n457_), .Z(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G15gat), .B(G43gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT31), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n374_), .A2(new_n286_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n374_), .A2(new_n286_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n461_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NOR3_X1   g264(.A1(new_n462_), .A2(new_n463_), .A3(new_n461_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n459_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n466_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(new_n458_), .A3(new_n464_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n454_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n423_), .A2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n471_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n451_), .ZN(new_n475_));
  NOR3_X1   g274(.A1(new_n435_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n434_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n475_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n443_), .A2(new_n448_), .A3(new_n451_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n478_), .A2(new_n479_), .A3(new_n470_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n474_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n413_), .ZN(new_n482_));
  OR2_X1    g281(.A1(new_n396_), .A2(KEYINPUT27), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n307_), .B(KEYINPUT99), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n419_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n485_), .A2(KEYINPUT27), .A3(new_n384_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .A4(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n473_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT13), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G120gat), .B(G148gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT5), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(G176gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(new_n353_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G57gat), .B(G64gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT11), .ZN(new_n495_));
  XOR2_X1   g294(.A(G71gat), .B(G78gat), .Z(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  OR2_X1    g296(.A1(new_n494_), .A2(KEYINPUT11), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G99gat), .A2(G106gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT6), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT6), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n502_), .A2(G99gat), .A3(G106gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT68), .ZN(new_n505_));
  INV_X1    g304(.A(G99gat), .ZN(new_n506_));
  INV_X1    g305(.A(G106gat), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(new_n507_), .A3(KEYINPUT66), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT7), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT7), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n510_), .A2(new_n506_), .A3(new_n507_), .A4(KEYINPUT66), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT68), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n501_), .A2(new_n503_), .A3(new_n512_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n505_), .A2(new_n509_), .A3(new_n511_), .A4(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G85gat), .B(G92gat), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n509_), .A2(new_n504_), .A3(KEYINPUT67), .A4(new_n511_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT8), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n509_), .A2(new_n504_), .A3(new_n511_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT67), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n515_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  AOI22_X1  g322(.A1(KEYINPUT8), .A2(new_n517_), .B1(new_n520_), .B2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT64), .B(G85gat), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT9), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  AOI22_X1  g326(.A1(new_n527_), .A2(G92gat), .B1(KEYINPUT9), .B2(G85gat), .ZN(new_n528_));
  NAND3_X1  g327(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT65), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(KEYINPUT10), .B(G99gat), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n504_), .B1(new_n532_), .B2(G106gat), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n499_), .B1(new_n524_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT69), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n497_), .A2(new_n498_), .ZN(new_n537_));
  OAI221_X1 g336(.A(new_n504_), .B1(G106gat), .B2(new_n532_), .C1(new_n528_), .C2(new_n530_), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n523_), .A2(new_n519_), .A3(new_n518_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n519_), .B1(new_n514_), .B2(new_n516_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n537_), .B(new_n538_), .C1(new_n539_), .C2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n535_), .A2(new_n536_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(G230gat), .ZN(new_n543_));
  INV_X1    g342(.A(G233gat), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  OAI211_X1 g344(.A(KEYINPUT69), .B(new_n499_), .C1(new_n524_), .C2(new_n534_), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n542_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n535_), .A2(KEYINPUT12), .A3(new_n541_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT12), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n549_), .B(new_n499_), .C1(new_n524_), .C2(new_n534_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n545_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n493_), .B1(new_n547_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n548_), .A2(new_n550_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n545_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n542_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n493_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n552_), .A2(new_n558_), .A3(KEYINPUT70), .ZN(new_n559_));
  AOI21_X1  g358(.A(KEYINPUT70), .B1(new_n552_), .B2(new_n558_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n489_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT71), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT70), .ZN(new_n563_));
  NOR3_X1   g362(.A1(new_n547_), .A2(new_n551_), .A3(new_n493_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n557_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n563_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n552_), .A2(new_n558_), .A3(KEYINPUT70), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(KEYINPUT13), .A3(new_n567_), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n561_), .A2(new_n562_), .A3(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n562_), .B1(new_n561_), .B2(new_n568_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n245_), .B(new_n488_), .C1(new_n569_), .C2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n229_), .B1(new_n524_), .B2(new_n534_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT73), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G232gat), .A2(G233gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT34), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n574_), .A2(KEYINPUT35), .A3(new_n576_), .ZN(new_n577_));
  OR3_X1    g376(.A1(new_n524_), .A2(new_n212_), .A3(new_n534_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n576_), .A2(KEYINPUT35), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n580_), .A2(KEYINPUT72), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(KEYINPUT72), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n578_), .A2(new_n572_), .A3(new_n581_), .A4(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n577_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G190gat), .B(G218gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(G134gat), .ZN(new_n587_));
  INV_X1    g386(.A(G162gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT36), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n577_), .A2(new_n583_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n585_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n577_), .A2(new_n583_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n589_), .ZN(new_n595_));
  OAI22_X1  g394(.A1(new_n594_), .A2(new_n584_), .B1(KEYINPUT36), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT37), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n593_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n597_), .B1(new_n593_), .B2(new_n596_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n499_), .B(new_n219_), .ZN(new_n602_));
  AND2_X1   g401(.A1(G231gat), .A2(G233gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G127gat), .B(G155gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT16), .ZN(new_n606_));
  INV_X1    g405(.A(G183gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(G211gat), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT17), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n610_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n604_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT75), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n604_), .A2(KEYINPUT74), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n604_), .A2(KEYINPUT74), .ZN(new_n616_));
  OR3_X1    g415(.A1(new_n615_), .A2(new_n616_), .A3(new_n611_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n614_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n601_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n571_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n622_), .A2(new_n214_), .A3(new_n413_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT38), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n593_), .A2(new_n596_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n619_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n571_), .A2(new_n482_), .A3(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n624_), .B1(new_n214_), .B2(new_n628_), .ZN(G1324gat));
  INV_X1    g428(.A(KEYINPUT40), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT39), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n483_), .A2(new_n486_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n571_), .A2(new_n633_), .A3(new_n627_), .ZN(new_n634_));
  OAI211_X1 g433(.A(KEYINPUT100), .B(new_n631_), .C1(new_n634_), .C2(new_n215_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n622_), .A2(new_n215_), .A3(new_n632_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n245_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n559_), .A2(new_n560_), .A3(new_n489_), .ZN(new_n638_));
  AOI21_X1  g437(.A(KEYINPUT13), .B1(new_n566_), .B2(new_n567_), .ZN(new_n639_));
  OAI21_X1  g438(.A(KEYINPUT71), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n561_), .A2(new_n568_), .A3(new_n562_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n637_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n642_), .A2(new_n632_), .A3(new_n488_), .A4(new_n626_), .ZN(new_n643_));
  OR2_X1    g442(.A1(new_n631_), .A2(KEYINPUT100), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n631_), .A2(KEYINPUT100), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n643_), .A2(G8gat), .A3(new_n644_), .A4(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n635_), .A2(new_n636_), .A3(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(KEYINPUT102), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT101), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT102), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n635_), .A2(new_n650_), .A3(new_n636_), .A4(new_n646_), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n648_), .A2(new_n649_), .A3(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n649_), .B1(new_n648_), .B2(new_n651_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n630_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n648_), .A2(new_n651_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(KEYINPUT101), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n648_), .A2(new_n649_), .A3(new_n651_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n656_), .A2(KEYINPUT40), .A3(new_n657_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n654_), .A2(new_n658_), .ZN(G1325gat));
  INV_X1    g458(.A(G15gat), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n571_), .A2(new_n627_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n661_), .B2(new_n471_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT41), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n622_), .A2(new_n660_), .A3(new_n471_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1326gat));
  INV_X1    g464(.A(G22gat), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n622_), .A2(new_n666_), .A3(new_n454_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n666_), .B1(new_n661_), .B2(new_n454_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n668_), .A2(new_n670_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n667_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT104), .Z(G1327gat));
  INV_X1    g473(.A(KEYINPUT107), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n600_), .B1(new_n473_), .B2(new_n487_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n676_), .B2(KEYINPUT106), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT43), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n676_), .A2(new_n675_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n675_), .B(new_n680_), .C1(new_n676_), .C2(KEYINPUT106), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n678_), .A2(new_n679_), .A3(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n640_), .A2(new_n641_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n683_), .A2(new_n245_), .A3(new_n619_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n642_), .A2(KEYINPUT105), .A3(new_n619_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n682_), .A2(new_n688_), .A3(KEYINPUT44), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT44), .B1(new_n682_), .B2(new_n688_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n689_), .A2(new_n690_), .A3(new_n482_), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n691_), .A2(KEYINPUT108), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(KEYINPUT108), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n692_), .A2(G29gat), .A3(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n619_), .A2(new_n625_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n571_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n482_), .A2(G29gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n694_), .B1(new_n697_), .B2(new_n698_), .ZN(G1328gat));
  NAND2_X1  g498(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT110), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT46), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(G36gat), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n689_), .A2(new_n690_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n705_), .B2(new_n632_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n696_), .A2(new_n704_), .A3(new_n632_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT109), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT109), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n696_), .A2(new_n709_), .A3(new_n704_), .A4(new_n632_), .ZN(new_n710_));
  AOI21_X1  g509(.A(KEYINPUT45), .B1(new_n708_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n708_), .A2(KEYINPUT45), .A3(new_n710_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n700_), .B(new_n703_), .C1(new_n706_), .C2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n690_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n682_), .A2(new_n688_), .A3(KEYINPUT44), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n716_), .A2(new_n632_), .A3(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(G36gat), .ZN(new_n719_));
  INV_X1    g518(.A(new_n713_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n720_), .A2(new_n711_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n719_), .A2(new_n721_), .A3(new_n701_), .A4(new_n702_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n715_), .A2(new_n722_), .ZN(G1329gat));
  NAND3_X1  g522(.A1(new_n705_), .A2(G43gat), .A3(new_n471_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n204_), .B1(new_n697_), .B2(new_n470_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g526(.A1(new_n696_), .A2(new_n202_), .A3(new_n454_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n705_), .A2(new_n454_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(new_n202_), .ZN(G1331gat));
  NOR2_X1   g529(.A1(new_n683_), .A2(new_n245_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(new_n488_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n732_), .A2(new_n621_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n482_), .B1(new_n734_), .B2(KEYINPUT111), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n735_), .B1(KEYINPUT111), .B2(new_n734_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n732_), .A2(new_n627_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n482_), .A2(new_n250_), .ZN(new_n738_));
  AOI22_X1  g537(.A1(new_n736_), .A2(new_n250_), .B1(new_n737_), .B2(new_n738_), .ZN(G1332gat));
  INV_X1    g538(.A(G64gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n737_), .B2(new_n632_), .ZN(new_n741_));
  XOR2_X1   g540(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n742_));
  XNOR2_X1  g541(.A(new_n741_), .B(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n733_), .A2(new_n740_), .A3(new_n632_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1333gat));
  INV_X1    g544(.A(G71gat), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n746_), .B1(new_n737_), .B2(new_n471_), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n747_), .B(KEYINPUT49), .Z(new_n748_));
  NAND3_X1  g547(.A1(new_n733_), .A2(new_n746_), .A3(new_n471_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1334gat));
  INV_X1    g549(.A(G78gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n737_), .B2(new_n454_), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n752_), .B(KEYINPUT50), .Z(new_n753_));
  NAND3_X1  g552(.A1(new_n733_), .A2(new_n751_), .A3(new_n454_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1335gat));
  NOR2_X1   g554(.A1(new_n732_), .A2(new_n695_), .ZN(new_n756_));
  AOI21_X1  g555(.A(G85gat), .B1(new_n756_), .B2(new_n413_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n682_), .A2(new_n619_), .A3(new_n731_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n482_), .A2(new_n525_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n757_), .B1(new_n758_), .B2(new_n759_), .ZN(G1336gat));
  AOI21_X1  g559(.A(G92gat), .B1(new_n756_), .B2(new_n632_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n632_), .A2(G92gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n758_), .B2(new_n762_), .ZN(G1337gat));
  NAND2_X1  g562(.A1(new_n758_), .A2(new_n471_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n470_), .A2(new_n532_), .ZN(new_n765_));
  AOI22_X1  g564(.A1(new_n764_), .A2(G99gat), .B1(new_n756_), .B2(new_n765_), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT51), .Z(G1338gat));
  XNOR2_X1  g566(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n682_), .A2(new_n454_), .A3(new_n619_), .A4(new_n731_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(G106gat), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT52), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n756_), .A2(new_n507_), .A3(new_n454_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n768_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n770_), .A2(KEYINPUT52), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n775_), .B1(new_n769_), .B2(G106gat), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n768_), .B(new_n772_), .C1(new_n774_), .C2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n773_), .A2(new_n778_), .ZN(G1339gat));
  INV_X1    g578(.A(G113gat), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n632_), .A2(new_n482_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n474_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n555_), .A2(KEYINPUT115), .A3(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n787_), .B1(new_n551_), .B2(KEYINPUT55), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n548_), .A2(new_n545_), .A3(new_n550_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n551_), .A2(KEYINPUT55), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n786_), .A2(new_n788_), .A3(new_n789_), .A4(new_n790_), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n791_), .A2(KEYINPUT56), .A3(new_n493_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT56), .B1(new_n791_), .B2(new_n493_), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n245_), .B(new_n558_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n230_), .A2(new_n222_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n220_), .A2(new_n221_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n241_), .A3(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n244_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT116), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n798_), .B(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n800_), .B1(new_n560_), .B2(new_n559_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n625_), .B1(new_n794_), .B2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT117), .B1(KEYINPUT118), .B2(KEYINPUT57), .ZN(new_n803_));
  OR2_X1    g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT118), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n802_), .B2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n804_), .B1(new_n807_), .B2(KEYINPUT57), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n800_), .B(new_n558_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT58), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n601_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n618_), .B1(new_n808_), .B2(new_n811_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n618_), .A2(new_n561_), .A3(new_n637_), .A4(new_n568_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n814_));
  OR2_X1    g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n814_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n601_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(KEYINPUT54), .ZN(new_n818_));
  OAI211_X1 g617(.A(KEYINPUT120), .B(new_n784_), .C1(new_n812_), .C2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT59), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n817_), .B(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n824_));
  AOI211_X1 g623(.A(KEYINPUT117), .B(new_n625_), .C1(new_n794_), .C2(new_n801_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n825_), .B2(new_n805_), .ZN(new_n826_));
  AOI22_X1  g625(.A1(new_n826_), .A2(new_n804_), .B1(new_n601_), .B2(new_n810_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n823_), .B1(new_n827_), .B2(new_n618_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n828_), .A2(KEYINPUT120), .A3(KEYINPUT59), .A4(new_n784_), .ZN(new_n829_));
  AOI211_X1 g628(.A(new_n780_), .B(new_n637_), .C1(new_n821_), .C2(new_n829_), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n245_), .B(new_n784_), .C1(new_n812_), .C2(new_n818_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n780_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n831_), .A2(KEYINPUT119), .A3(new_n780_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n830_), .A2(new_n836_), .ZN(G1340gat));
  NOR2_X1   g636(.A1(new_n812_), .A2(new_n818_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n838_), .A2(new_n783_), .ZN(new_n839_));
  XOR2_X1   g638(.A(KEYINPUT121), .B(G120gat), .Z(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n683_), .B2(KEYINPUT60), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n839_), .B(new_n841_), .C1(KEYINPUT60), .C2(new_n840_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n683_), .B1(new_n821_), .B2(new_n829_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n840_), .ZN(G1341gat));
  AOI21_X1  g643(.A(G127gat), .B1(new_n839_), .B2(new_n618_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n619_), .B1(new_n821_), .B2(new_n829_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g646(.A(G134gat), .B1(new_n839_), .B2(new_n625_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n600_), .B1(new_n821_), .B2(new_n829_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(G134gat), .ZN(G1343gat));
  INV_X1    g649(.A(new_n480_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n781_), .A2(new_n851_), .ZN(new_n852_));
  XOR2_X1   g651(.A(new_n852_), .B(KEYINPUT122), .Z(new_n853_));
  INV_X1    g652(.A(new_n812_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n853_), .B1(new_n854_), .B2(new_n823_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n245_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g656(.A(new_n683_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n855_), .A2(new_n858_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g659(.A1(new_n855_), .A2(new_n618_), .ZN(new_n861_));
  XOR2_X1   g660(.A(KEYINPUT61), .B(G155gat), .Z(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT123), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n861_), .B(new_n863_), .ZN(G1346gat));
  AOI21_X1  g663(.A(G162gat), .B1(new_n855_), .B2(new_n625_), .ZN(new_n865_));
  NOR4_X1   g664(.A1(new_n838_), .A2(new_n588_), .A3(new_n600_), .A4(new_n853_), .ZN(new_n866_));
  OAI21_X1  g665(.A(KEYINPUT124), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n855_), .A2(G162gat), .A3(new_n601_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT124), .ZN(new_n869_));
  INV_X1    g668(.A(new_n625_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n838_), .A2(new_n870_), .A3(new_n853_), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n868_), .B(new_n869_), .C1(new_n871_), .C2(G162gat), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n867_), .A2(new_n872_), .ZN(G1347gat));
  NOR2_X1   g672(.A1(new_n633_), .A2(new_n474_), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n482_), .B(new_n874_), .C1(new_n812_), .C2(new_n818_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT125), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT125), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n828_), .A2(new_n877_), .A3(new_n482_), .A4(new_n874_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(KEYINPUT22), .B(G169gat), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n876_), .A2(new_n878_), .A3(new_n245_), .A4(new_n879_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n828_), .A2(new_n482_), .A3(new_n245_), .A4(new_n874_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT62), .ZN(new_n882_));
  AND3_X1   g681(.A1(new_n881_), .A2(new_n882_), .A3(G169gat), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n881_), .B2(G169gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n880_), .B1(new_n883_), .B2(new_n884_), .ZN(G1348gat));
  NOR3_X1   g684(.A1(new_n875_), .A2(new_n322_), .A3(new_n683_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n876_), .A2(new_n878_), .A3(new_n858_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(new_n322_), .ZN(G1349gat));
  NOR2_X1   g687(.A1(new_n619_), .A2(new_n318_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n876_), .A2(new_n878_), .A3(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n607_), .B1(new_n875_), .B2(new_n619_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1350gat));
  NAND4_X1  g691(.A1(new_n876_), .A2(new_n878_), .A3(new_n319_), .A4(new_n625_), .ZN(new_n893_));
  AND3_X1   g692(.A1(new_n876_), .A2(new_n601_), .A3(new_n878_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n894_), .B2(new_n368_), .ZN(G1351gat));
  NAND2_X1  g694(.A1(new_n851_), .A2(new_n482_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(KEYINPUT126), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n828_), .A2(new_n632_), .A3(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n637_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(new_n240_), .ZN(G1352gat));
  NOR2_X1   g699(.A1(new_n898_), .A2(new_n683_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(new_n353_), .ZN(G1353gat));
  INV_X1    g701(.A(new_n898_), .ZN(new_n903_));
  XOR2_X1   g702(.A(KEYINPUT63), .B(G211gat), .Z(new_n904_));
  NAND3_X1  g703(.A1(new_n903_), .A2(new_n618_), .A3(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n906_), .B1(new_n898_), .B2(new_n619_), .ZN(new_n907_));
  AND2_X1   g706(.A1(new_n905_), .A2(new_n907_), .ZN(G1354gat));
  AOI21_X1  g707(.A(G218gat), .B1(new_n903_), .B2(new_n625_), .ZN(new_n909_));
  INV_X1    g708(.A(G218gat), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n600_), .A2(new_n910_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(KEYINPUT127), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n909_), .B1(new_n903_), .B2(new_n912_), .ZN(G1355gat));
endmodule


