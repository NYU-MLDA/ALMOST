//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1 0 0 0 1 1 0 0 0 1 1 0 1 1 0 0 1 0 1 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n836_, new_n837_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n856_, new_n857_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n890_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT64), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G57gat), .B(G64gat), .ZN(new_n205_));
  AND2_X1   g004(.A1(new_n205_), .A2(KEYINPUT11), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(KEYINPUT11), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G71gat), .B(G78gat), .ZN(new_n208_));
  OR3_X1    g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n205_), .A2(new_n208_), .A3(KEYINPUT11), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT7), .ZN(new_n213_));
  INV_X1    g012(.A(G99gat), .ZN(new_n214_));
  INV_X1    g013(.A(G106gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT69), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n218_));
  AND3_X1   g017(.A1(new_n216_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n217_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT68), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT6), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT67), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT67), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT6), .ZN(new_n226_));
  AND2_X1   g025(.A1(G99gat), .A2(G106gat), .ZN(new_n227_));
  AND3_X1   g026(.A1(new_n224_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n227_), .B1(new_n224_), .B2(new_n226_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n222_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n225_), .A2(KEYINPUT6), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n223_), .A2(KEYINPUT67), .ZN(new_n232_));
  OAI22_X1  g031(.A1(new_n231_), .A2(new_n232_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n224_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(KEYINPUT68), .A3(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n221_), .A2(new_n230_), .A3(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(G85gat), .B(G92gat), .Z(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT70), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n236_), .A2(KEYINPUT70), .A3(new_n237_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n240_), .A2(KEYINPUT8), .A3(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n228_), .A2(new_n229_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n243_), .A2(new_n218_), .A3(new_n216_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT8), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(new_n245_), .A3(new_n237_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n242_), .A2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT10), .B(G99gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT65), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n249_), .A2(new_n215_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n237_), .A2(KEYINPUT9), .ZN(new_n251_));
  NAND2_X1  g050(.A1(KEYINPUT66), .A2(G85gat), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n252_), .A2(KEYINPUT9), .ZN(new_n253_));
  NOR2_X1   g052(.A1(KEYINPUT66), .A2(G85gat), .ZN(new_n254_));
  OAI21_X1  g053(.A(G92gat), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n243_), .A2(new_n251_), .A3(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n250_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n212_), .B1(new_n247_), .B2(new_n258_), .ZN(new_n259_));
  AOI211_X1 g058(.A(new_n211_), .B(new_n257_), .C1(new_n242_), .C2(new_n246_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n204_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  AND3_X1   g060(.A1(new_n236_), .A2(KEYINPUT70), .A3(new_n237_), .ZN(new_n262_));
  AOI21_X1  g061(.A(KEYINPUT70), .B1(new_n236_), .B2(new_n237_), .ZN(new_n263_));
  NOR3_X1   g062(.A1(new_n262_), .A2(new_n263_), .A3(new_n245_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n246_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n258_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(new_n211_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n257_), .B1(new_n242_), .B2(new_n246_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(new_n212_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n267_), .A2(KEYINPUT12), .A3(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT12), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n259_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(KEYINPUT71), .B1(new_n273_), .B2(new_n203_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n275_));
  AOI211_X1 g074(.A(new_n275_), .B(new_n204_), .C1(new_n270_), .C2(new_n272_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n261_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT72), .B(G204gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G120gat), .B(G148gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT5), .B(G176gat), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n280_), .B(new_n281_), .Z(new_n282_));
  NAND2_X1  g081(.A1(new_n277_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n282_), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n261_), .B(new_n284_), .C1(new_n274_), .C2(new_n276_), .ZN(new_n285_));
  AOI21_X1  g084(.A(KEYINPUT13), .B1(new_n283_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n283_), .A2(KEYINPUT13), .A3(new_n285_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n289_), .B(KEYINPUT73), .Z(new_n290_));
  OR2_X1    g089(.A1(G169gat), .A2(G176gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(KEYINPUT24), .A3(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT26), .B(G190gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT25), .B(G183gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT23), .ZN(new_n298_));
  XOR2_X1   g097(.A(KEYINPUT86), .B(KEYINPUT23), .Z(new_n299_));
  OAI21_X1  g098(.A(new_n298_), .B1(new_n299_), .B2(new_n297_), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n291_), .A2(KEYINPUT24), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n302_), .A2(KEYINPUT95), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n302_), .A2(KEYINPUT95), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n293_), .B(new_n296_), .C1(new_n303_), .C2(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(G183gat), .A2(G190gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n299_), .A2(new_n297_), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n297_), .A2(KEYINPUT23), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n306_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT97), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT22), .B(G169gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT96), .ZN(new_n313_));
  INV_X1    g112(.A(G176gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n309_), .A2(new_n310_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n311_), .A2(new_n292_), .A3(new_n315_), .A4(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G211gat), .B(G218gat), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT92), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(G204gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT91), .B1(new_n321_), .B2(G197gat), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(KEYINPUT21), .A3(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G197gat), .B(G204gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  OR2_X1    g124(.A1(new_n320_), .A2(KEYINPUT21), .ZN(new_n326_));
  INV_X1    g125(.A(new_n324_), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n320_), .A2(KEYINPUT21), .A3(new_n327_), .A4(new_n322_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n325_), .A2(new_n326_), .A3(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n305_), .A2(new_n317_), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT20), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G226gat), .A2(G233gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT19), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n300_), .B1(G183gat), .B2(G190gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n312_), .A2(new_n314_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(new_n335_), .A3(new_n292_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n307_), .A2(new_n308_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT85), .ZN(new_n338_));
  INV_X1    g137(.A(G183gat), .ZN(new_n339_));
  OR3_X1    g138(.A1(new_n338_), .A2(new_n339_), .A3(KEYINPUT25), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT25), .B1(new_n338_), .B2(new_n339_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(new_n294_), .A3(new_n341_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n337_), .A2(new_n293_), .A3(new_n301_), .A4(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n336_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n345_), .A2(new_n329_), .ZN(new_n346_));
  OR3_X1    g145(.A1(new_n331_), .A2(new_n333_), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT20), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n305_), .A2(new_n317_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n329_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n348_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n345_), .A2(new_n329_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(new_n333_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT18), .B(G64gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(G92gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G8gat), .B(G36gat), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n356_), .B(new_n357_), .Z(new_n358_));
  NAND3_X1  g157(.A1(new_n347_), .A2(new_n354_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n358_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n333_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n361_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n331_), .A2(new_n333_), .A3(new_n346_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n360_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(KEYINPUT27), .B1(new_n359_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n359_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n351_), .A2(new_n361_), .A3(new_n352_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n331_), .A2(KEYINPUT102), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT102), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n369_), .B1(new_n330_), .B2(KEYINPUT20), .ZN(new_n370_));
  NOR3_X1   g169(.A1(new_n368_), .A2(new_n346_), .A3(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n367_), .B1(new_n371_), .B2(new_n361_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n366_), .B1(new_n372_), .B2(new_n360_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n365_), .B1(new_n373_), .B2(KEYINPUT27), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G225gat), .A2(G233gat), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT4), .ZN(new_n377_));
  AND2_X1   g176(.A1(G155gat), .A2(G162gat), .ZN(new_n378_));
  NOR2_X1   g177(.A1(G155gat), .A2(G162gat), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(G141gat), .A2(G148gat), .ZN(new_n381_));
  XOR2_X1   g180(.A(new_n381_), .B(KEYINPUT3), .Z(new_n382_));
  NAND2_X1  g181(.A1(G141gat), .A2(G148gat), .ZN(new_n383_));
  XOR2_X1   g182(.A(new_n383_), .B(KEYINPUT2), .Z(new_n384_));
  OAI21_X1  g183(.A(new_n380_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT1), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n381_), .B1(new_n380_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n378_), .A2(KEYINPUT1), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n387_), .A2(new_n388_), .A3(new_n383_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n385_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n391_), .A2(KEYINPUT98), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G127gat), .B(G134gat), .ZN(new_n393_));
  INV_X1    g192(.A(G113gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(G120gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n393_), .B(G113gat), .ZN(new_n397_));
  INV_X1    g196(.A(G120gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n396_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT98), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n400_), .B1(new_n390_), .B2(new_n401_), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n392_), .A2(new_n402_), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n391_), .A2(new_n400_), .A3(KEYINPUT98), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n377_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n400_), .A2(new_n377_), .A3(new_n390_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT99), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n376_), .B1(new_n406_), .B2(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n392_), .A2(new_n402_), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n411_), .A2(new_n376_), .A3(new_n404_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT0), .B(G57gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(G85gat), .ZN(new_n415_));
  XOR2_X1   g214(.A(G1gat), .B(G29gat), .Z(new_n416_));
  XOR2_X1   g215(.A(new_n415_), .B(new_n416_), .Z(new_n417_));
  NAND3_X1  g216(.A1(new_n410_), .A2(new_n413_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n417_), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT4), .B1(new_n411_), .B2(new_n404_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n375_), .B1(new_n420_), .B2(new_n408_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n419_), .B1(new_n421_), .B2(new_n412_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n418_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G227gat), .A2(G233gat), .ZN(new_n424_));
  INV_X1    g223(.A(G15gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G71gat), .B(G99gat), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n344_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n344_), .A2(new_n428_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n426_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n431_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n426_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(new_n429_), .A3(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT87), .B(KEYINPUT30), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(G43gat), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n432_), .A2(new_n435_), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n437_), .B1(new_n432_), .B2(new_n435_), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT88), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n432_), .A2(new_n435_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n437_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT88), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n444_), .A2(new_n445_), .A3(new_n438_), .ZN(new_n446_));
  XOR2_X1   g245(.A(new_n400_), .B(KEYINPUT31), .Z(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n441_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n449_));
  OAI211_X1 g248(.A(KEYINPUT88), .B(new_n447_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n390_), .A2(KEYINPUT29), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT90), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT93), .ZN(new_n454_));
  INV_X1    g253(.A(G228gat), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n455_), .A2(KEYINPUT89), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n455_), .A2(KEYINPUT89), .ZN(new_n457_));
  OAI21_X1  g256(.A(G233gat), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NOR3_X1   g257(.A1(new_n453_), .A2(new_n454_), .A3(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n452_), .A2(KEYINPUT93), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n350_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n458_), .B1(new_n453_), .B2(new_n329_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n390_), .A2(KEYINPUT29), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G22gat), .B(G50gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT28), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n464_), .A2(new_n466_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT94), .ZN(new_n469_));
  OR3_X1    g268(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n463_), .A2(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n469_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G78gat), .B(G106gat), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n473_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n471_), .A2(new_n476_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n463_), .A2(new_n474_), .A3(new_n470_), .A4(new_n475_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n451_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n449_), .A2(new_n479_), .A3(new_n450_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n423_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n372_), .A2(KEYINPUT32), .A3(new_n358_), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n358_), .A2(KEYINPUT32), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n347_), .A2(new_n354_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n484_), .B(new_n423_), .C1(new_n485_), .C2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n375_), .B1(new_n406_), .B2(new_n409_), .ZN(new_n488_));
  OR3_X1    g287(.A1(new_n411_), .A2(KEYINPUT100), .A3(new_n404_), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT100), .B1(new_n411_), .B2(new_n404_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(new_n376_), .A3(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n488_), .A2(new_n491_), .A3(KEYINPUT33), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(new_n417_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  OAI211_X1 g293(.A(KEYINPUT33), .B(new_n419_), .C1(new_n421_), .C2(new_n412_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT33), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n410_), .A2(new_n496_), .A3(new_n413_), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n495_), .A2(new_n497_), .A3(new_n359_), .A4(new_n364_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT101), .B1(new_n494_), .B2(new_n498_), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n497_), .A2(new_n359_), .A3(new_n364_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT101), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n500_), .A2(new_n501_), .A3(new_n493_), .A4(new_n495_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n487_), .A2(new_n499_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n451_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n504_), .A2(new_n480_), .ZN(new_n505_));
  AOI22_X1  g304(.A1(new_n374_), .A2(new_n483_), .B1(new_n503_), .B2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G29gat), .B(G36gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G43gat), .B(G50gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT15), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G15gat), .B(G22gat), .ZN(new_n514_));
  INV_X1    g313(.A(G1gat), .ZN(new_n515_));
  INV_X1    g314(.A(G8gat), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT14), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n514_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G1gat), .B(G8gat), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n518_), .B(new_n519_), .Z(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n513_), .A2(KEYINPUT82), .A3(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G229gat), .A2(G233gat), .ZN(new_n523_));
  INV_X1    g322(.A(new_n511_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(new_n520_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT82), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n526_), .B1(new_n512_), .B2(new_n520_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n522_), .A2(new_n523_), .A3(new_n525_), .A4(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n511_), .B(new_n521_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n523_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n528_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G169gat), .B(G197gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT83), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(G113gat), .ZN(new_n535_));
  XOR2_X1   g334(.A(new_n535_), .B(G141gat), .Z(new_n536_));
  NAND2_X1  g335(.A1(new_n532_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n536_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n528_), .A2(new_n531_), .A3(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT84), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT84), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT103), .B1(new_n506_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n503_), .A2(new_n505_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n481_), .A2(new_n482_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n423_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n548_), .A2(new_n374_), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n547_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT103), .ZN(new_n552_));
  INV_X1    g351(.A(new_n545_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n546_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G231gat), .A2(G233gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n520_), .B(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(new_n211_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G127gat), .B(G155gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G183gat), .B(G211gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n559_), .A2(KEYINPUT17), .A3(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n559_), .A2(KEYINPUT17), .ZN(new_n566_));
  OR2_X1    g365(.A1(KEYINPUT81), .A2(KEYINPUT17), .ZN(new_n567_));
  NAND2_X1  g366(.A1(KEYINPUT81), .A2(KEYINPUT17), .ZN(new_n568_));
  AOI21_X1  g367(.A(KEYINPUT79), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(KEYINPUT79), .A2(KEYINPUT81), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(KEYINPUT17), .ZN(new_n571_));
  AOI22_X1  g370(.A1(new_n566_), .A2(new_n569_), .B1(new_n571_), .B2(new_n559_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n565_), .B1(new_n572_), .B2(new_n564_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT37), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n266_), .A2(new_n513_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n268_), .A2(new_n524_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n578_), .B(KEYINPUT74), .Z(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT34), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n577_), .A2(KEYINPUT35), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(KEYINPUT35), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n580_), .A2(KEYINPUT35), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n575_), .A2(new_n576_), .A3(new_n582_), .A4(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(KEYINPUT77), .B(G134gat), .ZN(new_n586_));
  INV_X1    g385(.A(G162gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G190gat), .B(G218gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n591_), .A2(KEYINPUT36), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(KEYINPUT36), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n585_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n574_), .B1(new_n594_), .B2(KEYINPUT78), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n585_), .A2(new_n592_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(new_n594_), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n595_), .A2(new_n597_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NOR4_X1   g400(.A1(new_n290_), .A2(new_n556_), .A3(new_n573_), .A4(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n602_), .A2(new_n515_), .A3(new_n423_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT38), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n289_), .A2(new_n541_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n573_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n597_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n607_), .B1(new_n547_), .B2(new_n550_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n605_), .A2(KEYINPUT104), .A3(new_n606_), .A4(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT104), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n608_), .A2(new_n540_), .A3(new_n288_), .A4(new_n287_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n610_), .B1(new_n611_), .B2(new_n573_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n549_), .B1(new_n609_), .B2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n604_), .B1(new_n515_), .B2(new_n613_), .ZN(G1324gat));
  NOR2_X1   g413(.A1(new_n611_), .A2(new_n573_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n374_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n516_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT39), .Z(new_n618_));
  NAND3_X1  g417(.A1(new_n602_), .A2(new_n516_), .A3(new_n616_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g420(.A1(new_n602_), .A2(new_n425_), .A3(new_n504_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n612_), .A2(new_n609_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(new_n504_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT105), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n624_), .A2(new_n625_), .A3(G15gat), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n451_), .B1(new_n612_), .B2(new_n609_), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT105), .B1(new_n627_), .B2(new_n425_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n626_), .A2(new_n628_), .A3(KEYINPUT41), .ZN(new_n629_));
  AOI21_X1  g428(.A(KEYINPUT41), .B1(new_n626_), .B2(new_n628_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n622_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(KEYINPUT106), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT106), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n633_), .B(new_n622_), .C1(new_n629_), .C2(new_n630_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(G1326gat));
  INV_X1    g434(.A(G22gat), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n636_), .B1(new_n623_), .B2(new_n480_), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n637_), .B(KEYINPUT42), .Z(new_n638_));
  NAND3_X1  g437(.A1(new_n602_), .A2(new_n636_), .A3(new_n480_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(G1327gat));
  NOR2_X1   g439(.A1(new_n597_), .A2(new_n606_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n642_), .B1(new_n546_), .B2(new_n554_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n289_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(G29gat), .B1(new_n645_), .B2(new_n423_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT43), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n601_), .A2(new_n647_), .A3(new_n551_), .ZN(new_n648_));
  OAI21_X1  g447(.A(KEYINPUT43), .B1(new_n506_), .B2(new_n600_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n650_), .A2(KEYINPUT44), .A3(new_n573_), .A4(new_n605_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT107), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n654_), .A2(new_n549_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n650_), .A2(new_n573_), .A3(new_n605_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT44), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n658_), .A2(G29gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n646_), .B1(new_n655_), .B2(new_n659_), .ZN(G1328gat));
  NOR2_X1   g459(.A1(new_n374_), .A2(G36gat), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n555_), .A2(new_n644_), .A3(new_n641_), .A4(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(KEYINPUT108), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT108), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n643_), .A2(new_n664_), .A3(new_n644_), .A4(new_n661_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n663_), .A2(KEYINPUT45), .A3(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n663_), .A2(new_n665_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT45), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n658_), .A2(new_n616_), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n651_), .A2(new_n652_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n651_), .A2(new_n652_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n670_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(G36gat), .ZN(new_n674_));
  OAI211_X1 g473(.A(new_n666_), .B(new_n669_), .C1(new_n673_), .C2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(KEYINPUT46), .B1(new_n675_), .B2(KEYINPUT109), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n374_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n674_), .B1(new_n653_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n669_), .A2(new_n666_), .ZN(new_n679_));
  OAI211_X1 g478(.A(KEYINPUT109), .B(KEYINPUT46), .C1(new_n678_), .C2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n676_), .A2(new_n681_), .ZN(G1329gat));
  NAND4_X1  g481(.A1(new_n653_), .A2(G43gat), .A3(new_n504_), .A4(new_n658_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n645_), .A2(new_n504_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n683_), .B1(G43gat), .B2(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g485(.A(G50gat), .B1(new_n645_), .B2(new_n480_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n654_), .A2(new_n479_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n658_), .A2(G50gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n687_), .B1(new_n688_), .B2(new_n689_), .ZN(G1331gat));
  NOR4_X1   g489(.A1(new_n506_), .A2(new_n573_), .A3(new_n607_), .A4(new_n553_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n290_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(G57gat), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n692_), .A2(new_n693_), .A3(new_n549_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n289_), .A2(new_n606_), .A3(new_n600_), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n695_), .A2(KEYINPUT110), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(KEYINPUT110), .ZN(new_n697_));
  AND4_X1   g496(.A1(new_n551_), .A2(new_n696_), .A3(new_n541_), .A4(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(new_n423_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(new_n693_), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n700_), .A2(KEYINPUT111), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(KEYINPUT111), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n694_), .B1(new_n701_), .B2(new_n702_), .ZN(G1332gat));
  INV_X1    g502(.A(G64gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n698_), .A2(new_n704_), .A3(new_n616_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT48), .ZN(new_n706_));
  INV_X1    g505(.A(new_n692_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(new_n616_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n706_), .B1(new_n708_), .B2(G64gat), .ZN(new_n709_));
  AOI211_X1 g508(.A(KEYINPUT48), .B(new_n704_), .C1(new_n707_), .C2(new_n616_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n705_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT112), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n711_), .B(new_n712_), .ZN(G1333gat));
  INV_X1    g512(.A(G71gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n698_), .A2(new_n714_), .A3(new_n504_), .ZN(new_n715_));
  OAI21_X1  g514(.A(G71gat), .B1(new_n692_), .B2(new_n451_), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n716_), .A2(KEYINPUT113), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(KEYINPUT113), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n717_), .A2(KEYINPUT49), .A3(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT49), .B1(new_n717_), .B2(new_n718_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n715_), .B1(new_n719_), .B2(new_n720_), .ZN(G1334gat));
  NOR2_X1   g520(.A1(new_n479_), .A2(G78gat), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT114), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n698_), .A2(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(G78gat), .B1(new_n692_), .B2(new_n479_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n725_), .A2(KEYINPUT50), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n725_), .A2(KEYINPUT50), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n724_), .B1(new_n726_), .B2(new_n727_), .ZN(G1335gat));
  NOR3_X1   g527(.A1(new_n506_), .A2(new_n540_), .A3(new_n642_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n290_), .A2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(G85gat), .B1(new_n731_), .B2(new_n423_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n540_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n733_), .A2(new_n573_), .A3(new_n289_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n254_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n549_), .B1(new_n736_), .B2(new_n252_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT115), .Z(new_n738_));
  AOI21_X1  g537(.A(new_n732_), .B1(new_n735_), .B2(new_n738_), .ZN(G1336gat));
  AOI21_X1  g538(.A(G92gat), .B1(new_n731_), .B2(new_n616_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n734_), .A2(new_n374_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(G92gat), .B2(new_n741_), .ZN(G1337gat));
  INV_X1    g541(.A(KEYINPUT116), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n731_), .A2(new_n249_), .A3(new_n504_), .ZN(new_n744_));
  OAI21_X1  g543(.A(G99gat), .B1(new_n734_), .B2(new_n451_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n743_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n744_), .A2(new_n743_), .A3(new_n745_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g549(.A1(new_n731_), .A2(new_n215_), .A3(new_n480_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n733_), .A2(new_n573_), .A3(new_n480_), .A4(new_n289_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n752_), .A2(new_n753_), .A3(G106gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n752_), .B2(G106gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT117), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT117), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n751_), .B(new_n758_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n757_), .A2(KEYINPUT53), .A3(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT53), .B1(new_n757_), .B2(new_n759_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n760_), .A2(new_n761_), .ZN(G1339gat));
  AND3_X1   g561(.A1(new_n545_), .A2(KEYINPUT118), .A3(new_n606_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n289_), .A2(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(KEYINPUT118), .B1(new_n545_), .B2(new_n606_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n764_), .A2(new_n600_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT54), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT54), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n764_), .A2(new_n769_), .A3(new_n600_), .A4(new_n766_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n268_), .A2(KEYINPUT12), .A3(new_n212_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n259_), .A2(new_n260_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n773_), .B1(new_n774_), .B2(KEYINPUT12), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n275_), .B1(new_n775_), .B2(new_n204_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n204_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT71), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT55), .B1(new_n776_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(KEYINPUT55), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n780_), .B1(new_n203_), .B2(new_n273_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n282_), .B1(new_n779_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT56), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n785_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n273_), .A2(new_n203_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n787_), .B1(KEYINPUT55), .B2(new_n777_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n789_), .A2(KEYINPUT56), .A3(new_n282_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n784_), .A2(new_n790_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n522_), .A2(new_n530_), .A3(new_n525_), .A4(new_n527_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n529_), .A2(new_n523_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n792_), .A2(new_n536_), .A3(new_n793_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n794_), .A2(new_n539_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n285_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT119), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n285_), .A2(KEYINPUT119), .A3(new_n795_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n791_), .A2(new_n800_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n600_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  AND4_X1   g602(.A1(KEYINPUT121), .A2(new_n791_), .A3(KEYINPUT58), .A4(new_n800_), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n784_), .A2(new_n790_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT121), .B1(new_n805_), .B2(KEYINPUT58), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n803_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT122), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n285_), .A2(new_n540_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n810_), .B1(new_n784_), .B2(new_n790_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n795_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n812_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n597_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(KEYINPUT57), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n803_), .B(KEYINPUT122), .C1(new_n804_), .C2(new_n806_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n809_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n772_), .B1(new_n817_), .B2(new_n573_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n616_), .A2(new_n549_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n482_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(KEYINPUT123), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n818_), .A2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(G113gat), .B1(new_n824_), .B2(new_n540_), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT59), .B1(new_n818_), .B2(new_n823_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n823_), .A2(KEYINPUT59), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n606_), .B1(new_n815_), .B2(new_n807_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n827_), .B1(new_n828_), .B2(new_n772_), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n826_), .A2(G113gat), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n825_), .B1(new_n830_), .B2(new_n553_), .ZN(G1340gat));
  OAI21_X1  g630(.A(new_n398_), .B1(new_n644_), .B2(KEYINPUT60), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n824_), .B(new_n832_), .C1(KEYINPUT60), .C2(new_n398_), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n826_), .A2(new_n290_), .A3(new_n829_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n833_), .B1(new_n834_), .B2(new_n398_), .ZN(G1341gat));
  AOI21_X1  g634(.A(G127gat), .B1(new_n824_), .B2(new_n606_), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n826_), .A2(G127gat), .A3(new_n829_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(new_n606_), .ZN(G1342gat));
  NOR3_X1   g637(.A1(new_n818_), .A2(new_n597_), .A3(new_n823_), .ZN(new_n839_));
  OAI21_X1  g638(.A(KEYINPUT124), .B1(new_n839_), .B2(G134gat), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n817_), .A2(new_n573_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n771_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n842_), .A2(new_n607_), .A3(new_n822_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT124), .ZN(new_n844_));
  INV_X1    g643(.A(G134gat), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n843_), .A2(new_n844_), .A3(new_n845_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n826_), .A2(G134gat), .A3(new_n601_), .A4(new_n829_), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n840_), .A2(new_n846_), .A3(new_n847_), .ZN(G1343gat));
  INV_X1    g647(.A(new_n481_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n819_), .A2(new_n849_), .ZN(new_n850_));
  XOR2_X1   g649(.A(new_n850_), .B(KEYINPUT125), .Z(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(new_n841_), .B2(new_n771_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n540_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g654(.A1(new_n853_), .A2(new_n290_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(KEYINPUT126), .B(G148gat), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n856_), .B(new_n857_), .ZN(G1345gat));
  NAND2_X1  g657(.A1(new_n853_), .A2(new_n606_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(KEYINPUT61), .B(G155gat), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n859_), .B(new_n860_), .ZN(G1346gat));
  AOI21_X1  g660(.A(G162gat), .B1(new_n853_), .B2(new_n607_), .ZN(new_n862_));
  NOR4_X1   g661(.A1(new_n818_), .A2(new_n587_), .A3(new_n600_), .A4(new_n852_), .ZN(new_n863_));
  OAI21_X1  g662(.A(KEYINPUT127), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n842_), .A2(G162gat), .A3(new_n601_), .A4(new_n851_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT127), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n818_), .A2(new_n597_), .A3(new_n852_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n865_), .B(new_n866_), .C1(new_n867_), .C2(G162gat), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n864_), .A2(new_n868_), .ZN(G1347gat));
  NOR2_X1   g668(.A1(new_n374_), .A2(new_n423_), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n820_), .B(new_n870_), .C1(new_n828_), .C2(new_n772_), .ZN(new_n871_));
  OAI21_X1  g670(.A(G169gat), .B1(new_n871_), .B2(new_n541_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT62), .ZN(new_n873_));
  OR2_X1    g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n871_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n875_), .A2(new_n313_), .A3(new_n540_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n872_), .A2(new_n873_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n874_), .A2(new_n876_), .A3(new_n877_), .ZN(G1348gat));
  AOI21_X1  g677(.A(G176gat), .B1(new_n875_), .B2(new_n289_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n870_), .A2(new_n820_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n818_), .A2(new_n880_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n881_), .A2(new_n290_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n879_), .B1(new_n882_), .B2(G176gat), .ZN(G1349gat));
  NOR3_X1   g682(.A1(new_n871_), .A2(new_n573_), .A3(new_n295_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n881_), .A2(new_n606_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(new_n339_), .ZN(G1350gat));
  OAI21_X1  g685(.A(G190gat), .B1(new_n871_), .B2(new_n600_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n607_), .A2(new_n294_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n871_), .B2(new_n888_), .ZN(G1351gat));
  NAND4_X1  g688(.A1(new_n842_), .A2(new_n849_), .A3(new_n540_), .A4(new_n870_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(G197gat), .ZN(G1352gat));
  NAND4_X1  g690(.A1(new_n842_), .A2(new_n849_), .A3(new_n290_), .A4(new_n870_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g692(.A1(new_n818_), .A2(new_n481_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(KEYINPUT63), .B(G211gat), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n894_), .A2(new_n606_), .A3(new_n870_), .A4(new_n895_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n842_), .A2(new_n849_), .A3(new_n870_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n573_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n896_), .B1(new_n898_), .B2(new_n899_), .ZN(G1354gat));
  INV_X1    g699(.A(G218gat), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n897_), .A2(new_n901_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n894_), .A2(new_n607_), .A3(new_n870_), .ZN(new_n903_));
  AOI22_X1  g702(.A1(new_n902_), .A2(new_n601_), .B1(new_n903_), .B2(new_n901_), .ZN(G1355gat));
endmodule


