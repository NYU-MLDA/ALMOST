//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1 1 0 0 0 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 0 1 1 1 0 1 0 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n857_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT6), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(KEYINPUT10), .B(G99gat), .Z(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT64), .ZN(new_n206_));
  INV_X1    g005(.A(G106gat), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n204_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G85gat), .A2(G92gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G85gat), .A2(G92gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n209_), .B1(new_n211_), .B2(KEYINPUT9), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT9), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n213_), .B1(new_n210_), .B2(new_n214_), .ZN(new_n215_));
  AND3_X1   g014(.A1(new_n210_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n212_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n208_), .A2(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n211_), .A2(new_n209_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G99gat), .A2(G106gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT7), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n221_), .B1(new_n224_), .B2(new_n204_), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n225_), .A2(KEYINPUT8), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(KEYINPUT8), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n220_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G29gat), .B(G36gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT70), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G43gat), .B(G50gat), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n230_), .A2(KEYINPUT70), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n230_), .A2(KEYINPUT70), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(new_n236_), .A3(new_n232_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n234_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT15), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n234_), .A2(KEYINPUT15), .A3(new_n237_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n229_), .A2(new_n242_), .A3(KEYINPUT71), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(KEYINPUT71), .B1(new_n229_), .B2(new_n242_), .ZN(new_n245_));
  OAI22_X1  g044(.A1(new_n244_), .A2(new_n245_), .B1(new_n229_), .B2(new_n238_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n229_), .A2(new_n242_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT71), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(KEYINPUT72), .B1(new_n249_), .B2(new_n243_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G232gat), .A2(G233gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT35), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n246_), .B1(new_n250_), .B2(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n253_), .A2(KEYINPUT35), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT72), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n257_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n254_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n256_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n255_), .B1(new_n260_), .B2(new_n246_), .ZN(new_n261_));
  XOR2_X1   g060(.A(G134gat), .B(G162gat), .Z(new_n262_));
  XNOR2_X1  g061(.A(G190gat), .B(G218gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT36), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n266_), .B(KEYINPUT73), .Z(new_n267_));
  XOR2_X1   g066(.A(new_n267_), .B(KEYINPUT74), .Z(new_n268_));
  NAND2_X1  g067(.A1(new_n261_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n264_), .B(KEYINPUT36), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n255_), .B(new_n270_), .C1(new_n260_), .C2(new_n246_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT76), .B1(new_n272_), .B2(KEYINPUT37), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT76), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT37), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n269_), .A2(new_n274_), .A3(new_n275_), .A4(new_n271_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n273_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT75), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n269_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n261_), .A2(KEYINPUT75), .A3(new_n268_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(new_n271_), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT37), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n277_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G57gat), .B(G64gat), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n284_), .A2(KEYINPUT11), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(KEYINPUT11), .ZN(new_n286_));
  XOR2_X1   g085(.A(G71gat), .B(G78gat), .Z(new_n287_));
  NAND3_X1  g086(.A1(new_n285_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n286_), .A2(new_n287_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G231gat), .A2(G233gat), .ZN(new_n291_));
  XOR2_X1   g090(.A(new_n290_), .B(new_n291_), .Z(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT77), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G15gat), .B(G22gat), .ZN(new_n294_));
  INV_X1    g093(.A(G1gat), .ZN(new_n295_));
  INV_X1    g094(.A(G8gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT14), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n294_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G1gat), .B(G8gat), .ZN(new_n299_));
  XOR2_X1   g098(.A(new_n298_), .B(new_n299_), .Z(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n293_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT17), .ZN(new_n303_));
  XOR2_X1   g102(.A(G127gat), .B(G155gat), .Z(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT16), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G183gat), .B(G211gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  OR3_X1    g106(.A1(new_n302_), .A2(new_n303_), .A3(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(KEYINPUT17), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n302_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n283_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT78), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n229_), .A2(new_n289_), .A3(new_n288_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(KEYINPUT12), .ZN(new_n316_));
  AOI22_X1  g115(.A1(new_n219_), .A2(new_n208_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n317_));
  OR3_X1    g116(.A1(new_n317_), .A2(KEYINPUT12), .A3(new_n290_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G230gat), .A2(G233gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n321_), .B1(new_n317_), .B2(new_n290_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT68), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n323_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n319_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n317_), .A2(new_n290_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT67), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n315_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n329_), .B(new_n321_), .C1(new_n328_), .C2(new_n315_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G120gat), .B(G148gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT5), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G176gat), .B(G204gat), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n332_), .B(new_n333_), .Z(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n326_), .A2(new_n330_), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n335_), .B1(new_n326_), .B2(new_n330_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  OR2_X1    g138(.A1(new_n339_), .A2(KEYINPUT13), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(KEYINPUT13), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT79), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n344_), .B1(new_n238_), .B2(new_n301_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n300_), .A2(KEYINPUT79), .A3(new_n237_), .A4(new_n234_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n242_), .A2(new_n301_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G229gat), .A2(G233gat), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n347_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  AOI22_X1  g149(.A1(new_n345_), .A2(new_n346_), .B1(new_n238_), .B2(new_n301_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n350_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G113gat), .B(G141gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G169gat), .B(G197gat), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n353_), .B(new_n354_), .Z(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n352_), .A2(new_n356_), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n350_), .B(new_n355_), .C1(new_n349_), .C2(new_n351_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G141gat), .A2(G148gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT86), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT86), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(G141gat), .A3(G148gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(G141gat), .ZN(new_n366_));
  INV_X1    g165(.A(G148gat), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n365_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(G155gat), .A2(G162gat), .ZN(new_n369_));
  AND2_X1   g168(.A1(G155gat), .A2(G162gat), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT1), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n369_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NOR3_X1   g171(.A1(new_n370_), .A2(KEYINPUT87), .A3(new_n371_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT87), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G155gat), .A2(G162gat), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n374_), .B1(new_n375_), .B2(KEYINPUT1), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n372_), .B1(new_n373_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n368_), .A2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n370_), .A2(new_n369_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n365_), .A2(KEYINPUT2), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT3), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n381_), .A2(new_n366_), .A3(new_n367_), .A4(KEYINPUT88), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT88), .ZN(new_n383_));
  OAI22_X1  g182(.A1(new_n383_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n384_));
  NAND3_X1  g183(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n382_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n379_), .B1(new_n380_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT29), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n378_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n389_), .A2(KEYINPUT28), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(KEYINPUT28), .ZN(new_n391_));
  INV_X1    g190(.A(G233gat), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT89), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n393_), .A2(G228gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(G228gat), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n392_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT90), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n390_), .A2(new_n391_), .A3(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n398_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G211gat), .B(G218gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(G197gat), .ZN(new_n405_));
  AND2_X1   g204(.A1(KEYINPUT92), .A2(G204gat), .ZN(new_n406_));
  NOR2_X1   g205(.A1(KEYINPUT92), .A2(G204gat), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n405_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT93), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  OAI211_X1 g209(.A(KEYINPUT93), .B(new_n405_), .C1(new_n406_), .C2(new_n407_), .ZN(new_n411_));
  INV_X1    g210(.A(G204gat), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n405_), .A2(KEYINPUT91), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n405_), .A2(KEYINPUT91), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n412_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n410_), .A2(new_n411_), .A3(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n404_), .B1(new_n416_), .B2(KEYINPUT21), .ZN(new_n417_));
  INV_X1    g216(.A(new_n407_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(KEYINPUT92), .A2(G204gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT94), .B1(new_n420_), .B2(new_n405_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT21), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT91), .B(G197gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(G204gat), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT94), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n418_), .A2(new_n425_), .A3(G197gat), .A4(new_n419_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n421_), .A2(new_n422_), .A3(new_n424_), .A4(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n421_), .A2(new_n424_), .A3(new_n426_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n403_), .A2(new_n422_), .ZN(new_n429_));
  AOI22_X1  g228(.A1(new_n417_), .A2(new_n427_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n388_), .B1(new_n378_), .B2(new_n387_), .ZN(new_n431_));
  OAI21_X1  g230(.A(G78gat), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n416_), .A2(KEYINPUT21), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n433_), .A2(new_n427_), .A3(new_n403_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n428_), .A2(new_n429_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(G78gat), .ZN(new_n437_));
  INV_X1    g236(.A(new_n431_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n432_), .A2(new_n439_), .A3(G106gat), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(G106gat), .B1(new_n432_), .B2(new_n439_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G22gat), .B(G50gat), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n441_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n443_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n432_), .A2(new_n439_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n207_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n445_), .B1(new_n447_), .B2(new_n440_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n402_), .B1(new_n444_), .B2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n443_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n447_), .A2(new_n440_), .A3(new_n445_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n450_), .A2(new_n451_), .A3(new_n401_), .ZN(new_n452_));
  AND2_X1   g251(.A1(new_n449_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT22), .ZN(new_n454_));
  INV_X1    g253(.A(G169gat), .ZN(new_n455_));
  INV_X1    g254(.A(G176gat), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n454_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G183gat), .A2(G190gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT23), .ZN(new_n461_));
  OR2_X1    g260(.A1(KEYINPUT80), .A2(G183gat), .ZN(new_n462_));
  INV_X1    g261(.A(G190gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(KEYINPUT80), .A2(G183gat), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n459_), .B1(new_n461_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT23), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n460_), .B(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT24), .B1(new_n455_), .B2(new_n456_), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NOR3_X1   g270(.A1(KEYINPUT81), .A2(G169gat), .A3(G176gat), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n469_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  OR3_X1    g272(.A1(KEYINPUT81), .A2(G169gat), .A3(G176gat), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n474_), .A2(KEYINPUT24), .A3(new_n470_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n468_), .B1(new_n473_), .B2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT26), .B(G190gat), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT25), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n478_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n477_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n466_), .B1(new_n476_), .B2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT30), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT83), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G227gat), .A2(G233gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT82), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G71gat), .B(G99gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(G15gat), .B(G43gat), .Z(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n485_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n483_), .A2(new_n484_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n485_), .A2(new_n493_), .A3(new_n491_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  OR2_X1    g294(.A1(new_n495_), .A2(KEYINPUT85), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(KEYINPUT85), .ZN(new_n497_));
  XOR2_X1   g296(.A(G127gat), .B(G134gat), .Z(new_n498_));
  XOR2_X1   g297(.A(G113gat), .B(G120gat), .Z(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G127gat), .B(G134gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G113gat), .B(G120gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n500_), .A2(KEYINPUT84), .A3(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT84), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n501_), .A2(new_n502_), .A3(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT31), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n496_), .A2(new_n497_), .A3(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G1gat), .B(G29gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(G85gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT0), .B(G57gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n378_), .A2(new_n387_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(new_n507_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n500_), .A2(new_n503_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n378_), .A2(new_n387_), .A3(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n516_), .A2(KEYINPUT4), .A3(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G225gat), .A2(G233gat), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n520_), .B(KEYINPUT97), .Z(new_n521_));
  AOI22_X1  g320(.A1(new_n378_), .A2(new_n387_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT4), .ZN(new_n523_));
  AOI21_X1  g322(.A(KEYINPUT98), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  AND4_X1   g323(.A1(KEYINPUT98), .A2(new_n515_), .A3(new_n523_), .A4(new_n507_), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n519_), .B(new_n521_), .C1(new_n524_), .C2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n516_), .A2(new_n518_), .A3(new_n520_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n514_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n526_), .A2(new_n514_), .A3(new_n527_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n508_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n495_), .A2(KEYINPUT85), .A3(new_n533_), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n509_), .A2(new_n532_), .A3(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(G8gat), .B(G36gat), .Z(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT18), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G64gat), .B(G92gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT20), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT25), .B(G183gat), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n468_), .B1(new_n477_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n473_), .A2(new_n475_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n461_), .B1(G183gat), .B2(G190gat), .ZN(new_n544_));
  INV_X1    g343(.A(new_n459_), .ZN(new_n545_));
  AOI22_X1  g344(.A1(new_n542_), .A2(new_n543_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n540_), .B1(new_n430_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT96), .ZN(new_n548_));
  INV_X1    g347(.A(new_n482_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n548_), .B1(new_n436_), .B2(new_n549_), .ZN(new_n550_));
  AOI211_X1 g349(.A(KEYINPUT96), .B(new_n482_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n547_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G226gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT100), .ZN(new_n556_));
  INV_X1    g355(.A(new_n546_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n436_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n555_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n434_), .A2(new_n435_), .A3(new_n482_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n558_), .A2(KEYINPUT20), .A3(new_n559_), .A4(new_n560_), .ZN(new_n561_));
  AOI22_X1  g360(.A1(new_n552_), .A2(new_n555_), .B1(new_n556_), .B2(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n540_), .B1(new_n436_), .B2(new_n557_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n563_), .A2(KEYINPUT100), .A3(new_n559_), .A4(new_n560_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n539_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n559_), .B(new_n547_), .C1(new_n550_), .C2(new_n551_), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n560_), .B(KEYINPUT20), .C1(new_n430_), .C2(new_n546_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(new_n555_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n566_), .A2(new_n539_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT27), .ZN(new_n570_));
  OAI21_X1  g369(.A(KEYINPUT102), .B1(new_n565_), .B2(new_n570_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n569_), .A2(KEYINPUT27), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n556_), .B1(new_n567_), .B2(new_n555_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n434_), .A2(new_n435_), .A3(new_n546_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(KEYINPUT20), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT96), .B1(new_n430_), .B2(new_n482_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n436_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n575_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n573_), .B(new_n564_), .C1(new_n559_), .C2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n539_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT102), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n572_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n571_), .A2(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n539_), .B1(new_n566_), .B2(new_n568_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(KEYINPUT27), .B1(new_n586_), .B2(new_n569_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(KEYINPUT103), .B1(new_n584_), .B2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT103), .ZN(new_n590_));
  AOI211_X1 g389(.A(new_n590_), .B(new_n587_), .C1(new_n571_), .C2(new_n583_), .ZN(new_n591_));
  OAI211_X1 g390(.A(new_n453_), .B(new_n535_), .C1(new_n589_), .C2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n539_), .A2(KEYINPUT32), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n593_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n566_), .A2(new_n568_), .A3(new_n593_), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n526_), .A2(new_n514_), .A3(new_n527_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n595_), .B1(new_n596_), .B2(new_n528_), .ZN(new_n597_));
  OAI21_X1  g396(.A(KEYINPUT101), .B1(new_n594_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n593_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n579_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT101), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n600_), .A2(new_n601_), .A3(new_n531_), .A4(new_n595_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT99), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n603_), .A2(KEYINPUT33), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n520_), .B(new_n519_), .C1(new_n524_), .C2(new_n525_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n516_), .A2(new_n518_), .A3(new_n521_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n607_), .A2(new_n513_), .ZN(new_n608_));
  AOI22_X1  g407(.A1(new_n596_), .A2(new_n605_), .B1(new_n606_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n530_), .A2(new_n604_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n609_), .A2(new_n610_), .A3(new_n569_), .A4(new_n586_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n598_), .A2(new_n602_), .A3(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(new_n453_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n531_), .B1(new_n449_), .B2(new_n452_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n565_), .A2(KEYINPUT102), .A3(new_n570_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n582_), .B1(new_n572_), .B2(new_n581_), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n614_), .B(new_n588_), .C1(new_n615_), .C2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n613_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n509_), .A2(new_n534_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n360_), .B1(new_n592_), .B2(new_n620_), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n314_), .A2(new_n343_), .A3(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n622_), .A2(new_n295_), .A3(new_n531_), .ZN(new_n623_));
  XOR2_X1   g422(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n272_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n626_), .B1(new_n592_), .B2(new_n620_), .ZN(new_n627_));
  AND4_X1   g426(.A1(new_n627_), .A2(new_n312_), .A3(new_n359_), .A4(new_n343_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT105), .Z(new_n629_));
  OAI21_X1  g428(.A(G1gat), .B1(new_n629_), .B2(new_n532_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n625_), .A2(new_n630_), .ZN(G1324gat));
  NOR2_X1   g430(.A1(new_n589_), .A2(new_n591_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n622_), .A2(new_n296_), .A3(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n628_), .A2(new_n632_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(G8gat), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT106), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT39), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT106), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n634_), .A2(new_n638_), .A3(G8gat), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n636_), .A2(new_n637_), .A3(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n637_), .B1(new_n636_), .B2(new_n639_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n633_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT40), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(G1325gat));
  OAI21_X1  g443(.A(G15gat), .B1(new_n629_), .B2(new_n619_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT41), .Z(new_n646_));
  INV_X1    g445(.A(G15gat), .ZN(new_n647_));
  INV_X1    g446(.A(new_n619_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n622_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n649_), .ZN(G1326gat));
  OAI21_X1  g449(.A(G22gat), .B1(new_n629_), .B2(new_n453_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT42), .ZN(new_n652_));
  INV_X1    g451(.A(G22gat), .ZN(new_n653_));
  INV_X1    g452(.A(new_n453_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n622_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n652_), .A2(new_n655_), .ZN(G1327gat));
  AND4_X1   g455(.A1(new_n626_), .A2(new_n621_), .A3(new_n311_), .A4(new_n343_), .ZN(new_n657_));
  AOI21_X1  g456(.A(G29gat), .B1(new_n657_), .B2(new_n531_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n592_), .A2(new_n620_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT43), .ZN(new_n660_));
  AOI22_X1  g459(.A1(new_n273_), .A2(new_n276_), .B1(new_n281_), .B2(KEYINPUT37), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n659_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(KEYINPUT107), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT107), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n659_), .A2(new_n661_), .A3(new_n664_), .A4(new_n660_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n659_), .A2(new_n661_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(KEYINPUT43), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n663_), .A2(new_n665_), .A3(new_n667_), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n342_), .A2(new_n312_), .A3(new_n360_), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n668_), .A2(KEYINPUT44), .A3(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n669_), .ZN(new_n671_));
  AOI21_X1  g470(.A(KEYINPUT44), .B1(new_n671_), .B2(KEYINPUT108), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT108), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n668_), .A2(new_n673_), .A3(new_n669_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n670_), .B1(new_n672_), .B2(new_n674_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n531_), .A2(G29gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n658_), .B1(new_n675_), .B2(new_n676_), .ZN(G1328gat));
  INV_X1    g476(.A(KEYINPUT46), .ZN(new_n678_));
  INV_X1    g477(.A(G36gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n679_), .B1(new_n675_), .B2(new_n632_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT110), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n632_), .A2(KEYINPUT109), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n632_), .A2(KEYINPUT109), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n685_), .A2(G36gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n681_), .B1(new_n657_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n657_), .A2(new_n686_), .A3(new_n681_), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n688_), .A2(KEYINPUT45), .A3(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT45), .B1(new_n688_), .B2(new_n689_), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n678_), .B1(new_n680_), .B2(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n690_), .A2(new_n691_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n632_), .ZN(new_n695_));
  AOI211_X1 g494(.A(new_n695_), .B(new_n670_), .C1(new_n672_), .C2(new_n674_), .ZN(new_n696_));
  OAI211_X1 g495(.A(KEYINPUT46), .B(new_n694_), .C1(new_n696_), .C2(new_n679_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n693_), .A2(new_n697_), .ZN(G1329gat));
  AOI21_X1  g497(.A(G43gat), .B1(new_n657_), .B2(new_n648_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n648_), .A2(G43gat), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n699_), .B1(new_n675_), .B2(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n703_), .ZN(new_n705_));
  AOI211_X1 g504(.A(new_n700_), .B(new_n670_), .C1(new_n672_), .C2(new_n674_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(new_n706_), .B2(new_n699_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n704_), .A2(new_n707_), .ZN(G1330gat));
  AOI21_X1  g507(.A(G50gat), .B1(new_n657_), .B2(new_n654_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n654_), .A2(G50gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n675_), .B2(new_n710_), .ZN(G1331gat));
  AOI21_X1  g510(.A(new_n359_), .B1(new_n592_), .B2(new_n620_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n314_), .A2(new_n342_), .A3(new_n712_), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n713_), .A2(KEYINPUT112), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(KEYINPUT112), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(G57gat), .B1(new_n716_), .B2(new_n531_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n311_), .A2(new_n359_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n627_), .A2(new_n342_), .A3(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n719_), .A2(G57gat), .A3(new_n531_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT113), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n717_), .A2(new_n721_), .ZN(G1332gat));
  INV_X1    g521(.A(G64gat), .ZN(new_n723_));
  INV_X1    g522(.A(new_n685_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n716_), .A2(new_n723_), .A3(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n723_), .B1(new_n719_), .B2(new_n724_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT48), .Z(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(G1333gat));
  NOR2_X1   g527(.A1(new_n619_), .A2(G71gat), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT114), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n716_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(G71gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n719_), .B2(new_n648_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT49), .Z(new_n734_));
  NAND2_X1  g533(.A1(new_n731_), .A2(new_n734_), .ZN(G1334gat));
  NOR2_X1   g534(.A1(new_n453_), .A2(G78gat), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n714_), .A2(new_n715_), .A3(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n719_), .A2(new_n654_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(G78gat), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT50), .Z(new_n740_));
  OR3_X1    g539(.A1(new_n737_), .A2(KEYINPUT115), .A3(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(KEYINPUT115), .B1(new_n737_), .B2(new_n740_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1335gat));
  NOR3_X1   g542(.A1(new_n343_), .A2(new_n312_), .A3(new_n359_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n668_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(G85gat), .B1(new_n746_), .B2(new_n532_), .ZN(new_n747_));
  AND4_X1   g546(.A1(new_n626_), .A2(new_n712_), .A3(new_n311_), .A4(new_n342_), .ZN(new_n748_));
  INV_X1    g547(.A(G85gat), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n748_), .A2(new_n749_), .A3(new_n531_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n747_), .A2(new_n750_), .ZN(G1336gat));
  OAI21_X1  g550(.A(G92gat), .B1(new_n746_), .B2(new_n685_), .ZN(new_n752_));
  INV_X1    g551(.A(G92gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n748_), .A2(new_n753_), .A3(new_n632_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(G1337gat));
  NAND2_X1  g554(.A1(new_n745_), .A2(new_n648_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n648_), .A2(new_n206_), .ZN(new_n757_));
  AOI22_X1  g556(.A1(new_n756_), .A2(G99gat), .B1(new_n748_), .B2(new_n757_), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g558(.A1(new_n748_), .A2(new_n207_), .A3(new_n654_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n745_), .A2(new_n654_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n762_), .B2(G106gat), .ZN(new_n763_));
  AOI211_X1 g562(.A(KEYINPUT52), .B(new_n207_), .C1(new_n745_), .C2(new_n654_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n760_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT53), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n767_), .B(new_n760_), .C1(new_n763_), .C2(new_n764_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1339gat));
  INV_X1    g568(.A(KEYINPUT57), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n336_), .A2(new_n359_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT116), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n771_), .B(new_n772_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n319_), .A2(new_n324_), .A3(KEYINPUT55), .A4(new_n325_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT117), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  AOI22_X1  g575(.A1(new_n316_), .A2(new_n318_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n777_), .A2(KEYINPUT117), .A3(KEYINPUT55), .A4(new_n324_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n320_), .B1(new_n319_), .B2(new_n327_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(new_n326_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n779_), .A2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT56), .B1(new_n783_), .B2(new_n334_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT56), .ZN(new_n785_));
  AOI211_X1 g584(.A(new_n785_), .B(new_n335_), .C1(new_n779_), .C2(new_n782_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n773_), .B1(new_n784_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n349_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n347_), .A2(new_n348_), .A3(new_n788_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n789_), .B(new_n356_), .C1(new_n788_), .C2(new_n351_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n358_), .B(new_n790_), .C1(new_n337_), .C2(new_n338_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n787_), .A2(new_n791_), .ZN(new_n792_));
  OAI211_X1 g591(.A(KEYINPUT118), .B(new_n770_), .C1(new_n792_), .C2(new_n626_), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n336_), .A2(new_n358_), .A3(new_n790_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n794_), .B1(new_n784_), .B2(new_n786_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT58), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  OAI211_X1 g596(.A(KEYINPUT58), .B(new_n794_), .C1(new_n784_), .C2(new_n786_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n661_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n626_), .B1(new_n787_), .B2(new_n791_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT118), .ZN(new_n801_));
  OAI21_X1  g600(.A(KEYINPUT57), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n793_), .A2(new_n799_), .A3(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n343_), .A2(new_n718_), .ZN(new_n804_));
  OAI21_X1  g603(.A(KEYINPUT54), .B1(new_n804_), .B2(new_n661_), .ZN(new_n805_));
  OR3_X1    g604(.A1(new_n804_), .A2(new_n661_), .A3(KEYINPUT54), .ZN(new_n806_));
  AOI22_X1  g605(.A1(new_n803_), .A2(new_n311_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n695_), .A2(new_n531_), .A3(new_n453_), .A4(new_n648_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT119), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n807_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(G113gat), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(new_n359_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n803_), .A2(new_n311_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n806_), .A2(new_n805_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT120), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n809_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT59), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n817_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT120), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n819_), .B1(new_n807_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n811_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n360_), .B1(new_n820_), .B2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n813_), .B1(new_n824_), .B2(new_n812_), .ZN(G1340gat));
  INV_X1    g624(.A(G120gat), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n343_), .B2(KEYINPUT60), .ZN(new_n827_));
  XOR2_X1   g626(.A(new_n827_), .B(KEYINPUT121), .Z(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(KEYINPUT60), .B2(new_n826_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n818_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT122), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n830_), .B(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n343_), .B1(new_n820_), .B2(new_n823_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n832_), .B1(new_n826_), .B2(new_n833_), .ZN(G1341gat));
  INV_X1    g633(.A(KEYINPUT124), .ZN(new_n835_));
  NOR2_X1   g634(.A1(KEYINPUT123), .A2(G127gat), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n311_), .A2(KEYINPUT123), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(G127gat), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n839_), .B1(new_n820_), .B2(new_n823_), .ZN(new_n840_));
  AOI21_X1  g639(.A(G127gat), .B1(new_n811_), .B2(new_n312_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n835_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n822_), .A2(new_n811_), .ZN(new_n843_));
  AOI221_X4 g642(.A(new_n810_), .B1(new_n821_), .B2(new_n819_), .C1(new_n814_), .C2(new_n815_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n838_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n841_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(KEYINPUT124), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n842_), .A2(new_n847_), .ZN(G1342gat));
  INV_X1    g647(.A(G134gat), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n811_), .A2(new_n849_), .A3(new_n626_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n283_), .B1(new_n820_), .B2(new_n823_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n849_), .ZN(G1343gat));
  NOR2_X1   g651(.A1(new_n807_), .A2(new_n648_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n853_), .A2(new_n531_), .A3(new_n654_), .A4(new_n685_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(new_n360_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(new_n366_), .ZN(G1344gat));
  NOR2_X1   g655(.A1(new_n854_), .A2(new_n343_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(new_n367_), .ZN(G1345gat));
  NOR2_X1   g657(.A1(new_n854_), .A2(new_n311_), .ZN(new_n859_));
  XOR2_X1   g658(.A(KEYINPUT61), .B(G155gat), .Z(new_n860_));
  XNOR2_X1  g659(.A(new_n859_), .B(new_n860_), .ZN(G1346gat));
  OAI21_X1  g660(.A(G162gat), .B1(new_n854_), .B2(new_n283_), .ZN(new_n862_));
  OR2_X1    g661(.A1(new_n272_), .A2(G162gat), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n854_), .B2(new_n863_), .ZN(G1347gat));
  NOR2_X1   g663(.A1(new_n807_), .A2(new_n654_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n724_), .A2(new_n535_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(KEYINPUT125), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n865_), .A2(new_n867_), .A3(new_n359_), .ZN(new_n868_));
  OAI21_X1  g667(.A(KEYINPUT62), .B1(new_n868_), .B2(KEYINPUT22), .ZN(new_n869_));
  OAI21_X1  g668(.A(G169gat), .B1(new_n868_), .B2(KEYINPUT62), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n871_), .B1(new_n455_), .B2(new_n869_), .ZN(G1348gat));
  NAND2_X1  g671(.A1(new_n865_), .A2(new_n867_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(G176gat), .B1(new_n874_), .B2(new_n342_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n865_), .B(KEYINPUT126), .ZN(new_n876_));
  AND3_X1   g675(.A1(new_n867_), .A2(G176gat), .A3(new_n342_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n875_), .B1(new_n876_), .B2(new_n877_), .ZN(G1349gat));
  NOR3_X1   g677(.A1(new_n873_), .A2(new_n541_), .A3(new_n311_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n876_), .A2(new_n312_), .A3(new_n867_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n462_), .A2(new_n464_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n879_), .B1(new_n880_), .B2(new_n882_), .ZN(G1350gat));
  OAI21_X1  g682(.A(G190gat), .B1(new_n873_), .B2(new_n283_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n626_), .A2(new_n477_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(KEYINPUT127), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n884_), .B1(new_n873_), .B2(new_n886_), .ZN(G1351gat));
  NOR3_X1   g686(.A1(new_n685_), .A2(new_n531_), .A3(new_n453_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n853_), .A2(new_n888_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n889_), .A2(new_n360_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(new_n405_), .ZN(G1352gat));
  NOR2_X1   g690(.A1(new_n889_), .A2(new_n343_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(G204gat), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n893_), .B1(new_n420_), .B2(new_n892_), .ZN(G1353gat));
  NAND3_X1  g693(.A1(new_n853_), .A2(new_n312_), .A3(new_n888_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n896_));
  AND2_X1   g695(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n895_), .A2(new_n896_), .A3(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n898_), .B1(new_n895_), .B2(new_n896_), .ZN(G1354gat));
  OAI21_X1  g698(.A(G218gat), .B1(new_n889_), .B2(new_n283_), .ZN(new_n900_));
  OR2_X1    g699(.A1(new_n272_), .A2(G218gat), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n889_), .B2(new_n901_), .ZN(G1355gat));
endmodule


