//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n861_, new_n862_, new_n863_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_;
  XOR2_X1   g000(.A(G57gat), .B(G64gat), .Z(new_n202_));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G57gat), .B(G64gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT11), .ZN(new_n206_));
  XOR2_X1   g005(.A(G71gat), .B(G78gat), .Z(new_n207_));
  NAND3_X1  g006(.A1(new_n204_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n206_), .A2(new_n207_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G231gat), .A2(G233gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT80), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n210_), .B(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT78), .B(KEYINPUT79), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G1gat), .B(G8gat), .ZN(new_n215_));
  XOR2_X1   g014(.A(new_n214_), .B(new_n215_), .Z(new_n216_));
  XNOR2_X1  g015(.A(G15gat), .B(G22gat), .ZN(new_n217_));
  INV_X1    g016(.A(G1gat), .ZN(new_n218_));
  INV_X1    g017(.A(G8gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT14), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n217_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n216_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n214_), .B(new_n215_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(new_n221_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n213_), .B(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT16), .B(G183gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(G211gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G127gat), .B(G155gat), .ZN(new_n230_));
  XOR2_X1   g029(.A(new_n229_), .B(new_n230_), .Z(new_n231_));
  INV_X1    g030(.A(KEYINPUT17), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n227_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT81), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n231_), .A2(new_n232_), .ZN(new_n237_));
  OR3_X1    g036(.A1(new_n227_), .A2(new_n233_), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n240_));
  AND3_X1   g039(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n241_));
  AOI21_X1  g040(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n240_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G99gat), .A2(G106gat), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT6), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n246_), .A2(KEYINPUT66), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(G99gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT10), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT10), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(G99gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT64), .B(G106gat), .ZN(new_n254_));
  AOI22_X1  g053(.A1(new_n243_), .A2(new_n248_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  AND2_X1   g054(.A1(G85gat), .A2(G92gat), .ZN(new_n256_));
  NOR2_X1   g055(.A1(G85gat), .A2(G92gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT9), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT65), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT9), .ZN(new_n260_));
  INV_X1    g059(.A(G85gat), .ZN(new_n261_));
  INV_X1    g060(.A(G92gat), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n260_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n258_), .A2(new_n259_), .A3(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n259_), .B1(new_n258_), .B2(new_n263_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n255_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT70), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n255_), .B(new_n268_), .C1(new_n264_), .C2(new_n265_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NOR3_X1   g071(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT68), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT67), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n275_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n246_), .A2(KEYINPUT67), .A3(new_n247_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT7), .ZN(new_n278_));
  INV_X1    g077(.A(G106gat), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(new_n249_), .A3(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT68), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n280_), .A2(new_n281_), .A3(new_n271_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n274_), .A2(new_n276_), .A3(new_n277_), .A4(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n256_), .A2(new_n257_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n283_), .A2(KEYINPUT8), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT8), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n280_), .A2(new_n271_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n287_), .B1(new_n243_), .B2(new_n248_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n284_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n286_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n285_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n270_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(G50gat), .ZN(new_n293_));
  INV_X1    g092(.A(G29gat), .ZN(new_n294_));
  INV_X1    g093(.A(G36gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(G43gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G29gat), .A2(G36gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n297_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n293_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n301_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n303_), .A2(G50gat), .A3(new_n299_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT15), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT15), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n305_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n292_), .A2(new_n310_), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n306_), .A2(new_n285_), .A3(new_n290_), .A4(new_n266_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT75), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G232gat), .A2(G233gat), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n316_), .B(KEYINPUT71), .Z(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT34), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT72), .B(KEYINPUT35), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n318_), .A2(new_n319_), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n311_), .A2(new_n315_), .A3(new_n320_), .A4(new_n321_), .ZN(new_n322_));
  AOI22_X1  g121(.A1(new_n270_), .A2(new_n291_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n319_), .B(new_n318_), .C1(new_n323_), .C2(new_n314_), .ZN(new_n324_));
  XOR2_X1   g123(.A(KEYINPUT74), .B(KEYINPUT36), .Z(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT73), .B(G190gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(G218gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G134gat), .B(G162gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n322_), .A2(new_n324_), .A3(new_n325_), .A4(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT77), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n322_), .A2(new_n324_), .A3(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n329_), .B(KEYINPUT76), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT36), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n332_), .A2(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n331_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n330_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT37), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n322_), .A2(new_n324_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(new_n335_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(KEYINPUT37), .A3(new_n330_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n340_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(G197gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(G204gat), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(G204gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(G197gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT93), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n348_), .A2(KEYINPUT93), .A3(G197gat), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n347_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G211gat), .B(G218gat), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT95), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT21), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  AOI211_X1 g155(.A(new_n353_), .B(new_n356_), .C1(new_n355_), .C2(new_n354_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G183gat), .A2(G190gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT23), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT83), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT23), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(G183gat), .A3(G190gat), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n359_), .A2(KEYINPUT83), .A3(KEYINPUT23), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n362_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(G183gat), .A2(G190gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G169gat), .A2(G176gat), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT22), .B(G169gat), .ZN(new_n372_));
  INV_X1    g171(.A(G176gat), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n371_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n369_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(G169gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n373_), .ZN(new_n377_));
  OR2_X1    g176(.A1(new_n377_), .A2(KEYINPUT24), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n360_), .A2(new_n364_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n377_), .A2(new_n370_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT25), .B(G183gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT26), .B(G190gat), .ZN(new_n383_));
  AOI22_X1  g182(.A1(new_n381_), .A2(KEYINPUT24), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n380_), .A2(new_n384_), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n375_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n354_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT21), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n387_), .B1(new_n353_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT94), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n345_), .A2(G204gat), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT91), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n388_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n346_), .A2(new_n349_), .A3(KEYINPUT91), .ZN(new_n394_));
  AOI21_X1  g193(.A(KEYINPUT92), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n393_), .A2(KEYINPUT92), .A3(new_n394_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n389_), .B(new_n390_), .C1(new_n395_), .C2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n393_), .A2(new_n394_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT92), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n393_), .A2(KEYINPUT92), .A3(new_n394_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n390_), .B1(new_n403_), .B2(new_n389_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n358_), .B(new_n386_), .C1(new_n398_), .C2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n389_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT94), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n357_), .B1(new_n407_), .B2(new_n397_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n366_), .A2(new_n378_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT84), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT84), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n366_), .A2(new_n411_), .A3(new_n378_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n410_), .A2(new_n384_), .A3(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(KEYINPUT22), .B1(new_n376_), .B2(KEYINPUT85), .ZN(new_n414_));
  OR2_X1    g213(.A1(new_n376_), .A2(KEYINPUT22), .ZN(new_n415_));
  OAI211_X1 g214(.A(new_n373_), .B(new_n414_), .C1(new_n415_), .C2(KEYINPUT85), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n379_), .A2(new_n368_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(new_n417_), .A3(new_n370_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n413_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n405_), .B(KEYINPUT20), .C1(new_n408_), .C2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G226gat), .A2(G233gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT19), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT99), .B1(new_n421_), .B2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n358_), .B1(new_n398_), .B2(new_n404_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT20), .B1(new_n425_), .B2(new_n419_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n408_), .A2(new_n386_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n423_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT20), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n429_), .B1(new_n408_), .B2(new_n386_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT99), .ZN(new_n431_));
  INV_X1    g230(.A(new_n423_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n425_), .A2(new_n419_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .A4(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n424_), .A2(new_n428_), .A3(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT18), .B(G64gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(G92gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G8gat), .B(G36gat), .ZN(new_n438_));
  XOR2_X1   g237(.A(new_n437_), .B(new_n438_), .Z(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n435_), .A2(new_n440_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n424_), .A2(new_n439_), .A3(new_n428_), .A4(new_n434_), .ZN(new_n442_));
  AOI21_X1  g241(.A(KEYINPUT27), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT27), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n405_), .A2(KEYINPUT20), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n407_), .A2(new_n397_), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n446_), .A2(new_n358_), .B1(new_n418_), .B2(new_n413_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n423_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n429_), .B1(new_n408_), .B2(new_n420_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n386_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n425_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(new_n432_), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n448_), .A2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n444_), .B1(new_n453_), .B2(new_n440_), .ZN(new_n454_));
  AND3_X1   g253(.A1(new_n454_), .A2(KEYINPUT102), .A3(new_n442_), .ZN(new_n455_));
  AOI21_X1  g254(.A(KEYINPUT102), .B1(new_n454_), .B2(new_n442_), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n443_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G225gat), .A2(G233gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G127gat), .B(G134gat), .ZN(new_n459_));
  INV_X1    g258(.A(G113gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(G120gat), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT3), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT88), .ZN(new_n464_));
  NOR2_X1   g263(.A1(G141gat), .A2(G148gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G141gat), .A2(G148gat), .ZN(new_n467_));
  AND2_X1   g266(.A1(KEYINPUT89), .A2(KEYINPUT2), .ZN(new_n468_));
  NOR2_X1   g267(.A1(KEYINPUT89), .A2(KEYINPUT2), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n467_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n466_), .B(new_n470_), .C1(new_n467_), .C2(new_n469_), .ZN(new_n471_));
  AND2_X1   g270(.A1(G155gat), .A2(G162gat), .ZN(new_n472_));
  NOR2_X1   g271(.A1(G155gat), .A2(G162gat), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n471_), .A2(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n465_), .B1(new_n472_), .B2(KEYINPUT1), .ZN(new_n476_));
  INV_X1    g275(.A(new_n474_), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n476_), .B(new_n467_), .C1(KEYINPUT1), .C2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n475_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT100), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n462_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(G120gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n461_), .B(new_n482_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n483_), .A2(KEYINPUT100), .A3(new_n475_), .A4(new_n478_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n481_), .A2(new_n484_), .A3(KEYINPUT4), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT4), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n479_), .A2(new_n462_), .A3(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n458_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT0), .B(G57gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(G85gat), .ZN(new_n491_));
  XOR2_X1   g290(.A(G1gat), .B(G29gat), .Z(new_n492_));
  XOR2_X1   g291(.A(new_n491_), .B(new_n492_), .Z(new_n493_));
  INV_X1    g292(.A(new_n458_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n494_), .B1(new_n481_), .B2(new_n484_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n489_), .A2(new_n493_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT101), .ZN(new_n498_));
  INV_X1    g297(.A(new_n493_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n499_), .B1(new_n488_), .B2(new_n495_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n497_), .A2(new_n498_), .A3(new_n500_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n489_), .A2(KEYINPUT101), .A3(new_n493_), .A4(new_n496_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT86), .B(KEYINPUT87), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G71gat), .B(G99gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT30), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n413_), .A2(new_n508_), .A3(new_n418_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n508_), .B1(new_n413_), .B2(new_n418_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n462_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n419_), .A2(KEYINPUT30), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n513_), .A2(new_n483_), .A3(new_n509_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G15gat), .B(G43gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT31), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G227gat), .A2(G233gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n512_), .A2(new_n514_), .A3(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n518_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n507_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n518_), .ZN(new_n522_));
  NOR3_X1   g321(.A1(new_n510_), .A2(new_n511_), .A3(new_n462_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n483_), .B1(new_n513_), .B2(new_n509_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n522_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n512_), .A2(new_n514_), .A3(new_n518_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n525_), .A2(new_n506_), .A3(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n521_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT98), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n479_), .A2(KEYINPUT29), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G22gat), .B(G50gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT28), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n531_), .B(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(G78gat), .B(G106gat), .Z(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G228gat), .A2(G233gat), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n538_), .B(KEYINPUT90), .Z(new_n539_));
  NAND2_X1  g338(.A1(new_n479_), .A2(KEYINPUT29), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n425_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(KEYINPUT96), .B(KEYINPUT29), .Z(new_n542_));
  NAND2_X1  g341(.A1(new_n479_), .A2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n539_), .B1(new_n425_), .B2(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n537_), .B1(new_n541_), .B2(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n535_), .B1(new_n545_), .B2(KEYINPUT97), .ZN(new_n546_));
  INV_X1    g345(.A(new_n539_), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n479_), .A2(new_n542_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n547_), .B1(new_n408_), .B2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n425_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(new_n536_), .A3(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n536_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT97), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n551_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n530_), .B1(new_n546_), .B2(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n534_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n545_), .A2(KEYINPUT97), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n556_), .A2(new_n557_), .A3(KEYINPUT98), .A4(new_n551_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n555_), .A2(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n535_), .B1(new_n545_), .B2(new_n551_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n529_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n562_));
  AOI211_X1 g361(.A(new_n560_), .B(new_n528_), .C1(new_n555_), .C2(new_n558_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n457_), .B(new_n503_), .C1(new_n562_), .C2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n500_), .B(KEYINPUT33), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n485_), .A2(new_n458_), .A3(new_n487_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n481_), .A2(new_n484_), .A3(new_n494_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(new_n493_), .A3(new_n567_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n565_), .A2(new_n442_), .A3(new_n441_), .A4(new_n568_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n439_), .A2(KEYINPUT32), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n435_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n453_), .A2(new_n570_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n571_), .A2(new_n502_), .A3(new_n501_), .A4(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n569_), .A2(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n560_), .B1(new_n555_), .B2(new_n558_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n574_), .A2(new_n575_), .A3(new_n528_), .ZN(new_n576_));
  AOI211_X1 g375(.A(new_n239_), .B(new_n344_), .C1(new_n564_), .C2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G120gat), .B(G148gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(new_n348_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT5), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(new_n373_), .ZN(new_n581_));
  AND4_X1   g380(.A1(new_n210_), .A2(new_n285_), .A3(new_n290_), .A4(new_n266_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n208_), .A2(new_n209_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT12), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n582_), .B1(new_n292_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G230gat), .A2(G233gat), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n285_), .A2(new_n290_), .A3(new_n266_), .ZN(new_n588_));
  AOI21_X1  g387(.A(KEYINPUT12), .B1(new_n588_), .B2(new_n583_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n586_), .A2(new_n587_), .A3(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n291_), .A2(new_n210_), .A3(new_n266_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT69), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n588_), .A2(new_n583_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n592_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n587_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n588_), .A2(KEYINPUT69), .A3(new_n583_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n595_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n581_), .B1(new_n591_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n591_), .A2(new_n598_), .A3(new_n581_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n602_), .A2(KEYINPUT13), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(KEYINPUT13), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n226_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(new_n306_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(G229gat), .A2(G233gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n305_), .B(KEYINPUT15), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n608_), .B(new_n609_), .C1(new_n607_), .C2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n609_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n226_), .A2(new_n305_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n306_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n612_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n611_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G113gat), .B(G141gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(new_n376_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(new_n345_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n616_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n619_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n611_), .A2(new_n615_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(KEYINPUT82), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT82), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n623_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n606_), .A2(new_n628_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n577_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n503_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n630_), .A2(new_n218_), .A3(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n338_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n564_), .B2(new_n576_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n239_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n606_), .A2(new_n624_), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n636_), .A2(new_n637_), .A3(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n218_), .B1(new_n639_), .B2(new_n631_), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n634_), .A2(new_n640_), .ZN(G1324gat));
  INV_X1    g440(.A(new_n457_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n630_), .A2(new_n219_), .A3(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n639_), .A2(new_n642_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(G8gat), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n645_), .A2(KEYINPUT39), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(KEYINPUT39), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n643_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g448(.A(G15gat), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n650_), .B1(new_n639_), .B2(new_n529_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT41), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n630_), .A2(new_n650_), .A3(new_n529_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1326gat));
  INV_X1    g453(.A(G22gat), .ZN(new_n655_));
  INV_X1    g454(.A(new_n575_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n630_), .A2(new_n655_), .A3(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n639_), .A2(new_n656_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(G22gat), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n659_), .A2(KEYINPUT42), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(KEYINPUT42), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n657_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT104), .Z(G1327gat));
  NOR3_X1   g462(.A1(new_n606_), .A2(new_n637_), .A3(new_n624_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT43), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n564_), .A2(new_n576_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n666_), .B2(new_n344_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n344_), .ZN(new_n668_));
  AOI211_X1 g467(.A(KEYINPUT43), .B(new_n668_), .C1(new_n564_), .C2(new_n576_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n664_), .B1(new_n667_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  OAI211_X1 g471(.A(KEYINPUT44), .B(new_n664_), .C1(new_n667_), .C2(new_n669_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n672_), .A2(new_n631_), .A3(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n338_), .B1(new_n564_), .B2(new_n576_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n675_), .A2(new_n239_), .A3(new_n629_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n503_), .A2(G29gat), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT105), .ZN(new_n678_));
  OAI22_X1  g477(.A1(new_n674_), .A2(new_n294_), .B1(new_n676_), .B2(new_n678_), .ZN(G1328gat));
  NAND3_X1  g478(.A1(new_n672_), .A2(new_n642_), .A3(new_n673_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT106), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n672_), .A2(new_n682_), .A3(new_n642_), .A4(new_n673_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n681_), .A2(G36gat), .A3(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n676_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n685_), .A2(new_n295_), .A3(new_n642_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT45), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n684_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT46), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n684_), .A2(KEYINPUT46), .A3(new_n687_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1329gat));
  NAND4_X1  g491(.A1(new_n672_), .A2(G43gat), .A3(new_n529_), .A4(new_n673_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n297_), .B1(new_n676_), .B2(new_n528_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(KEYINPUT107), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n693_), .A2(new_n697_), .A3(new_n694_), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n696_), .A2(KEYINPUT47), .A3(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(KEYINPUT47), .B1(new_n696_), .B2(new_n698_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1330gat));
  NAND3_X1  g500(.A1(new_n672_), .A2(new_n656_), .A3(new_n673_), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n702_), .A2(KEYINPUT108), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(KEYINPUT108), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n703_), .A2(G50gat), .A3(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n685_), .A2(new_n293_), .A3(new_n656_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1331gat));
  AOI21_X1  g506(.A(new_n239_), .B1(new_n625_), .B2(new_n627_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n636_), .A2(new_n606_), .A3(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(G57gat), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n709_), .A2(new_n710_), .A3(new_n503_), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n577_), .A2(new_n624_), .A3(new_n606_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n631_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n711_), .B1(new_n713_), .B2(new_n710_), .ZN(G1332gat));
  OAI21_X1  g513(.A(G64gat), .B1(new_n709_), .B2(new_n457_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT48), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n457_), .A2(G64gat), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT109), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n712_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n716_), .A2(new_n719_), .ZN(G1333gat));
  OAI21_X1  g519(.A(G71gat), .B1(new_n709_), .B2(new_n528_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT49), .ZN(new_n722_));
  INV_X1    g521(.A(G71gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n712_), .A2(new_n723_), .A3(new_n529_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(G1334gat));
  OAI21_X1  g524(.A(G78gat), .B1(new_n709_), .B2(new_n575_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT50), .ZN(new_n727_));
  INV_X1    g526(.A(G78gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n712_), .A2(new_n728_), .A3(new_n656_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1335gat));
  NOR3_X1   g529(.A1(new_n605_), .A2(new_n637_), .A3(new_n623_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n675_), .A2(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(G85gat), .B1(new_n732_), .B2(new_n631_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT110), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n667_), .A2(new_n669_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(new_n731_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n503_), .A2(new_n261_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(G1336gat));
  AOI21_X1  g538(.A(G92gat), .B1(new_n732_), .B2(new_n642_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n457_), .A2(new_n262_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n737_), .B2(new_n741_), .ZN(G1337gat));
  OAI21_X1  g541(.A(G99gat), .B1(new_n736_), .B2(new_n528_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n732_), .A2(new_n253_), .A3(new_n529_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g545(.A(G106gat), .B1(new_n736_), .B2(new_n575_), .ZN(new_n747_));
  XOR2_X1   g546(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n732_), .A2(new_n254_), .A3(new_n656_), .ZN(new_n751_));
  OAI211_X1 g550(.A(G106gat), .B(new_n748_), .C1(new_n736_), .C2(new_n575_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n750_), .A2(new_n751_), .A3(new_n752_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g553(.A(KEYINPUT112), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n605_), .A2(new_n708_), .A3(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n605_), .B2(new_n708_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n668_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT54), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n608_), .B(new_n612_), .C1(new_n607_), .C2(new_n610_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n609_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(new_n761_), .A3(new_n619_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n622_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n601_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n581_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n584_), .B1(new_n270_), .B2(new_n291_), .ZN(new_n766_));
  NOR4_X1   g565(.A1(new_n766_), .A2(new_n589_), .A3(new_n596_), .A4(new_n582_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n285_), .A2(new_n290_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n768_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n592_), .B1(new_n769_), .B2(new_n584_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n596_), .B1(new_n770_), .B2(new_n589_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n767_), .B1(new_n771_), .B2(KEYINPUT55), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n773_));
  NOR4_X1   g572(.A1(new_n770_), .A2(new_n773_), .A3(new_n596_), .A4(new_n589_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n765_), .B1(new_n772_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT56), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  OAI211_X1 g576(.A(KEYINPUT56), .B(new_n765_), .C1(new_n772_), .C2(new_n774_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n764_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n344_), .B1(new_n779_), .B2(KEYINPUT58), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT114), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n779_), .A2(KEYINPUT58), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n344_), .B(KEYINPUT114), .C1(new_n779_), .C2(KEYINPUT58), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n782_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n602_), .A2(new_n763_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT113), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n788_));
  INV_X1    g587(.A(new_n601_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n763_), .B(new_n788_), .C1(new_n789_), .C2(new_n599_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n787_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n623_), .A2(new_n601_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n792_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n338_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT57), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n777_), .A2(new_n778_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n792_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n788_), .B1(new_n602_), .B2(new_n763_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n790_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n799_), .A2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n803_), .A2(KEYINPUT57), .A3(new_n338_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n796_), .A2(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n239_), .B1(new_n785_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n759_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT59), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n457_), .A2(new_n631_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n563_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n807_), .A2(new_n808_), .A3(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT115), .B1(new_n785_), .B2(new_n805_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n782_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n815_), .A2(new_n816_), .A3(new_n796_), .A4(new_n804_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n814_), .A2(new_n239_), .A3(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n811_), .B1(new_n818_), .B2(new_n759_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n813_), .B1(new_n819_), .B2(new_n808_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  OAI211_X1 g621(.A(KEYINPUT116), .B(new_n813_), .C1(new_n819_), .C2(new_n808_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n628_), .A2(new_n460_), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n822_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(G113gat), .B1(new_n819_), .B2(new_n623_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(G1340gat));
  OAI21_X1  g626(.A(G120gat), .B1(new_n820_), .B2(new_n605_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n482_), .B1(new_n605_), .B2(KEYINPUT60), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n819_), .B(new_n829_), .C1(KEYINPUT60), .C2(new_n482_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(G1341gat));
  XNOR2_X1  g630(.A(KEYINPUT118), .B(G127gat), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n822_), .A2(new_n637_), .A3(new_n823_), .A4(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n818_), .A2(new_n759_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n834_), .A2(new_n637_), .A3(new_n812_), .ZN(new_n835_));
  INV_X1    g634(.A(G127gat), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n835_), .A2(KEYINPUT117), .A3(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(KEYINPUT117), .B1(new_n835_), .B2(new_n836_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n833_), .A2(new_n839_), .ZN(G1342gat));
  XOR2_X1   g639(.A(KEYINPUT119), .B(G134gat), .Z(new_n841_));
  NAND4_X1  g640(.A1(new_n822_), .A2(new_n344_), .A3(new_n823_), .A4(new_n841_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n819_), .A2(new_n635_), .ZN(new_n843_));
  OR2_X1    g642(.A1(new_n843_), .A2(G134gat), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n842_), .A2(new_n844_), .ZN(G1343gat));
  INV_X1    g644(.A(new_n562_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n846_), .B1(new_n818_), .B2(new_n759_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT120), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(new_n848_), .A3(new_n810_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n848_), .B1(new_n847_), .B2(new_n810_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n623_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(G141gat), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n834_), .A2(new_n562_), .A3(new_n810_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(KEYINPUT120), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n849_), .ZN(new_n856_));
  INV_X1    g655(.A(G141gat), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n856_), .A2(new_n857_), .A3(new_n623_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n853_), .A2(new_n858_), .ZN(G1344gat));
  OAI21_X1  g658(.A(new_n606_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(G148gat), .ZN(new_n861_));
  INV_X1    g660(.A(G148gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n856_), .A2(new_n862_), .A3(new_n606_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n863_), .ZN(G1345gat));
  XNOR2_X1  g663(.A(KEYINPUT61), .B(G155gat), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n865_), .B1(new_n856_), .B2(new_n637_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n865_), .ZN(new_n867_));
  AOI211_X1 g666(.A(new_n239_), .B(new_n867_), .C1(new_n855_), .C2(new_n849_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n866_), .A2(new_n868_), .ZN(G1346gat));
  AOI21_X1  g668(.A(G162gat), .B1(new_n856_), .B2(new_n635_), .ZN(new_n870_));
  INV_X1    g669(.A(G162gat), .ZN(new_n871_));
  AOI211_X1 g670(.A(new_n871_), .B(new_n668_), .C1(new_n855_), .C2(new_n849_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n870_), .A2(new_n872_), .ZN(G1347gat));
  AOI21_X1  g672(.A(new_n656_), .B1(new_n759_), .B2(new_n806_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n642_), .A2(new_n503_), .A3(new_n529_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(KEYINPUT121), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(G169gat), .B1(new_n877_), .B2(new_n624_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT62), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n874_), .A2(new_n372_), .A3(new_n623_), .A4(new_n876_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n878_), .A2(new_n879_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n880_), .A2(new_n881_), .A3(new_n882_), .ZN(G1348gat));
  AOI21_X1  g682(.A(new_n656_), .B1(new_n818_), .B2(new_n759_), .ZN(new_n884_));
  AND4_X1   g683(.A1(G176gat), .A2(new_n884_), .A3(new_n606_), .A4(new_n876_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n373_), .B1(new_n877_), .B2(new_n605_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n887_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n885_), .B1(new_n888_), .B2(new_n889_), .ZN(G1349gat));
  INV_X1    g689(.A(new_n382_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n876_), .A2(new_n637_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n874_), .A2(new_n891_), .A3(new_n893_), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n894_), .B(KEYINPUT123), .Z(new_n895_));
  AOI21_X1  g694(.A(G183gat), .B1(new_n884_), .B2(new_n893_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n895_), .A2(new_n896_), .ZN(G1350gat));
  OAI21_X1  g696(.A(G190gat), .B1(new_n877_), .B2(new_n668_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n635_), .A2(new_n383_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n877_), .B2(new_n899_), .ZN(G1351gat));
  NOR3_X1   g699(.A1(new_n846_), .A2(KEYINPUT124), .A3(new_n631_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n901_), .A2(new_n457_), .ZN(new_n902_));
  OAI21_X1  g701(.A(KEYINPUT124), .B1(new_n846_), .B2(new_n631_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n834_), .A2(new_n623_), .A3(new_n902_), .A4(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n345_), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n905_), .A2(KEYINPUT126), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(KEYINPUT126), .ZN(new_n907_));
  OR3_X1    g706(.A1(new_n904_), .A2(KEYINPUT125), .A3(new_n345_), .ZN(new_n908_));
  OAI21_X1  g707(.A(KEYINPUT125), .B1(new_n904_), .B2(new_n345_), .ZN(new_n909_));
  AOI22_X1  g708(.A1(new_n906_), .A2(new_n907_), .B1(new_n908_), .B2(new_n909_), .ZN(G1352gat));
  AND3_X1   g709(.A1(new_n834_), .A2(new_n902_), .A3(new_n903_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n606_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G204gat), .ZN(G1353gat));
  XOR2_X1   g712(.A(KEYINPUT63), .B(G211gat), .Z(new_n914_));
  AND3_X1   g713(.A1(new_n911_), .A2(new_n637_), .A3(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n911_), .A2(new_n637_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n915_), .B1(new_n916_), .B2(new_n917_), .ZN(G1354gat));
  NAND2_X1  g717(.A1(new_n911_), .A2(new_n635_), .ZN(new_n919_));
  XOR2_X1   g718(.A(KEYINPUT127), .B(G218gat), .Z(new_n920_));
  NOR2_X1   g719(.A1(new_n668_), .A2(new_n920_), .ZN(new_n921_));
  AOI22_X1  g720(.A1(new_n919_), .A2(new_n920_), .B1(new_n911_), .B2(new_n921_), .ZN(G1355gat));
endmodule


