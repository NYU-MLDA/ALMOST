//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 1 0 0 0 0 1 1 0 1 1 0 1 0 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n607_, new_n608_, new_n609_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n814_, new_n816_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n844_,
    new_n846_, new_n847_, new_n848_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT95), .B(KEYINPUT27), .Z(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G197gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G204gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT85), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G204gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G197gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n205_), .A2(KEYINPUT85), .A3(G204gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n208_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n212_), .A2(KEYINPUT21), .ZN(new_n213_));
  XOR2_X1   g012(.A(G211gat), .B(G218gat), .Z(new_n214_));
  NAND2_X1  g013(.A1(new_n206_), .A2(new_n210_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n214_), .B1(KEYINPUT21), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  AND2_X1   g016(.A1(new_n214_), .A2(KEYINPUT21), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(new_n212_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(KEYINPUT23), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT79), .B(G183gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n222_), .B1(G190gat), .B2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(G169gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  OR2_X1    g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(KEYINPUT24), .A3(new_n229_), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n222_), .B(new_n230_), .C1(KEYINPUT24), .C2(new_n228_), .ZN(new_n231_));
  XOR2_X1   g030(.A(KEYINPUT26), .B(G190gat), .Z(new_n232_));
  NAND2_X1  g031(.A1(new_n223_), .A2(KEYINPUT25), .ZN(new_n233_));
  OR2_X1    g032(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n232_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n227_), .B1(new_n231_), .B2(new_n235_), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n220_), .A2(new_n236_), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n217_), .A2(new_n219_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n222_), .B1(KEYINPUT24), .B2(new_n228_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT25), .B(G183gat), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n230_), .B1(new_n241_), .B2(new_n232_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n239_), .B1(KEYINPUT87), .B2(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n242_), .A2(KEYINPUT87), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n222_), .B1(G183gat), .B2(G190gat), .ZN(new_n245_));
  AOI22_X1  g044(.A1(new_n243_), .A2(new_n244_), .B1(new_n226_), .B2(new_n245_), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n237_), .B(KEYINPUT20), .C1(new_n238_), .C2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G226gat), .A2(G233gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT19), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n220_), .A2(new_n236_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT88), .ZN(new_n252_));
  INV_X1    g051(.A(new_n249_), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n253_), .A2(KEYINPUT20), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n246_), .A2(new_n238_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT89), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n246_), .A2(KEYINPUT89), .A3(new_n238_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n250_), .B1(new_n255_), .B2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G8gat), .B(G36gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT18), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G64gat), .B(G92gat), .ZN(new_n264_));
  XOR2_X1   g063(.A(new_n263_), .B(new_n264_), .Z(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  AND2_X1   g065(.A1(new_n261_), .A2(new_n266_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n250_), .B(new_n265_), .C1(new_n255_), .C2(new_n260_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n204_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n256_), .A2(KEYINPUT20), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n253_), .B1(new_n252_), .B2(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n247_), .A2(new_n249_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n268_), .B(KEYINPUT27), .C1(new_n274_), .C2(new_n265_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n270_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT97), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT97), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n270_), .A2(new_n278_), .A3(new_n275_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G141gat), .A2(G148gat), .ZN(new_n282_));
  INV_X1    g081(.A(G141gat), .ZN(new_n283_));
  INV_X1    g082(.A(G148gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G155gat), .A2(G162gat), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT84), .B1(new_n286_), .B2(KEYINPUT1), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(KEYINPUT1), .ZN(new_n288_));
  OR2_X1    g087(.A1(G155gat), .A2(G162gat), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n287_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  NOR3_X1   g089(.A1(new_n286_), .A2(KEYINPUT84), .A3(KEYINPUT1), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n282_), .B(new_n285_), .C1(new_n290_), .C2(new_n291_), .ZN(new_n292_));
  OR3_X1    g091(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT2), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n282_), .A2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n293_), .A2(new_n295_), .A3(new_n296_), .A4(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(new_n286_), .A3(new_n289_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n292_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT29), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT28), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G22gat), .B(G50gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G228gat), .A2(G233gat), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n220_), .B(new_n306_), .C1(new_n301_), .C2(new_n300_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n292_), .A2(new_n299_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT86), .B(KEYINPUT29), .ZN(new_n309_));
  AOI22_X1  g108(.A1(new_n217_), .A2(new_n219_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n307_), .B1(new_n310_), .B2(new_n306_), .ZN(new_n311_));
  XOR2_X1   g110(.A(G78gat), .B(G106gat), .Z(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n305_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n305_), .A2(new_n313_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G127gat), .B(G134gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT83), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G113gat), .B(G120gat), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n317_), .A2(KEYINPUT83), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n317_), .A2(KEYINPUT83), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n322_), .A2(new_n323_), .A3(new_n319_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n321_), .A2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(new_n300_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT4), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G225gat), .A2(G233gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT4), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n325_), .A2(new_n330_), .A3(new_n308_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n327_), .A2(KEYINPUT90), .A3(new_n329_), .A4(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n326_), .A2(new_n328_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n327_), .A2(new_n329_), .A3(new_n331_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT90), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n334_), .A2(new_n337_), .ZN(new_n338_));
  XOR2_X1   g137(.A(G1gat), .B(G29gat), .Z(new_n339_));
  XNOR2_X1  g138(.A(G57gat), .B(G85gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT91), .B(KEYINPUT0), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n338_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n343_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n334_), .A2(new_n345_), .A3(new_n337_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G227gat), .A2(G233gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(G15gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT81), .B(G43gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  XOR2_X1   g151(.A(G71gat), .B(G99gat), .Z(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(KEYINPUT80), .B(KEYINPUT30), .Z(new_n355_));
  XNOR2_X1  g154(.A(new_n236_), .B(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n354_), .B1(new_n356_), .B2(KEYINPUT82), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(KEYINPUT82), .ZN(new_n358_));
  XOR2_X1   g157(.A(new_n357_), .B(new_n358_), .Z(new_n359_));
  XOR2_X1   g158(.A(new_n325_), .B(KEYINPUT31), .Z(new_n360_));
  XOR2_X1   g159(.A(new_n359_), .B(new_n360_), .Z(new_n361_));
  NAND2_X1  g160(.A1(new_n348_), .A2(new_n361_), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n281_), .A2(new_n316_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n316_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n265_), .A2(KEYINPUT32), .ZN(new_n365_));
  MUX2_X1   g164(.A(new_n274_), .B(new_n261_), .S(new_n365_), .Z(new_n366_));
  NAND2_X1  g165(.A1(new_n347_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT94), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT94), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n347_), .A2(new_n369_), .A3(new_n366_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n267_), .A2(new_n269_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n327_), .A2(new_n328_), .A3(new_n331_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n345_), .B1(new_n326_), .B2(new_n329_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT93), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT33), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n372_), .B(new_n376_), .C1(new_n377_), .C2(new_n346_), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n346_), .A2(KEYINPUT92), .A3(new_n377_), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT92), .B1(new_n346_), .B2(new_n377_), .ZN(new_n380_));
  NOR3_X1   g179(.A1(new_n378_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n364_), .B1(new_n371_), .B2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n316_), .A2(new_n344_), .A3(new_n346_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n276_), .A2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT96), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n382_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n361_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n363_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G1gat), .B(G8gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT74), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G15gat), .B(G22gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G1gat), .A2(G8gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT14), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  OR2_X1    g193(.A1(new_n390_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n390_), .A2(new_n394_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G29gat), .B(G36gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G43gat), .B(G50gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n397_), .B(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G229gat), .A2(G233gat), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n400_), .B(KEYINPUT15), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n405_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n397_), .A2(new_n400_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(new_n407_), .A3(new_n402_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n404_), .A2(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(new_n409_), .B(KEYINPUT77), .Z(new_n410_));
  XNOR2_X1  g209(.A(G113gat), .B(G141gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G169gat), .B(G197gat), .ZN(new_n412_));
  XOR2_X1   g211(.A(new_n411_), .B(new_n412_), .Z(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n414_), .A2(KEYINPUT76), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n410_), .B(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT78), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n388_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G85gat), .A2(G92gat), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(G85gat), .A2(G92gat), .ZN(new_n422_));
  INV_X1    g221(.A(G92gat), .ZN(new_n423_));
  OAI22_X1  g222(.A1(new_n421_), .A2(new_n422_), .B1(KEYINPUT9), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n422_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT9), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n426_), .A3(new_n420_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT64), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n424_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  AND2_X1   g228(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n430_));
  NOR2_X1   g229(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(G106gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G99gat), .A2(G106gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT6), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT6), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(G99gat), .A3(G106gat), .ZN(new_n437_));
  AOI22_X1  g236(.A1(new_n432_), .A2(new_n433_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n429_), .A2(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n428_), .B1(new_n424_), .B2(new_n427_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(G99gat), .A2(G106gat), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT7), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT65), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT65), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n445_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  AOI22_X1  g246(.A1(new_n435_), .A2(new_n437_), .B1(new_n443_), .B2(new_n442_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n421_), .A2(new_n422_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT8), .ZN(new_n452_));
  AOI22_X1  g251(.A1(new_n439_), .A2(new_n441_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n451_), .A2(new_n452_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n405_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G232gat), .A2(G233gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT35), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n429_), .A2(new_n438_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n425_), .A2(new_n420_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n464_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n465_));
  OAI22_X1  g264(.A1(new_n463_), .A2(new_n440_), .B1(new_n465_), .B2(KEYINPUT8), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n466_), .A2(new_n454_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(new_n400_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n457_), .A2(new_n462_), .A3(new_n468_), .ZN(new_n469_));
  OR2_X1    g268(.A1(new_n460_), .A2(new_n461_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT73), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G190gat), .B(G218gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G134gat), .B(G162gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n476_), .A2(KEYINPUT36), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n473_), .A2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n471_), .A2(new_n472_), .A3(new_n477_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n471_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n482_), .A2(KEYINPUT36), .A3(new_n476_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n484_), .A2(KEYINPUT37), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(KEYINPUT37), .ZN(new_n486_));
  OR2_X1    g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT68), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT67), .ZN(new_n489_));
  INV_X1    g288(.A(G57gat), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n490_), .A2(G64gat), .ZN(new_n491_));
  INV_X1    g290(.A(G64gat), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n492_), .A2(G57gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT66), .B1(new_n491_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(G57gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n490_), .A2(G64gat), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT66), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n494_), .A2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n489_), .B1(new_n499_), .B2(KEYINPUT11), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT11), .ZN(new_n501_));
  AOI211_X1 g300(.A(KEYINPUT67), .B(new_n501_), .C1(new_n494_), .C2(new_n498_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n494_), .A2(new_n501_), .A3(new_n498_), .ZN(new_n503_));
  XOR2_X1   g302(.A(G71gat), .B(G78gat), .Z(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NOR3_X1   g304(.A1(new_n500_), .A2(new_n502_), .A3(new_n505_), .ZN(new_n506_));
  AND3_X1   g305(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n497_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT11), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT67), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n499_), .A2(new_n489_), .A3(KEYINPUT11), .ZN(new_n511_));
  AOI22_X1  g310(.A1(new_n510_), .A2(new_n511_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n488_), .B1(new_n506_), .B2(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n505_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n510_), .A2(new_n511_), .A3(new_n503_), .A4(new_n504_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(new_n515_), .A3(KEYINPUT68), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n513_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(new_n467_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n513_), .A2(new_n456_), .A3(new_n516_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(KEYINPUT69), .A3(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G230gat), .A2(G233gat), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n520_), .B(new_n522_), .C1(KEYINPUT69), .C2(new_n518_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n522_), .B1(new_n517_), .B2(new_n467_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT12), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n519_), .A2(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n506_), .A2(new_n512_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT70), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n527_), .A2(new_n528_), .A3(new_n456_), .A4(KEYINPUT12), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT12), .B1(new_n466_), .B2(new_n454_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n514_), .A2(new_n515_), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT70), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n524_), .A2(new_n526_), .A3(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(G120gat), .B(G148gat), .Z(new_n535_));
  XNOR2_X1  g334(.A(G176gat), .B(G204gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n523_), .A2(new_n534_), .A3(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n539_), .B1(new_n523_), .B2(new_n534_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n543_), .A2(KEYINPUT13), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(KEYINPUT13), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G231gat), .A2(G233gat), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n397_), .B(new_n547_), .Z(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(new_n531_), .ZN(new_n549_));
  XOR2_X1   g348(.A(KEYINPUT75), .B(KEYINPUT17), .Z(new_n550_));
  XNOR2_X1  g349(.A(G127gat), .B(G155gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT16), .ZN(new_n552_));
  XOR2_X1   g351(.A(G183gat), .B(G211gat), .Z(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  OR3_X1    g353(.A1(new_n549_), .A2(new_n550_), .A3(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n554_), .B(KEYINPUT17), .Z(new_n556_));
  INV_X1    g355(.A(new_n517_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n556_), .B1(new_n557_), .B2(new_n548_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n558_), .B1(new_n548_), .B2(new_n557_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n555_), .A2(new_n559_), .ZN(new_n560_));
  NOR3_X1   g359(.A1(new_n487_), .A2(new_n546_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n419_), .A2(new_n561_), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n348_), .A2(G1gat), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n202_), .B1(new_n564_), .B2(KEYINPUT38), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT38), .ZN(new_n566_));
  NOR4_X1   g365(.A1(new_n562_), .A2(KEYINPUT98), .A3(new_n566_), .A4(new_n563_), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n566_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT100), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n388_), .A2(new_n484_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n416_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n546_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n560_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT99), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n571_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(G1gat), .B1(new_n578_), .B2(new_n348_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n568_), .A2(new_n570_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT101), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n568_), .A2(new_n570_), .A3(KEYINPUT101), .A4(new_n579_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(G1324gat));
  XNOR2_X1  g383(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n577_), .A2(new_n281_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(G8gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT39), .ZN(new_n588_));
  OR3_X1    g387(.A1(new_n562_), .A2(G8gat), .A3(new_n280_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n585_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n587_), .A2(KEYINPUT39), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT39), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n592_), .B1(new_n586_), .B2(G8gat), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n589_), .B(new_n585_), .C1(new_n591_), .C2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n590_), .A2(new_n595_), .ZN(G1325gat));
  NAND2_X1  g395(.A1(new_n577_), .A2(new_n361_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(G15gat), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n598_), .A2(KEYINPUT103), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(KEYINPUT103), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT41), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  OR3_X1    g402(.A1(new_n562_), .A2(G15gat), .A3(new_n387_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n599_), .A2(KEYINPUT41), .A3(new_n600_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n603_), .A2(new_n604_), .A3(new_n605_), .ZN(G1326gat));
  OAI21_X1  g405(.A(G22gat), .B1(new_n578_), .B2(new_n364_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT42), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n364_), .A2(G22gat), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n608_), .B1(new_n562_), .B2(new_n609_), .ZN(G1327gat));
  INV_X1    g409(.A(new_n484_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n546_), .A2(new_n611_), .A3(new_n574_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n419_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(G29gat), .B1(new_n614_), .B2(new_n347_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n485_), .A2(new_n486_), .ZN(new_n616_));
  OAI21_X1  g415(.A(KEYINPUT43), .B1(new_n388_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT43), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n361_), .B1(new_n382_), .B2(new_n385_), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n618_), .B(new_n487_), .C1(new_n619_), .C2(new_n363_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n617_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n573_), .A2(new_n560_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT44), .B1(new_n621_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT44), .ZN(new_n625_));
  AOI211_X1 g424(.A(new_n625_), .B(new_n622_), .C1(new_n617_), .C2(new_n620_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n347_), .A2(G29gat), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n615_), .B1(new_n627_), .B2(new_n628_), .ZN(G1328gat));
  NAND2_X1  g428(.A1(new_n621_), .A2(new_n623_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(new_n625_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n621_), .A2(KEYINPUT44), .A3(new_n623_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n631_), .A2(new_n281_), .A3(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(G36gat), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n280_), .A2(G36gat), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  OR3_X1    g435(.A1(new_n613_), .A2(KEYINPUT45), .A3(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(KEYINPUT45), .B1(new_n613_), .B2(new_n636_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n640_));
  AOI22_X1  g439(.A1(new_n634_), .A2(new_n639_), .B1(KEYINPUT104), .B2(new_n640_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n624_), .A2(new_n626_), .A3(new_n280_), .ZN(new_n642_));
  INV_X1    g441(.A(G36gat), .ZN(new_n643_));
  OAI211_X1 g442(.A(KEYINPUT104), .B(new_n639_), .C1(new_n642_), .C2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT105), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT46), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n641_), .B1(new_n645_), .B2(new_n646_), .ZN(G1329gat));
  NAND3_X1  g446(.A1(new_n627_), .A2(G43gat), .A3(new_n361_), .ZN(new_n648_));
  AOI21_X1  g447(.A(G43gat), .B1(new_n614_), .B2(new_n361_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g451(.A(G50gat), .B1(new_n614_), .B2(new_n316_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n316_), .A2(G50gat), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n653_), .B1(new_n627_), .B2(new_n654_), .ZN(G1331gat));
  INV_X1    g454(.A(new_n546_), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n388_), .A2(new_n416_), .A3(new_n656_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n657_), .A2(new_n616_), .A3(new_n574_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n658_), .A2(new_n490_), .A3(new_n347_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n571_), .A2(new_n418_), .A3(new_n574_), .A4(new_n546_), .ZN(new_n660_));
  OAI21_X1  g459(.A(G57gat), .B1(new_n660_), .B2(new_n348_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n661_), .ZN(G1332gat));
  OAI21_X1  g461(.A(G64gat), .B1(new_n660_), .B2(new_n280_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT48), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n281_), .A2(new_n492_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT106), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n658_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n664_), .A2(new_n667_), .ZN(G1333gat));
  OAI21_X1  g467(.A(G71gat), .B1(new_n660_), .B2(new_n387_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT49), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n387_), .A2(G71gat), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT107), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n658_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n670_), .A2(new_n673_), .ZN(G1334gat));
  OAI21_X1  g473(.A(G78gat), .B1(new_n660_), .B2(new_n364_), .ZN(new_n675_));
  XOR2_X1   g474(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n676_));
  XNOR2_X1  g475(.A(new_n675_), .B(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(G78gat), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n658_), .A2(new_n678_), .A3(new_n316_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(G1335gat));
  AND3_X1   g479(.A1(new_n657_), .A2(new_n484_), .A3(new_n560_), .ZN(new_n681_));
  INV_X1    g480(.A(G85gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n681_), .A2(new_n682_), .A3(new_n347_), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n617_), .A2(KEYINPUT109), .A3(new_n620_), .ZN(new_n684_));
  AOI21_X1  g483(.A(KEYINPUT109), .B1(new_n617_), .B2(new_n620_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n546_), .A2(new_n572_), .A3(new_n560_), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n686_), .A2(new_n348_), .A3(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n683_), .B1(new_n688_), .B2(new_n682_), .ZN(G1336gat));
  NAND3_X1  g488(.A1(new_n681_), .A2(new_n423_), .A3(new_n281_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n686_), .A2(new_n280_), .A3(new_n687_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n690_), .B1(new_n691_), .B2(new_n423_), .ZN(G1337gat));
  INV_X1    g491(.A(new_n687_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n361_), .B(new_n693_), .C1(new_n684_), .C2(new_n685_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n694_), .A2(KEYINPUT110), .A3(G99gat), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n361_), .A2(new_n432_), .ZN(new_n696_));
  AOI21_X1  g495(.A(KEYINPUT111), .B1(new_n681_), .B2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(KEYINPUT110), .B1(new_n694_), .B2(G99gat), .ZN(new_n699_));
  OAI21_X1  g498(.A(KEYINPUT51), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n699_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT51), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n701_), .A2(new_n702_), .A3(new_n695_), .A4(new_n697_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n700_), .A2(new_n703_), .ZN(G1338gat));
  NAND3_X1  g503(.A1(new_n681_), .A2(new_n433_), .A3(new_n316_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n687_), .A2(new_n364_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n433_), .B1(new_n621_), .B2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT52), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n707_), .A2(new_n708_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n705_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g511(.A(KEYINPUT59), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n281_), .A2(new_n316_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n714_), .A2(new_n347_), .A3(new_n361_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n416_), .A2(new_n540_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT56), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n524_), .A2(new_n526_), .A3(new_n533_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n526_), .A2(new_n533_), .A3(new_n518_), .ZN(new_n720_));
  AOI22_X1  g519(.A1(new_n719_), .A2(KEYINPUT55), .B1(new_n522_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT55), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT113), .B1(new_n534_), .B2(new_n722_), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n534_), .A2(KEYINPUT113), .A3(new_n722_), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n721_), .B(KEYINPUT114), .C1(new_n723_), .C2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n539_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT113), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n728_), .B1(new_n719_), .B2(KEYINPUT55), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n534_), .A2(KEYINPUT113), .A3(new_n722_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(KEYINPUT114), .B1(new_n731_), .B2(new_n721_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n718_), .B1(new_n727_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT114), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n724_), .A2(new_n723_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n721_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n734_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n737_), .A2(KEYINPUT56), .A3(new_n726_), .A4(new_n725_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n717_), .B1(new_n733_), .B2(new_n738_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n409_), .A2(new_n414_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n401_), .A2(new_n402_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(new_n414_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n742_), .A2(KEYINPUT115), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n406_), .A2(new_n407_), .A3(new_n403_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n744_), .B1(new_n742_), .B2(KEYINPUT115), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n740_), .B1(new_n743_), .B2(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n746_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT116), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n747_), .B(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n611_), .B1(new_n739_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT57), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  OAI211_X1 g551(.A(KEYINPUT57), .B(new_n611_), .C1(new_n739_), .C2(new_n749_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n733_), .A2(new_n738_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n746_), .A2(new_n540_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT58), .ZN(new_n759_));
  OAI21_X1  g558(.A(KEYINPUT117), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n616_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT117), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n755_), .A2(new_n762_), .A3(KEYINPUT58), .A4(new_n757_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n760_), .A2(new_n761_), .A3(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n574_), .B1(new_n754_), .B2(new_n764_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(KEYINPUT112), .A2(KEYINPUT54), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n656_), .A2(new_n616_), .A3(new_n574_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n766_), .B1(new_n767_), .B2(new_n417_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n766_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n561_), .A2(new_n418_), .A3(new_n769_), .ZN(new_n770_));
  AOI22_X1  g569(.A1(new_n768_), .A2(new_n770_), .B1(KEYINPUT112), .B2(KEYINPUT54), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n713_), .B(new_n716_), .C1(new_n765_), .C2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT118), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n773_), .B1(new_n765_), .B2(new_n771_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n771_), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n760_), .A2(new_n761_), .A3(new_n763_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n752_), .A2(new_n753_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n560_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n775_), .A2(new_n778_), .A3(KEYINPUT118), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n715_), .B1(new_n774_), .B2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n772_), .B1(new_n780_), .B2(new_n713_), .ZN(new_n781_));
  OAI21_X1  g580(.A(G113gat), .B1(new_n781_), .B2(new_n418_), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n765_), .A2(new_n773_), .A3(new_n771_), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT118), .B1(new_n775_), .B2(new_n778_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n716_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  OR2_X1    g584(.A1(new_n572_), .A2(G113gat), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n782_), .B1(new_n785_), .B2(new_n786_), .ZN(G1340gat));
  OAI21_X1  g586(.A(G120gat), .B1(new_n781_), .B2(new_n656_), .ZN(new_n788_));
  INV_X1    g587(.A(G120gat), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n789_), .B1(new_n656_), .B2(KEYINPUT60), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n790_), .B1(KEYINPUT60), .B2(new_n789_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n788_), .B1(new_n785_), .B2(new_n791_), .ZN(G1341gat));
  INV_X1    g591(.A(G127gat), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n560_), .A2(new_n793_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n772_), .B(new_n794_), .C1(new_n780_), .C2(new_n713_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n574_), .B(new_n716_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n793_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT119), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT119), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n795_), .A2(new_n797_), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(G1342gat));
  INV_X1    g601(.A(G134gat), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n803_), .B1(new_n785_), .B2(new_n611_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT120), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  OAI211_X1 g605(.A(KEYINPUT120), .B(new_n803_), .C1(new_n785_), .C2(new_n611_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n781_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n616_), .A2(new_n803_), .ZN(new_n809_));
  AOI22_X1  g608(.A1(new_n806_), .A2(new_n807_), .B1(new_n808_), .B2(new_n809_), .ZN(G1343gat));
  NOR3_X1   g609(.A1(new_n281_), .A2(new_n364_), .A3(new_n348_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n387_), .B(new_n811_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n812_), .A2(new_n572_), .ZN(new_n813_));
  XOR2_X1   g612(.A(KEYINPUT121), .B(G141gat), .Z(new_n814_));
  XNOR2_X1  g613(.A(new_n813_), .B(new_n814_), .ZN(G1344gat));
  NOR2_X1   g614(.A1(new_n812_), .A2(new_n656_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(new_n284_), .ZN(G1345gat));
  NOR2_X1   g616(.A1(new_n812_), .A2(new_n560_), .ZN(new_n818_));
  XOR2_X1   g617(.A(KEYINPUT61), .B(G155gat), .Z(new_n819_));
  XNOR2_X1  g618(.A(new_n818_), .B(new_n819_), .ZN(G1346gat));
  INV_X1    g619(.A(G162gat), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n812_), .A2(new_n821_), .A3(new_n616_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n812_), .B2(new_n611_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT122), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT122), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n825_), .B(new_n821_), .C1(new_n812_), .C2(new_n611_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n822_), .B1(new_n824_), .B2(new_n826_), .ZN(G1347gat));
  NOR2_X1   g626(.A1(new_n765_), .A2(new_n771_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n280_), .A2(new_n362_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n364_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n416_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT123), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(new_n833_), .A3(G169gat), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n828_), .A2(new_n572_), .A3(new_n830_), .ZN(new_n835_));
  INV_X1    g634(.A(G169gat), .ZN(new_n836_));
  OAI21_X1  g635(.A(KEYINPUT123), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n834_), .A2(KEYINPUT62), .A3(new_n837_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(KEYINPUT22), .B(G169gat), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n835_), .A2(new_n839_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n838_), .B(new_n840_), .C1(KEYINPUT62), .C2(new_n837_), .ZN(G1348gat));
  AOI21_X1  g640(.A(G176gat), .B1(new_n831_), .B2(new_n546_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n316_), .B1(new_n774_), .B2(new_n779_), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n829_), .A2(G176gat), .A3(new_n546_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n842_), .B1(new_n843_), .B2(new_n844_), .ZN(G1349gat));
  NAND3_X1  g644(.A1(new_n843_), .A2(new_n574_), .A3(new_n829_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n223_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n560_), .A2(new_n240_), .ZN(new_n848_));
  AOI22_X1  g647(.A1(new_n846_), .A2(new_n847_), .B1(new_n831_), .B2(new_n848_), .ZN(G1350gat));
  NOR2_X1   g648(.A1(new_n611_), .A2(new_n232_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n831_), .A2(new_n850_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n828_), .A2(new_n616_), .A3(new_n830_), .ZN(new_n852_));
  INV_X1    g651(.A(G190gat), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n851_), .B1(new_n852_), .B2(new_n853_), .ZN(G1351gat));
  AOI21_X1  g653(.A(new_n361_), .B1(new_n774_), .B2(new_n779_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n280_), .A2(new_n383_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(new_n416_), .A3(new_n856_), .ZN(new_n857_));
  XOR2_X1   g656(.A(KEYINPUT124), .B(G197gat), .Z(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(G1352gat));
  OR2_X1    g658(.A1(new_n209_), .A2(KEYINPUT125), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n855_), .A2(new_n546_), .A3(new_n856_), .A4(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n209_), .A2(KEYINPUT125), .ZN(new_n862_));
  XOR2_X1   g661(.A(new_n862_), .B(KEYINPUT126), .Z(new_n863_));
  XNOR2_X1  g662(.A(new_n861_), .B(new_n863_), .ZN(G1353gat));
  NAND2_X1  g663(.A1(new_n855_), .A2(new_n856_), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT127), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(KEYINPUT127), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n868_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n574_), .A2(new_n869_), .ZN(new_n870_));
  OR3_X1    g669(.A1(new_n865_), .A2(new_n867_), .A3(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n867_), .B1(new_n865_), .B2(new_n870_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(G1354gat));
  OAI21_X1  g672(.A(G218gat), .B1(new_n865_), .B2(new_n616_), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n611_), .A2(G218gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n865_), .B2(new_n875_), .ZN(G1355gat));
endmodule


