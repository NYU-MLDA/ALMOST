//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 0 0 0 1 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n794_, new_n795_,
    new_n796_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n806_, new_n808_, new_n809_, new_n810_, new_n812_,
    new_n813_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n839_, new_n840_, new_n841_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_;
  XNOR2_X1  g000(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT25), .B(G183gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT26), .B(G190gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT83), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT23), .ZN(new_n209_));
  INV_X1    g008(.A(G169gat), .ZN(new_n210_));
  INV_X1    g009(.A(G176gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT24), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  MUX2_X1   g012(.A(new_n212_), .B(KEYINPUT24), .S(new_n213_), .Z(new_n214_));
  NAND3_X1  g013(.A1(new_n207_), .A2(new_n209_), .A3(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n210_), .A2(new_n211_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT22), .B(G169gat), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n216_), .B1(new_n217_), .B2(new_n211_), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n208_), .A2(KEYINPUT23), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n219_), .A2(KEYINPUT84), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n220_), .B1(KEYINPUT84), .B2(new_n209_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n218_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n215_), .A2(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(G211gat), .B(G218gat), .Z(new_n225_));
  XOR2_X1   g024(.A(G197gat), .B(G204gat), .Z(new_n226_));
  AOI21_X1  g025(.A(new_n225_), .B1(KEYINPUT21), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT86), .ZN(new_n228_));
  INV_X1    g027(.A(G204gat), .ZN(new_n229_));
  NOR3_X1   g028(.A1(new_n228_), .A2(new_n229_), .A3(G197gat), .ZN(new_n230_));
  INV_X1    g029(.A(G197gat), .ZN(new_n231_));
  AOI21_X1  g030(.A(KEYINPUT86), .B1(new_n231_), .B2(G204gat), .ZN(new_n232_));
  OAI22_X1  g031(.A1(new_n230_), .A2(new_n232_), .B1(new_n231_), .B2(G204gat), .ZN(new_n233_));
  XOR2_X1   g032(.A(KEYINPUT87), .B(KEYINPUT21), .Z(new_n234_));
  OAI21_X1  g033(.A(new_n227_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT88), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n225_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n225_), .A2(new_n236_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n233_), .A2(new_n238_), .A3(KEYINPUT21), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n235_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n224_), .A2(new_n240_), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n209_), .A2(KEYINPUT84), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n214_), .B(new_n206_), .C1(new_n242_), .C2(new_n220_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n209_), .B1(G183gat), .B2(G190gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(new_n218_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n241_), .B(KEYINPUT20), .C1(new_n240_), .C2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G226gat), .A2(G233gat), .ZN(new_n248_));
  XOR2_X1   g047(.A(new_n248_), .B(KEYINPUT90), .Z(new_n249_));
  XOR2_X1   g048(.A(new_n249_), .B(KEYINPUT19), .Z(new_n250_));
  OR2_X1    g049(.A1(new_n247_), .A2(new_n250_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n246_), .A2(new_n240_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT91), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n224_), .A2(new_n240_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n254_), .A2(KEYINPUT20), .ZN(new_n255_));
  AND2_X1   g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n250_), .ZN(new_n257_));
  OAI211_X1 g056(.A(KEYINPUT92), .B(new_n251_), .C1(new_n256_), .C2(new_n257_), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n251_), .A2(KEYINPUT92), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  XOR2_X1   g059(.A(G8gat), .B(G36gat), .Z(new_n261_));
  XNOR2_X1  g060(.A(G64gat), .B(G92gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n264_));
  XOR2_X1   g063(.A(new_n263_), .B(new_n264_), .Z(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n260_), .A2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n258_), .A2(new_n265_), .A3(new_n259_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(KEYINPUT94), .A3(new_n268_), .ZN(new_n269_));
  OR3_X1    g068(.A1(new_n260_), .A2(KEYINPUT94), .A3(new_n266_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT27), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  AND3_X1   g071(.A1(new_n253_), .A2(new_n255_), .A3(new_n257_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT99), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n247_), .A2(new_n250_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n273_), .A2(new_n274_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n266_), .A2(KEYINPUT100), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n266_), .A2(KEYINPUT100), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n278_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n281_), .A2(KEYINPUT27), .A3(new_n267_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n272_), .A2(new_n282_), .ZN(new_n283_));
  AND2_X1   g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284_));
  NOR2_X1   g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(G141gat), .A2(G148gat), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n287_), .B(KEYINPUT3), .Z(new_n288_));
  NAND2_X1  g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n289_), .B(KEYINPUT2), .Z(new_n290_));
  OAI21_X1  g089(.A(new_n286_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT1), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n287_), .B1(new_n286_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n284_), .A2(KEYINPUT1), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n293_), .A2(new_n294_), .A3(new_n289_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n291_), .A2(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n296_), .A2(KEYINPUT29), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G22gat), .B(G50gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT28), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n297_), .B(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT89), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n296_), .A2(KEYINPUT29), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(new_n240_), .ZN(new_n303_));
  INV_X1    g102(.A(G228gat), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n304_), .A2(KEYINPUT85), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n304_), .A2(KEYINPUT85), .ZN(new_n306_));
  OAI21_X1  g105(.A(G233gat), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n303_), .B(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(G78gat), .B(G106gat), .Z(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  MUX2_X1   g109(.A(new_n300_), .B(new_n301_), .S(new_n310_), .Z(new_n311_));
  OR2_X1    g110(.A1(new_n308_), .A2(new_n309_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n312_), .A2(new_n301_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n283_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G127gat), .B(G134gat), .ZN(new_n317_));
  INV_X1    g116(.A(G113gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(G120gat), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n320_), .A2(new_n296_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n296_), .ZN(new_n322_));
  AND2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G225gat), .A2(G233gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  OR2_X1    g124(.A1(new_n325_), .A2(KEYINPUT97), .ZN(new_n326_));
  INV_X1    g125(.A(new_n324_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT4), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n322_), .A2(KEYINPUT95), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n328_), .B1(new_n330_), .B2(new_n321_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n329_), .A2(KEYINPUT4), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n327_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n325_), .A2(KEYINPUT97), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n326_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  XOR2_X1   g134(.A(G1gat), .B(G29gat), .Z(new_n336_));
  XNOR2_X1  g135(.A(G57gat), .B(G85gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n338_), .B(new_n339_), .Z(new_n340_));
  NAND2_X1  g139(.A1(new_n335_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n340_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n326_), .A2(new_n333_), .A3(new_n334_), .A4(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n224_), .B(KEYINPUT30), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(new_n320_), .ZN(new_n347_));
  XOR2_X1   g146(.A(G15gat), .B(G43gat), .Z(new_n348_));
  XOR2_X1   g147(.A(new_n348_), .B(KEYINPUT31), .Z(new_n349_));
  XNOR2_X1  g148(.A(new_n347_), .B(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G71gat), .B(G99gat), .Z(new_n351_));
  NAND2_X1  g150(.A1(G227gat), .A2(G233gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  OR2_X1    g153(.A1(new_n350_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n350_), .A2(new_n354_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n316_), .A2(new_n345_), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n324_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(new_n340_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n361_), .B1(new_n327_), .B2(new_n323_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n362_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(KEYINPUT98), .A2(KEYINPUT33), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n343_), .B(new_n364_), .Z(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n315_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n260_), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n266_), .A2(KEYINPUT32), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n344_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n278_), .A2(new_n369_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n366_), .A2(new_n367_), .A3(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n357_), .B1(new_n283_), .B2(new_n315_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n367_), .A2(new_n345_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n374_), .A2(new_n375_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT101), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n372_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n376_), .B1(new_n381_), .B2(new_n367_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n382_), .A2(KEYINPUT101), .A3(new_n375_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n359_), .B1(new_n380_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT64), .ZN(new_n385_));
  XOR2_X1   g184(.A(KEYINPUT10), .B(G99gat), .Z(new_n386_));
  INV_X1    g185(.A(G106gat), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n385_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT10), .B(G99gat), .ZN(new_n389_));
  NOR3_X1   g188(.A1(new_n389_), .A2(KEYINPUT64), .A3(G106gat), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G99gat), .A2(G106gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT6), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT6), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n394_), .A2(G99gat), .A3(G106gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT9), .ZN(new_n397_));
  OR2_X1    g196(.A1(G85gat), .A2(G92gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G85gat), .A2(G92gat), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n397_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT65), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  OR3_X1    g201(.A1(new_n400_), .A2(KEYINPUT65), .A3(new_n401_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n391_), .A2(new_n396_), .A3(new_n402_), .A4(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT8), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n398_), .A2(new_n399_), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n393_), .A2(new_n395_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT7), .ZN(new_n408_));
  INV_X1    g207(.A(G99gat), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(new_n409_), .A3(new_n387_), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n405_), .B(new_n406_), .C1(new_n407_), .C2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT66), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n396_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n416_), .A2(KEYINPUT66), .A3(new_n405_), .A4(new_n406_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT67), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n396_), .A2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n393_), .A2(new_n395_), .A3(KEYINPUT67), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n420_), .A2(new_n410_), .A3(new_n411_), .A4(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n405_), .B1(new_n422_), .B2(new_n406_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n404_), .B1(new_n418_), .B2(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G43gat), .B(G50gat), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  AND2_X1   g225(.A1(G29gat), .A2(G36gat), .ZN(new_n427_));
  NOR2_X1   g226(.A1(G29gat), .A2(G36gat), .ZN(new_n428_));
  NOR3_X1   g227(.A1(new_n427_), .A2(new_n428_), .A3(KEYINPUT72), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT72), .ZN(new_n430_));
  INV_X1    g229(.A(G29gat), .ZN(new_n431_));
  INV_X1    g230(.A(G36gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G29gat), .A2(G36gat), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n430_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n426_), .B1(new_n429_), .B2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT72), .B1(new_n427_), .B2(new_n428_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n433_), .A2(new_n430_), .A3(new_n434_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(new_n425_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n436_), .A2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT15), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n424_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G232gat), .A2(G233gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT34), .ZN(new_n444_));
  INV_X1    g243(.A(new_n440_), .ZN(new_n445_));
  OAI221_X1 g244(.A(new_n442_), .B1(KEYINPUT35), .B2(new_n444_), .C1(new_n445_), .C2(new_n424_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(KEYINPUT35), .ZN(new_n447_));
  XOR2_X1   g246(.A(new_n446_), .B(new_n447_), .Z(new_n448_));
  XNOR2_X1  g247(.A(G190gat), .B(G218gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(G134gat), .ZN(new_n450_));
  INV_X1    g249(.A(G162gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT36), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n448_), .A2(new_n454_), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n452_), .A2(new_n453_), .ZN(new_n456_));
  OR2_X1    g255(.A1(new_n448_), .A2(new_n456_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n455_), .B(new_n457_), .C1(KEYINPUT73), .C2(KEYINPUT37), .ZN(new_n458_));
  NAND2_X1  g257(.A1(KEYINPUT73), .A2(KEYINPUT37), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(G127gat), .B(G155gat), .Z(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT75), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G183gat), .B(G211gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  XOR2_X1   g263(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT17), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G57gat), .B(G64gat), .ZN(new_n469_));
  OR2_X1    g268(.A1(new_n469_), .A2(KEYINPUT11), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(KEYINPUT11), .ZN(new_n471_));
  XOR2_X1   g270(.A(G71gat), .B(G78gat), .Z(new_n472_));
  NAND3_X1  g271(.A1(new_n470_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n471_), .A2(new_n472_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G15gat), .B(G22gat), .ZN(new_n476_));
  INV_X1    g275(.A(G1gat), .ZN(new_n477_));
  INV_X1    g276(.A(G8gat), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT14), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n476_), .A2(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(G1gat), .B(G8gat), .Z(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n475_), .B(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G231gat), .A2(G233gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n468_), .A2(new_n485_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n466_), .A2(KEYINPUT17), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n468_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n486_), .B1(new_n489_), .B2(new_n485_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n460_), .A2(new_n491_), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n492_), .B(KEYINPUT76), .Z(new_n493_));
  NOR2_X1   g292(.A1(new_n384_), .A2(new_n493_), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n404_), .B(new_n475_), .C1(new_n418_), .C2(new_n423_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G230gat), .A2(G233gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT69), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n475_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n424_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT12), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n424_), .A2(KEYINPUT12), .A3(new_n500_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n495_), .A2(KEYINPUT69), .A3(new_n496_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n499_), .A2(new_n503_), .A3(new_n504_), .A4(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(KEYINPUT68), .B1(new_n424_), .B2(new_n500_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(new_n495_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n506_), .B1(new_n508_), .B2(new_n496_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT70), .B(G204gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G120gat), .B(G148gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT5), .B(G176gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n509_), .B(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT13), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n516_), .B(KEYINPUT71), .Z(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G229gat), .A2(G233gat), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT77), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n437_), .A2(new_n438_), .A3(new_n425_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n425_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n521_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n436_), .A2(KEYINPUT77), .A3(new_n439_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n524_), .A2(new_n482_), .A3(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT78), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT78), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n524_), .A2(new_n482_), .A3(new_n525_), .A4(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n482_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(KEYINPUT79), .B1(new_n530_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT79), .ZN(new_n534_));
  AOI211_X1 g333(.A(new_n534_), .B(new_n531_), .C1(new_n527_), .C2(new_n529_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n520_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT80), .ZN(new_n537_));
  INV_X1    g336(.A(new_n482_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n441_), .A2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n530_), .A2(new_n539_), .A3(new_n519_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT80), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n541_), .B(new_n520_), .C1(new_n533_), .C2(new_n535_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n537_), .A2(new_n540_), .A3(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G113gat), .B(G141gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(G197gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT81), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(new_n210_), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n543_), .A2(new_n547_), .ZN(new_n548_));
  AND2_X1   g347(.A1(new_n537_), .A2(new_n542_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT82), .ZN(new_n550_));
  INV_X1    g349(.A(new_n547_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n549_), .A2(new_n550_), .A3(new_n540_), .A4(new_n551_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n537_), .A2(new_n540_), .A3(new_n542_), .A4(new_n551_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT82), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n548_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n518_), .A2(new_n555_), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n494_), .A2(new_n477_), .A3(new_n556_), .ZN(new_n557_));
  AND3_X1   g356(.A1(new_n557_), .A2(KEYINPUT102), .A3(new_n344_), .ZN(new_n558_));
  AOI21_X1  g357(.A(KEYINPUT102), .B1(new_n557_), .B2(new_n344_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n203_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT104), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  OR3_X1    g361(.A1(new_n558_), .A2(new_n559_), .A3(new_n203_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n383_), .ZN(new_n564_));
  AOI21_X1  g363(.A(KEYINPUT101), .B1(new_n382_), .B2(new_n375_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n358_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n457_), .A2(new_n455_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n516_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n568_), .A2(new_n555_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n566_), .A2(new_n567_), .A3(new_n491_), .A4(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(G1gat), .B1(new_n570_), .B2(new_n345_), .ZN(new_n571_));
  OAI211_X1 g370(.A(KEYINPUT104), .B(new_n203_), .C1(new_n558_), .C2(new_n559_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n562_), .A2(new_n563_), .A3(new_n571_), .A4(new_n572_), .ZN(G1324gat));
  INV_X1    g372(.A(KEYINPUT40), .ZN(new_n574_));
  INV_X1    g373(.A(new_n283_), .ZN(new_n575_));
  OAI21_X1  g374(.A(G8gat), .B1(new_n570_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT39), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT39), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n578_), .B(G8gat), .C1(new_n570_), .C2(new_n575_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT105), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n494_), .A2(new_n556_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n582_), .A2(new_n478_), .A3(new_n283_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n580_), .A2(new_n581_), .A3(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n581_), .B1(new_n580_), .B2(new_n583_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n574_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n579_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n567_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n384_), .A2(new_n589_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n590_), .A2(new_n283_), .A3(new_n491_), .A4(new_n569_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n578_), .B1(new_n591_), .B2(G8gat), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n583_), .B1(new_n588_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT105), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(KEYINPUT40), .A3(new_n584_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n587_), .A2(new_n595_), .ZN(G1325gat));
  INV_X1    g395(.A(new_n357_), .ZN(new_n597_));
  OAI21_X1  g396(.A(G15gat), .B1(new_n570_), .B2(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT41), .Z(new_n599_));
  INV_X1    g398(.A(G15gat), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n582_), .A2(new_n600_), .A3(new_n357_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(G1326gat));
  OAI21_X1  g401(.A(G22gat), .B1(new_n570_), .B2(new_n367_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT42), .ZN(new_n604_));
  INV_X1    g403(.A(G22gat), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n582_), .A2(new_n605_), .A3(new_n315_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(G1327gat));
  NAND2_X1  g406(.A1(new_n569_), .A2(new_n490_), .ZN(new_n608_));
  NOR3_X1   g407(.A1(new_n384_), .A2(new_n567_), .A3(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(G29gat), .B1(new_n609_), .B2(new_n344_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n608_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT43), .ZN(new_n612_));
  INV_X1    g411(.A(new_n460_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n612_), .B1(new_n566_), .B2(new_n613_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n384_), .A2(KEYINPUT43), .A3(new_n460_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n611_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT44), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n616_), .A2(KEYINPUT106), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT106), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n566_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n620_));
  OAI21_X1  g419(.A(KEYINPUT43), .B1(new_n384_), .B2(new_n460_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n608_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n619_), .B1(new_n622_), .B2(KEYINPUT44), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n345_), .B1(new_n618_), .B2(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n431_), .B1(new_n622_), .B2(KEYINPUT44), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n610_), .B1(new_n624_), .B2(new_n625_), .ZN(G1328gat));
  INV_X1    g425(.A(KEYINPUT107), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n627_), .A2(KEYINPUT46), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n618_), .A2(new_n623_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n575_), .B1(new_n622_), .B2(KEYINPUT44), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n432_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n609_), .A2(new_n432_), .A3(new_n283_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT45), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n628_), .B1(new_n631_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n628_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n622_), .A2(KEYINPUT44), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(new_n283_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n638_), .B1(new_n623_), .B2(new_n618_), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n636_), .B(new_n633_), .C1(new_n639_), .C2(new_n432_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n635_), .A2(new_n640_), .ZN(G1329gat));
  INV_X1    g440(.A(G43gat), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n642_), .B1(new_n622_), .B2(KEYINPUT44), .ZN(new_n643_));
  AOI21_X1  g442(.A(KEYINPUT106), .B1(new_n616_), .B2(new_n617_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n622_), .A2(new_n619_), .A3(KEYINPUT44), .ZN(new_n645_));
  OAI211_X1 g444(.A(new_n357_), .B(new_n643_), .C1(new_n644_), .C2(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(G43gat), .B1(new_n609_), .B2(new_n357_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT108), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(KEYINPUT47), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT47), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n646_), .A2(new_n651_), .A3(new_n648_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(G1330gat));
  INV_X1    g452(.A(G50gat), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n315_), .A2(new_n654_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT109), .Z(new_n656_));
  NAND2_X1  g455(.A1(new_n609_), .A2(new_n656_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n629_), .A2(new_n315_), .A3(new_n637_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n657_), .B1(new_n658_), .B2(new_n654_), .ZN(G1331gat));
  NAND2_X1  g458(.A1(new_n568_), .A2(new_n555_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n384_), .A2(new_n493_), .A3(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(G57gat), .B1(new_n661_), .B2(new_n344_), .ZN(new_n662_));
  AND4_X1   g461(.A1(new_n491_), .A2(new_n590_), .A3(new_n555_), .A4(new_n518_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n663_), .A2(new_n344_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n662_), .B1(new_n664_), .B2(G57gat), .ZN(G1332gat));
  INV_X1    g464(.A(G64gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(new_n663_), .B2(new_n283_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT48), .Z(new_n668_));
  NAND3_X1  g467(.A1(new_n661_), .A2(new_n666_), .A3(new_n283_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1333gat));
  INV_X1    g469(.A(G71gat), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n671_), .B1(new_n663_), .B2(new_n357_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT49), .Z(new_n673_));
  NAND2_X1  g472(.A1(new_n357_), .A2(new_n671_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT110), .Z(new_n675_));
  NAND2_X1  g474(.A1(new_n661_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n673_), .A2(new_n676_), .ZN(G1334gat));
  INV_X1    g476(.A(G78gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n678_), .B1(new_n663_), .B2(new_n315_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT50), .Z(new_n680_));
  NAND3_X1  g479(.A1(new_n661_), .A2(new_n678_), .A3(new_n315_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1335gat));
  NAND3_X1  g481(.A1(new_n518_), .A2(new_n490_), .A3(new_n555_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n384_), .A2(new_n567_), .A3(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G85gat), .B1(new_n684_), .B2(new_n344_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n660_), .A2(new_n491_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT111), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n689_), .A2(new_n344_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n685_), .B1(new_n690_), .B2(G85gat), .ZN(G1336gat));
  INV_X1    g490(.A(G92gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n689_), .B2(new_n283_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n684_), .A2(new_n692_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n283_), .B2(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT112), .ZN(G1337gat));
  NAND3_X1  g495(.A1(new_n684_), .A2(new_n357_), .A3(new_n386_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n689_), .A2(new_n357_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n697_), .B1(new_n698_), .B2(new_n409_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g499(.A1(new_n684_), .A2(new_n387_), .A3(new_n315_), .ZN(new_n701_));
  OAI211_X1 g500(.A(new_n315_), .B(new_n687_), .C1(new_n614_), .C2(new_n615_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT52), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n702_), .A2(new_n703_), .A3(G106gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n702_), .B2(G106gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n701_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g506(.A1(new_n460_), .A2(new_n491_), .A3(new_n555_), .A4(new_n516_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT54), .Z(new_n709_));
  NOR2_X1   g508(.A1(new_n509_), .A2(new_n514_), .ZN(new_n710_));
  OAI21_X1  g509(.A(KEYINPUT113), .B1(new_n555_), .B2(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n503_), .A2(new_n504_), .A3(new_n495_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n496_), .ZN(new_n714_));
  AOI22_X1  g513(.A1(new_n506_), .A2(new_n712_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT115), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT55), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(new_n506_), .B2(new_n717_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n503_), .A2(new_n504_), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n495_), .A2(KEYINPUT69), .A3(new_n496_), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT69), .B1(new_n495_), .B2(new_n496_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n719_), .A2(new_n722_), .A3(KEYINPUT115), .A4(KEYINPUT55), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n715_), .A2(new_n718_), .A3(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT116), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT116), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n715_), .A2(new_n718_), .A3(new_n726_), .A4(new_n723_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n725_), .A2(new_n514_), .A3(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT117), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT56), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n543_), .A2(new_n547_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n553_), .A2(KEYINPUT82), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n553_), .A2(KEYINPUT82), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n732_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT113), .ZN(new_n736_));
  INV_X1    g535(.A(new_n710_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n735_), .A2(new_n736_), .A3(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n728_), .A2(KEYINPUT117), .A3(KEYINPUT56), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n711_), .A2(new_n731_), .A3(new_n738_), .A4(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT118), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n728_), .A2(KEYINPUT117), .A3(KEYINPUT56), .ZN(new_n743_));
  AOI21_X1  g542(.A(KEYINPUT56), .B1(new_n728_), .B2(KEYINPUT117), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n745_), .A2(KEYINPUT118), .A3(new_n711_), .A4(new_n738_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n519_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n530_), .A2(new_n539_), .A3(new_n520_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  AOI22_X1  g548(.A1(new_n552_), .A2(new_n554_), .B1(new_n547_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n515_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n742_), .A2(new_n746_), .A3(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(new_n567_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT57), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n752_), .A2(KEYINPUT57), .A3(new_n567_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n728_), .A2(KEYINPUT56), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n757_), .A2(new_n750_), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n728_), .A2(KEYINPUT56), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n758_), .A2(new_n737_), .A3(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT58), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n758_), .A2(KEYINPUT58), .A3(new_n737_), .A4(new_n759_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n762_), .A2(new_n613_), .A3(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n755_), .A2(new_n756_), .A3(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n709_), .B1(new_n765_), .B2(new_n490_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n316_), .A2(new_n344_), .A3(new_n357_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(G113gat), .B1(new_n768_), .B2(new_n735_), .ZN(new_n769_));
  OAI21_X1  g568(.A(KEYINPUT59), .B1(new_n766_), .B2(new_n767_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n755_), .A2(KEYINPUT119), .A3(new_n764_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT119), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT57), .B1(new_n752_), .B2(new_n567_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n764_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n772_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n771_), .A2(new_n756_), .A3(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n709_), .B1(new_n776_), .B2(new_n490_), .ZN(new_n777_));
  OR2_X1    g576(.A1(new_n767_), .A2(KEYINPUT59), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n770_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n779_), .B1(KEYINPUT120), .B2(new_n318_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT120), .ZN(new_n781_));
  OAI21_X1  g580(.A(G113gat), .B1(new_n555_), .B2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n769_), .B1(new_n780_), .B2(new_n782_), .ZN(G1340gat));
  XOR2_X1   g582(.A(KEYINPUT121), .B(G120gat), .Z(new_n784_));
  OAI21_X1  g583(.A(new_n784_), .B1(new_n779_), .B2(new_n517_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n784_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n786_), .B1(new_n516_), .B2(KEYINPUT60), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n768_), .B(new_n787_), .C1(KEYINPUT60), .C2(new_n786_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n785_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT122), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n785_), .A2(KEYINPUT122), .A3(new_n788_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(G1341gat));
  AOI21_X1  g592(.A(G127gat), .B1(new_n768_), .B2(new_n491_), .ZN(new_n794_));
  INV_X1    g593(.A(G127gat), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n779_), .A2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n794_), .B1(new_n796_), .B2(new_n491_), .ZN(G1342gat));
  AOI21_X1  g596(.A(G134gat), .B1(new_n768_), .B2(new_n589_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n779_), .A2(new_n460_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(G134gat), .ZN(G1343gat));
  NOR2_X1   g599(.A1(new_n766_), .A2(new_n283_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n377_), .A2(new_n357_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n803_), .A2(new_n555_), .ZN(new_n804_));
  XOR2_X1   g603(.A(new_n804_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g604(.A1(new_n803_), .A2(new_n517_), .ZN(new_n806_));
  XOR2_X1   g605(.A(new_n806_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g606(.A1(new_n803_), .A2(new_n490_), .ZN(new_n808_));
  XOR2_X1   g607(.A(KEYINPUT61), .B(G155gat), .Z(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT123), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n808_), .B(new_n810_), .ZN(G1346gat));
  NOR3_X1   g610(.A1(new_n803_), .A2(new_n451_), .A3(new_n460_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n801_), .A2(new_n589_), .A3(new_n802_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n451_), .B2(new_n813_), .ZN(G1347gat));
  NAND2_X1  g613(.A1(new_n776_), .A2(new_n490_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n709_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n283_), .A2(new_n345_), .A3(new_n357_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n818_), .A2(new_n315_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n817_), .A2(new_n735_), .A3(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(G169gat), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT124), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT62), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n821_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n756_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n755_), .A2(new_n764_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(new_n772_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n491_), .B1(new_n827_), .B2(new_n771_), .ZN(new_n828_));
  OAI211_X1 g627(.A(KEYINPUT125), .B(new_n819_), .C1(new_n828_), .C2(new_n709_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT125), .ZN(new_n830_));
  INV_X1    g629(.A(new_n819_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n777_), .B2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n829_), .A2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n833_), .A2(new_n217_), .A3(new_n735_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n822_), .A2(new_n823_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n820_), .A2(G169gat), .A3(new_n835_), .A4(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n824_), .A2(new_n834_), .A3(new_n837_), .ZN(G1348gat));
  OR2_X1    g637(.A1(new_n766_), .A2(new_n315_), .ZN(new_n839_));
  NOR4_X1   g638(.A1(new_n839_), .A2(new_n211_), .A3(new_n517_), .A4(new_n818_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n833_), .A2(new_n568_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n840_), .B1(new_n841_), .B2(new_n211_), .ZN(G1349gat));
  NOR2_X1   g641(.A1(new_n839_), .A2(new_n818_), .ZN(new_n843_));
  AOI21_X1  g642(.A(G183gat), .B1(new_n843_), .B2(new_n491_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n204_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n490_), .B1(new_n829_), .B2(new_n832_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n844_), .B1(new_n845_), .B2(new_n846_), .ZN(G1350gat));
  NAND3_X1  g646(.A1(new_n833_), .A2(new_n205_), .A3(new_n589_), .ZN(new_n848_));
  AOI21_X1  g647(.A(KEYINPUT125), .B1(new_n817_), .B2(new_n819_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n777_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n613_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT126), .B1(new_n851_), .B2(G190gat), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n460_), .B1(new_n829_), .B2(new_n832_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT126), .ZN(new_n854_));
  INV_X1    g653(.A(G190gat), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n853_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n848_), .B1(new_n852_), .B2(new_n856_), .ZN(G1351gat));
  NOR3_X1   g656(.A1(new_n766_), .A2(new_n344_), .A3(new_n575_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n357_), .A2(new_n367_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n858_), .A2(new_n735_), .A3(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(KEYINPUT127), .A2(G197gat), .ZN(new_n861_));
  OR2_X1    g660(.A1(KEYINPUT127), .A2(G197gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n860_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(new_n860_), .B2(new_n862_), .ZN(G1352gat));
  NAND2_X1  g663(.A1(new_n858_), .A2(new_n859_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n865_), .A2(new_n517_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(new_n229_), .ZN(G1353gat));
  NOR2_X1   g666(.A1(new_n865_), .A2(new_n490_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n868_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n869_));
  XOR2_X1   g668(.A(KEYINPUT63), .B(G211gat), .Z(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(new_n868_), .B2(new_n870_), .ZN(G1354gat));
  NOR2_X1   g670(.A1(new_n865_), .A2(new_n567_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n872_), .A2(G218gat), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n865_), .A2(new_n460_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n873_), .B1(G218gat), .B2(new_n874_), .ZN(G1355gat));
endmodule


