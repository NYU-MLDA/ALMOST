//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 0 1 1 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 1 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n816_,
    new_n817_, new_n819_, new_n820_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_;
  NAND2_X1  g000(.A1(G1gat), .A2(G8gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT14), .ZN(new_n203_));
  INV_X1    g002(.A(G22gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G15gat), .ZN(new_n205_));
  INV_X1    g004(.A(G15gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G22gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n203_), .A2(new_n205_), .A3(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT72), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(G1gat), .B(G8gat), .Z(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G29gat), .B(G36gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G43gat), .B(G50gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n211_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n210_), .B(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n215_), .B(KEYINPUT15), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G229gat), .A2(G233gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n216_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT75), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n215_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n218_), .A2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n212_), .A2(new_n215_), .ZN(new_n227_));
  OAI211_X1 g026(.A(G229gat), .B(G233gat), .C1(new_n226_), .C2(new_n227_), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n216_), .A2(new_n220_), .A3(KEYINPUT75), .A4(new_n221_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n224_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G113gat), .B(G141gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G169gat), .B(G197gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n230_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n233_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n224_), .A2(new_n228_), .A3(new_n229_), .A4(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(G155gat), .A2(G162gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G155gat), .A2(G162gat), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n239_), .B1(KEYINPUT1), .B2(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n241_), .B1(KEYINPUT1), .B2(new_n240_), .ZN(new_n242_));
  INV_X1    g041(.A(G141gat), .ZN(new_n243_));
  INV_X1    g042(.A(G148gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G141gat), .A2(G148gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n242_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT84), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n243_), .A2(new_n244_), .A3(KEYINPUT3), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n250_), .B1(G141gat), .B2(G148gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n246_), .A2(KEYINPUT2), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT2), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n254_), .A2(G141gat), .A3(G148gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n252_), .A2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G155gat), .B(G162gat), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n248_), .B1(new_n257_), .B2(new_n259_), .ZN(new_n260_));
  AOI211_X1 g059(.A(KEYINPUT84), .B(new_n258_), .C1(new_n252_), .C2(new_n256_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n247_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT85), .ZN(new_n263_));
  XOR2_X1   g062(.A(G127gat), .B(G134gat), .Z(new_n264_));
  XNOR2_X1  g063(.A(G113gat), .B(G120gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT85), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n267_), .B(new_n247_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n263_), .A2(new_n266_), .A3(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT89), .B1(new_n262_), .B2(new_n266_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n263_), .A2(KEYINPUT89), .A3(new_n266_), .A4(new_n268_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(KEYINPUT4), .A3(new_n272_), .ZN(new_n273_));
  OR2_X1    g072(.A1(new_n269_), .A2(KEYINPUT4), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G225gat), .A2(G233gat), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  XOR2_X1   g077(.A(G57gat), .B(G85gat), .Z(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT90), .B(KEYINPUT0), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G1gat), .B(G29gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT91), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n281_), .B(new_n283_), .Z(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n277_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n278_), .A2(KEYINPUT92), .A3(new_n285_), .A4(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n276_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n284_), .B1(new_n289_), .B2(new_n286_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n286_), .B1(new_n275_), .B2(new_n277_), .ZN(new_n292_));
  AOI21_X1  g091(.A(KEYINPUT92), .B1(new_n292_), .B2(new_n285_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G71gat), .B(G99gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT81), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(G43gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G227gat), .A2(G233gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(new_n206_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n297_), .B(new_n299_), .ZN(new_n300_));
  OR2_X1    g099(.A1(KEYINPUT79), .A2(G176gat), .ZN(new_n301_));
  INV_X1    g100(.A(G169gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT22), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT22), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(G169gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(KEYINPUT79), .A2(G176gat), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n301_), .A2(new_n303_), .A3(new_n305_), .A4(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT80), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT78), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(KEYINPUT78), .A2(G183gat), .A3(G190gat), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n313_), .A2(KEYINPUT23), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT23), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n316_), .A2(G183gat), .A3(G190gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(G183gat), .ZN(new_n319_));
  INV_X1    g118(.A(G190gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n318_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT80), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n307_), .A2(new_n323_), .A3(new_n308_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n310_), .A2(new_n322_), .A3(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n313_), .A2(new_n316_), .A3(new_n314_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT76), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n329_), .B1(new_n320_), .B2(KEYINPUT26), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT25), .B(G183gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT26), .B(G190gat), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n330_), .B(new_n331_), .C1(new_n332_), .C2(new_n329_), .ZN(new_n333_));
  INV_X1    g132(.A(G176gat), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n302_), .A2(new_n334_), .A3(KEYINPUT77), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT77), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n336_), .B1(G169gat), .B2(G176gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT24), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n335_), .A2(new_n337_), .A3(KEYINPUT24), .A4(new_n308_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n328_), .A2(new_n333_), .A3(new_n340_), .A4(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n325_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT30), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n300_), .A2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT82), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n346_), .B1(new_n300_), .B2(new_n344_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n266_), .B(KEYINPUT31), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n348_), .A2(KEYINPUT83), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n347_), .B(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT94), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n263_), .A2(new_n268_), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n352_), .A2(KEYINPUT29), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n353_), .B(KEYINPUT28), .Z(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n263_), .A2(KEYINPUT29), .A3(new_n268_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT86), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n263_), .A2(KEYINPUT86), .A3(KEYINPUT29), .A4(new_n268_), .ZN(new_n359_));
  XOR2_X1   g158(.A(G197gat), .B(G204gat), .Z(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G211gat), .B(G218gat), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n361_), .A2(KEYINPUT21), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT21), .ZN(new_n364_));
  INV_X1    g163(.A(G218gat), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n365_), .A2(G211gat), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n365_), .A2(G211gat), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n364_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n362_), .A2(KEYINPUT21), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(new_n369_), .A3(new_n360_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n363_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G228gat), .A2(G233gat), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n358_), .A2(new_n359_), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n371_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n375_), .B1(new_n262_), .B2(KEYINPUT29), .ZN(new_n376_));
  OR2_X1    g175(.A1(new_n376_), .A2(new_n372_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G78gat), .B(G106gat), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n374_), .A2(new_n377_), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n379_), .B1(new_n374_), .B2(new_n377_), .ZN(new_n382_));
  XOR2_X1   g181(.A(G22gat), .B(G50gat), .Z(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NOR3_X1   g183(.A1(new_n381_), .A2(new_n382_), .A3(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n374_), .A2(new_n377_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(new_n378_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n383_), .B1(new_n387_), .B2(new_n380_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n355_), .B1(new_n385_), .B2(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n384_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n387_), .A2(new_n380_), .A3(new_n383_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(new_n391_), .A3(new_n354_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n389_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT20), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n303_), .A2(new_n305_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT88), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n301_), .A2(new_n306_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT88), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n303_), .A2(new_n305_), .A3(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n396_), .A2(new_n398_), .A3(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n326_), .A2(new_n327_), .A3(new_n321_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(new_n402_), .A3(new_n308_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n332_), .A2(new_n331_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n318_), .A2(new_n340_), .A3(new_n341_), .A4(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n394_), .B1(new_n406_), .B2(new_n371_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n375_), .A2(new_n342_), .A3(new_n325_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G226gat), .A2(G233gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n409_), .A2(new_n413_), .ZN(new_n414_));
  XOR2_X1   g213(.A(G8gat), .B(G36gat), .Z(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT18), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G64gat), .B(G92gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n343_), .A2(new_n371_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n375_), .A2(new_n403_), .A3(new_n405_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(KEYINPUT20), .A3(new_n421_), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n414_), .B(new_n419_), .C1(new_n413_), .C2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n409_), .A2(new_n412_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n420_), .A2(new_n421_), .A3(KEYINPUT20), .A4(new_n413_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n424_), .A2(new_n418_), .A3(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n423_), .A2(KEYINPUT27), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT27), .ZN(new_n429_));
  INV_X1    g228(.A(new_n425_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n413_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n431_));
  NOR3_X1   g230(.A1(new_n430_), .A2(new_n419_), .A3(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n418_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n429_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT93), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n419_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n426_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT93), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(new_n429_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n428_), .B1(new_n435_), .B2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n351_), .B1(new_n393_), .B2(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n438_), .B1(new_n437_), .B2(new_n429_), .ZN(new_n442_));
  AOI211_X1 g241(.A(KEYINPUT93), .B(KEYINPUT27), .C1(new_n436_), .C2(new_n426_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n427_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  AOI211_X1 g243(.A(KEYINPUT94), .B(new_n444_), .C1(new_n389_), .C2(new_n392_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n294_), .B(new_n350_), .C1(new_n441_), .C2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n350_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n292_), .A2(new_n285_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT92), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n440_), .A2(new_n450_), .A3(new_n288_), .A4(new_n290_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n393_), .A2(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n414_), .B1(new_n422_), .B2(new_n413_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n424_), .A2(new_n425_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n418_), .A2(KEYINPUT32), .ZN(new_n455_));
  MUX2_X1   g254(.A(new_n453_), .B(new_n454_), .S(new_n455_), .Z(new_n456_));
  OAI21_X1  g255(.A(new_n456_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT33), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n290_), .A2(new_n458_), .ZN(new_n459_));
  OAI211_X1 g258(.A(KEYINPUT33), .B(new_n284_), .C1(new_n289_), .C2(new_n286_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n437_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n277_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n276_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n285_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .A4(new_n464_), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n457_), .A2(new_n465_), .B1(new_n392_), .B2(new_n389_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n447_), .B1(new_n452_), .B2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n238_), .B1(new_n446_), .B2(new_n467_), .ZN(new_n468_));
  XOR2_X1   g267(.A(G85gat), .B(G92gat), .Z(new_n469_));
  INV_X1    g268(.A(KEYINPUT9), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT65), .ZN(new_n471_));
  OR2_X1    g270(.A1(new_n470_), .A2(KEYINPUT65), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n469_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(KEYINPUT10), .B(G99gat), .Z(new_n474_));
  INV_X1    g273(.A(G106gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n470_), .A2(KEYINPUT65), .A3(G85gat), .A4(G92gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G99gat), .A2(G106gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT6), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n473_), .A2(new_n476_), .A3(new_n477_), .A4(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT7), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT66), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(KEYINPUT66), .ZN(new_n483_));
  INV_X1    g282(.A(G99gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n475_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n482_), .B1(new_n483_), .B2(new_n485_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n479_), .B(new_n486_), .C1(new_n485_), .C2(new_n482_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT67), .ZN(new_n488_));
  AOI21_X1  g287(.A(KEYINPUT8), .B1(new_n469_), .B2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n469_), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n489_), .B1(new_n487_), .B2(new_n469_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n480_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G232gat), .A2(G233gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT34), .ZN(new_n495_));
  OAI22_X1  g294(.A1(new_n493_), .A2(new_n225_), .B1(KEYINPUT35), .B2(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n496_), .B1(new_n219_), .B2(new_n493_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(KEYINPUT35), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G190gat), .B(G218gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G134gat), .B(G162gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n502_), .B(KEYINPUT36), .Z(new_n503_));
  NAND2_X1  g302(.A1(new_n499_), .A2(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n502_), .A2(KEYINPUT36), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n504_), .B1(new_n505_), .B2(new_n499_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT97), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT12), .ZN(new_n509_));
  INV_X1    g308(.A(new_n480_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n487_), .A2(new_n469_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n489_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n510_), .B1(new_n513_), .B2(new_n490_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G57gat), .B(G64gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT11), .ZN(new_n516_));
  XOR2_X1   g315(.A(G71gat), .B(G78gat), .Z(new_n517_));
  OR2_X1    g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n515_), .A2(KEYINPUT11), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n516_), .A2(new_n517_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n518_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n509_), .B1(new_n514_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT69), .ZN(new_n523_));
  INV_X1    g322(.A(new_n521_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n493_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT69), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n525_), .A2(new_n526_), .A3(new_n509_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n523_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n493_), .A2(KEYINPUT12), .A3(new_n524_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT68), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT68), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n493_), .A2(new_n531_), .A3(KEYINPUT12), .A4(new_n524_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G230gat), .A2(G233gat), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n534_), .B(KEYINPUT64), .Z(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n514_), .A2(new_n521_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n528_), .A2(new_n533_), .A3(new_n536_), .A4(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n525_), .A2(new_n537_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(new_n535_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(G120gat), .B(G148gat), .Z(new_n542_));
  XNOR2_X1  g341(.A(G176gat), .B(G204gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n544_), .B(new_n545_), .Z(new_n546_));
  NAND2_X1  g345(.A1(new_n541_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n546_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n538_), .A2(new_n540_), .A3(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n550_), .A2(KEYINPUT13), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(KEYINPUT13), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G231gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n521_), .B(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(new_n218_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G127gat), .B(G155gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G183gat), .B(G211gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XOR2_X1   g359(.A(KEYINPUT73), .B(KEYINPUT16), .Z(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(KEYINPUT17), .B1(new_n557_), .B2(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n562_), .B1(new_n557_), .B2(KEYINPUT74), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n508_), .A2(new_n554_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n468_), .A2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(G1gat), .B1(new_n568_), .B2(new_n294_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT95), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n468_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n468_), .A2(new_n570_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n553_), .B(KEYINPUT71), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n506_), .B(KEYINPUT37), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(new_n565_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n573_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT96), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT96), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n573_), .A2(new_n581_), .A3(new_n578_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n294_), .A2(G1gat), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n580_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n584_), .A2(KEYINPUT38), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(KEYINPUT38), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n569_), .B1(new_n585_), .B2(new_n586_), .ZN(G1324gat));
  NOR2_X1   g386(.A1(new_n440_), .A2(G8gat), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n580_), .A2(new_n582_), .A3(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(G8gat), .B1(new_n568_), .B2(new_n440_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT39), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT40), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n589_), .A2(new_n591_), .A3(KEYINPUT40), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(G1325gat));
  INV_X1    g395(.A(new_n579_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n597_), .A2(new_n206_), .A3(new_n350_), .ZN(new_n598_));
  OAI21_X1  g397(.A(G15gat), .B1(new_n568_), .B2(new_n447_), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n599_), .A2(KEYINPUT41), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(KEYINPUT41), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n598_), .A2(new_n600_), .A3(new_n601_), .ZN(G1326gat));
  OAI21_X1  g401(.A(G22gat), .B1(new_n568_), .B2(new_n393_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT42), .ZN(new_n604_));
  INV_X1    g403(.A(new_n393_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(new_n204_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n604_), .B1(new_n579_), .B2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT98), .ZN(G1327gat));
  NOR2_X1   g407(.A1(new_n506_), .A2(new_n565_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n553_), .A2(new_n609_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n573_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n294_), .ZN(new_n612_));
  AOI21_X1  g411(.A(G29gat), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n554_), .A2(new_n238_), .A3(new_n565_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT43), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n446_), .A2(new_n467_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n506_), .B(KEYINPUT37), .Z(new_n617_));
  AOI21_X1  g416(.A(new_n615_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  AOI211_X1 g417(.A(KEYINPUT43), .B(new_n576_), .C1(new_n446_), .C2(new_n467_), .ZN(new_n619_));
  OAI211_X1 g418(.A(KEYINPUT44), .B(new_n614_), .C1(new_n618_), .C2(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n614_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT44), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n623_), .A2(G29gat), .A3(new_n612_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n613_), .B1(new_n620_), .B2(new_n624_), .ZN(G1328gat));
  NOR2_X1   g424(.A1(new_n440_), .A2(G36gat), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n571_), .A2(new_n572_), .A3(new_n610_), .A4(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT45), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT99), .ZN(new_n629_));
  INV_X1    g428(.A(G36gat), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n440_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n631_));
  AOI211_X1 g430(.A(new_n629_), .B(new_n630_), .C1(new_n631_), .C2(new_n620_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n623_), .A2(new_n444_), .A3(new_n620_), .ZN(new_n633_));
  AOI21_X1  g432(.A(KEYINPUT99), .B1(new_n633_), .B2(G36gat), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n628_), .B1(new_n632_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT46), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  OAI211_X1 g436(.A(KEYINPUT46), .B(new_n628_), .C1(new_n632_), .C2(new_n634_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(G1329gat));
  NAND2_X1  g438(.A1(new_n611_), .A2(new_n350_), .ZN(new_n640_));
  INV_X1    g439(.A(G43gat), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n623_), .A2(G43gat), .A3(new_n350_), .A4(new_n620_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(KEYINPUT100), .B(KEYINPUT47), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n642_), .A2(new_n643_), .A3(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n644_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n645_), .A2(new_n646_), .ZN(G1330gat));
  AOI21_X1  g446(.A(G50gat), .B1(new_n611_), .B2(new_n605_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n623_), .A2(G50gat), .A3(new_n605_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n620_), .B2(new_n649_), .ZN(G1331gat));
  AND3_X1   g449(.A1(new_n575_), .A2(new_n616_), .A3(new_n238_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n651_), .A2(new_n565_), .A3(new_n507_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT101), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(G57gat), .B1(new_n655_), .B2(new_n294_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n554_), .A2(new_n238_), .ZN(new_n657_));
  AOI211_X1 g456(.A(new_n577_), .B(new_n657_), .C1(new_n446_), .C2(new_n467_), .ZN(new_n658_));
  INV_X1    g457(.A(G57gat), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n658_), .A2(new_n659_), .A3(new_n612_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n656_), .A2(new_n660_), .ZN(G1332gat));
  OAI21_X1  g460(.A(G64gat), .B1(new_n655_), .B2(new_n440_), .ZN(new_n662_));
  XOR2_X1   g461(.A(KEYINPUT102), .B(KEYINPUT48), .Z(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n663_), .ZN(new_n665_));
  OAI211_X1 g464(.A(G64gat), .B(new_n665_), .C1(new_n655_), .C2(new_n440_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n440_), .A2(G64gat), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT103), .Z(new_n668_));
  NAND2_X1  g467(.A1(new_n658_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n664_), .A2(new_n666_), .A3(new_n669_), .ZN(G1333gat));
  NAND2_X1  g469(.A1(new_n654_), .A2(new_n350_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(G71gat), .ZN(new_n672_));
  XOR2_X1   g471(.A(KEYINPUT104), .B(KEYINPUT49), .Z(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n673_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n671_), .A2(G71gat), .A3(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(G71gat), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n658_), .A2(new_n677_), .A3(new_n350_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n674_), .A2(new_n676_), .A3(new_n678_), .ZN(G1334gat));
  INV_X1    g478(.A(G78gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n658_), .A2(new_n680_), .A3(new_n605_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT50), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n654_), .A2(new_n605_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n682_), .B1(new_n683_), .B2(G78gat), .ZN(new_n684_));
  AOI211_X1 g483(.A(KEYINPUT50), .B(new_n680_), .C1(new_n654_), .C2(new_n605_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n681_), .B1(new_n684_), .B2(new_n685_), .ZN(G1335gat));
  NOR2_X1   g485(.A1(new_n657_), .A2(new_n565_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n687_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n688_), .A2(KEYINPUT105), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(KEYINPUT105), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(G85gat), .B1(new_n691_), .B2(new_n294_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n651_), .A2(new_n609_), .ZN(new_n693_));
  INV_X1    g492(.A(G85gat), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(new_n694_), .A3(new_n612_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n692_), .A2(new_n695_), .ZN(G1336gat));
  OAI21_X1  g495(.A(G92gat), .B1(new_n691_), .B2(new_n440_), .ZN(new_n697_));
  INV_X1    g496(.A(G92gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n693_), .A2(new_n698_), .A3(new_n444_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(G1337gat));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n701_), .A2(KEYINPUT51), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(KEYINPUT51), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n688_), .B(KEYINPUT105), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n484_), .B1(new_n704_), .B2(new_n350_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n693_), .A2(new_n350_), .A3(new_n474_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n702_), .B(new_n703_), .C1(new_n705_), .C2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(G99gat), .B1(new_n691_), .B2(new_n447_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n709_), .A2(new_n701_), .A3(KEYINPUT51), .A4(new_n706_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n708_), .A2(new_n710_), .ZN(G1338gat));
  NAND3_X1  g510(.A1(new_n693_), .A2(new_n475_), .A3(new_n605_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT52), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n605_), .B(new_n687_), .C1(new_n618_), .C2(new_n619_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n714_), .B2(G106gat), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n714_), .A2(new_n713_), .A3(G106gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n718_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n712_), .B1(new_n717_), .B2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(KEYINPUT53), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT53), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n722_), .B(new_n712_), .C1(new_n717_), .C2(new_n719_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(G1339gat));
  INV_X1    g523(.A(G113gat), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n441_), .A2(new_n445_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n726_), .A2(new_n447_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n237_), .A2(new_n549_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT109), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n237_), .A2(new_n549_), .A3(KEYINPUT109), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT55), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n538_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n528_), .A2(new_n533_), .A3(new_n537_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(new_n535_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n734_), .B1(new_n538_), .B2(new_n733_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n546_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT56), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  OAI211_X1 g541(.A(KEYINPUT56), .B(new_n546_), .C1(new_n738_), .C2(new_n739_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n732_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n227_), .A2(new_n226_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n235_), .B1(new_n745_), .B2(new_n221_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n216_), .A2(new_n220_), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n747_), .A2(KEYINPUT111), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(KEYINPUT111), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n746_), .B1(new_n750_), .B2(new_n221_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT112), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT112), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n753_), .B(new_n746_), .C1(new_n750_), .C2(new_n221_), .ZN(new_n754_));
  AND4_X1   g553(.A1(new_n236_), .A2(new_n550_), .A3(new_n752_), .A4(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n506_), .B1(new_n744_), .B2(new_n755_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT57), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n752_), .A2(new_n549_), .A3(new_n754_), .A4(new_n236_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n617_), .B1(new_n759_), .B2(KEYINPUT58), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT113), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT113), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n617_), .B(new_n762_), .C1(new_n759_), .C2(KEYINPUT58), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n759_), .A2(KEYINPUT58), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n761_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n565_), .B1(new_n757_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n565_), .A2(new_n238_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT108), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n617_), .A2(new_n554_), .A3(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT54), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n612_), .B(new_n727_), .C1(new_n766_), .C2(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n725_), .B1(new_n771_), .B2(new_n238_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT114), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n774_), .B(new_n725_), .C1(new_n771_), .C2(new_n238_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT115), .B1(new_n771_), .B2(KEYINPUT59), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n771_), .A2(KEYINPUT115), .A3(KEYINPUT59), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT59), .ZN(new_n780_));
  INV_X1    g579(.A(new_n771_), .ZN(new_n781_));
  AOI22_X1  g580(.A1(new_n778_), .A2(new_n779_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n238_), .A2(new_n725_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n776_), .B1(new_n782_), .B2(new_n783_), .ZN(G1340gat));
  NAND2_X1  g583(.A1(new_n781_), .A2(new_n780_), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n771_), .A2(KEYINPUT115), .A3(KEYINPUT59), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n575_), .B(new_n785_), .C1(new_n786_), .C2(new_n777_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(G120gat), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT60), .ZN(new_n789_));
  INV_X1    g588(.A(G120gat), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n554_), .A2(new_n789_), .A3(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n791_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n781_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n788_), .A2(new_n793_), .ZN(G1341gat));
  AOI21_X1  g593(.A(G127gat), .B1(new_n781_), .B2(new_n565_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT116), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n565_), .A2(new_n796_), .A3(G127gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n797_), .B1(new_n796_), .B2(G127gat), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n795_), .B1(new_n782_), .B2(new_n798_), .ZN(G1342gat));
  INV_X1    g598(.A(G134gat), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n800_), .B1(new_n771_), .B2(new_n507_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT117), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  OAI211_X1 g602(.A(KEYINPUT117), .B(new_n800_), .C1(new_n771_), .C2(new_n507_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n576_), .A2(new_n800_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n782_), .B2(new_n806_), .ZN(G1343gat));
  OR2_X1    g606(.A1(new_n766_), .A2(new_n770_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n393_), .A2(new_n350_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n810_), .A2(new_n444_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n808_), .A2(new_n612_), .A3(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n812_), .A2(new_n238_), .ZN(new_n813_));
  XOR2_X1   g612(.A(KEYINPUT118), .B(G141gat), .Z(new_n814_));
  XNOR2_X1  g613(.A(new_n813_), .B(new_n814_), .ZN(G1344gat));
  NOR2_X1   g614(.A1(new_n812_), .A2(new_n574_), .ZN(new_n816_));
  XOR2_X1   g615(.A(KEYINPUT119), .B(G148gat), .Z(new_n817_));
  XNOR2_X1  g616(.A(new_n816_), .B(new_n817_), .ZN(G1345gat));
  NOR2_X1   g617(.A1(new_n812_), .A2(new_n566_), .ZN(new_n819_));
  XOR2_X1   g618(.A(KEYINPUT61), .B(G155gat), .Z(new_n820_));
  XNOR2_X1  g619(.A(new_n819_), .B(new_n820_), .ZN(G1346gat));
  INV_X1    g620(.A(G162gat), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n822_), .B1(new_n812_), .B2(new_n507_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT120), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  OAI211_X1 g624(.A(KEYINPUT120), .B(new_n822_), .C1(new_n812_), .C2(new_n507_), .ZN(new_n826_));
  OR3_X1    g625(.A1(new_n812_), .A2(new_n822_), .A3(new_n576_), .ZN(new_n827_));
  AND3_X1   g626(.A1(new_n825_), .A2(new_n826_), .A3(new_n827_), .ZN(G1347gat));
  NOR4_X1   g627(.A1(new_n605_), .A2(new_n447_), .A3(new_n612_), .A4(new_n440_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n808_), .A2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(G169gat), .B1(new_n830_), .B2(new_n238_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(KEYINPUT121), .B(KEYINPUT62), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n832_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n830_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n835_), .A2(new_n396_), .A3(new_n400_), .A4(new_n237_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n833_), .A2(new_n834_), .A3(new_n836_), .ZN(G1348gat));
  AOI21_X1  g636(.A(new_n397_), .B1(new_n835_), .B2(new_n554_), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n830_), .A2(new_n334_), .A3(new_n574_), .ZN(new_n839_));
  OAI21_X1  g638(.A(KEYINPUT122), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n835_), .A2(G176gat), .A3(new_n575_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT122), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n398_), .B1(new_n830_), .B2(new_n553_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n841_), .A2(new_n842_), .A3(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n840_), .A2(new_n844_), .ZN(G1349gat));
  AOI21_X1  g644(.A(new_n319_), .B1(new_n835_), .B2(new_n565_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n331_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n830_), .A2(new_n847_), .A3(new_n566_), .ZN(new_n848_));
  OAI21_X1  g647(.A(KEYINPUT123), .B1(new_n846_), .B2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n835_), .A2(new_n331_), .A3(new_n565_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT123), .ZN(new_n851_));
  OAI21_X1  g650(.A(G183gat), .B1(new_n830_), .B2(new_n566_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n850_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n849_), .A2(new_n853_), .ZN(G1350gat));
  INV_X1    g653(.A(KEYINPUT124), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n320_), .B1(new_n835_), .B2(new_n617_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n332_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n830_), .A2(new_n857_), .A3(new_n507_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n855_), .B1(new_n856_), .B2(new_n858_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n835_), .A2(new_n332_), .A3(new_n508_), .ZN(new_n860_));
  OAI21_X1  g659(.A(G190gat), .B1(new_n830_), .B2(new_n576_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(KEYINPUT124), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n859_), .A2(new_n862_), .ZN(G1351gat));
  INV_X1    g662(.A(KEYINPUT126), .ZN(new_n864_));
  INV_X1    g663(.A(G197gat), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n810_), .A2(new_n612_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n866_), .A2(KEYINPUT125), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(KEYINPUT125), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n867_), .A2(new_n868_), .A3(new_n440_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n808_), .A2(new_n869_), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n864_), .B(new_n865_), .C1(new_n870_), .C2(new_n238_), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n808_), .A2(new_n869_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n237_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n871_), .B1(new_n873_), .B2(new_n865_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n864_), .B1(new_n873_), .B2(new_n865_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n874_), .A2(new_n875_), .ZN(G1352gat));
  AOI21_X1  g675(.A(new_n574_), .B1(KEYINPUT127), .B2(G204gat), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n872_), .A2(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n879_));
  XOR2_X1   g678(.A(new_n878_), .B(new_n879_), .Z(G1353gat));
  NOR2_X1   g679(.A1(new_n870_), .A2(new_n566_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n882_));
  AND2_X1   g681(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n881_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(new_n881_), .B2(new_n882_), .ZN(G1354gat));
  NAND3_X1  g684(.A1(new_n872_), .A2(new_n365_), .A3(new_n508_), .ZN(new_n886_));
  OAI21_X1  g685(.A(G218gat), .B1(new_n870_), .B2(new_n576_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1355gat));
endmodule


