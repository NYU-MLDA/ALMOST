//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 0 1 1 0 1 1 1 0 1 0 0 0 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n919_, new_n920_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n952_, new_n953_,
    new_n954_, new_n956_, new_n957_, new_n958_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n968_,
    new_n969_, new_n970_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n977_, new_n978_, new_n979_;
  INV_X1    g000(.A(KEYINPUT15), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G29gat), .B(G36gat), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n204_), .A2(KEYINPUT71), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(KEYINPUT71), .ZN(new_n206_));
  AOI21_X1  g005(.A(new_n203_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n204_), .A2(KEYINPUT71), .ZN(new_n208_));
  INV_X1    g007(.A(G36gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G29gat), .ZN(new_n210_));
  INV_X1    g009(.A(G29gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G36gat), .ZN(new_n212_));
  AND3_X1   g011(.A1(new_n210_), .A2(new_n212_), .A3(KEYINPUT71), .ZN(new_n213_));
  INV_X1    g012(.A(new_n203_), .ZN(new_n214_));
  NOR3_X1   g013(.A1(new_n208_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n202_), .B1(new_n207_), .B2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n205_), .A2(new_n206_), .A3(new_n203_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n214_), .B1(new_n208_), .B2(new_n213_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(new_n218_), .A3(KEYINPUT15), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G15gat), .B(G22gat), .ZN(new_n221_));
  INV_X1    g020(.A(G1gat), .ZN(new_n222_));
  INV_X1    g021(.A(G8gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT14), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n221_), .A2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G1gat), .B(G8gat), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n226_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n220_), .A2(new_n229_), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n217_), .A2(new_n227_), .A3(new_n218_), .A4(new_n228_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G229gat), .A2(G233gat), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n230_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n217_), .A2(new_n218_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(new_n229_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(new_n231_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n232_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n234_), .A2(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(G113gat), .B(G141gat), .Z(new_n241_));
  XOR2_X1   g040(.A(G169gat), .B(G197gat), .Z(new_n242_));
  XOR2_X1   g041(.A(new_n241_), .B(new_n242_), .Z(new_n243_));
  OR2_X1    g042(.A1(new_n240_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n234_), .A2(new_n239_), .A3(new_n243_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT79), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n234_), .A2(KEYINPUT79), .A3(new_n239_), .A4(new_n243_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n244_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NOR3_X1   g050(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G169gat), .A2(G176gat), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n252_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G183gat), .A2(G190gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT23), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n260_));
  XOR2_X1   g059(.A(KEYINPUT81), .B(G190gat), .Z(new_n261_));
  AOI21_X1  g060(.A(new_n260_), .B1(new_n261_), .B2(KEYINPUT26), .ZN(new_n262_));
  NOR2_X1   g061(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n263_));
  XOR2_X1   g062(.A(KEYINPUT80), .B(G183gat), .Z(new_n264_));
  AOI21_X1  g063(.A(new_n263_), .B1(new_n264_), .B2(KEYINPUT25), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n259_), .B1(new_n262_), .B2(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n258_), .B1(new_n261_), .B2(new_n264_), .ZN(new_n267_));
  INV_X1    g066(.A(G176gat), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT22), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT82), .B1(new_n269_), .B2(G169gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT22), .B(G169gat), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n268_), .B(new_n270_), .C1(new_n271_), .C2(KEYINPUT82), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n267_), .A2(new_n255_), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n266_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G71gat), .B(G99gat), .ZN(new_n275_));
  XOR2_X1   g074(.A(new_n275_), .B(G43gat), .Z(new_n276_));
  XNOR2_X1  g075(.A(new_n274_), .B(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G227gat), .A2(G233gat), .ZN(new_n278_));
  INV_X1    g077(.A(G15gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT30), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT31), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n277_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n277_), .A2(new_n283_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT83), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(G127gat), .B(G134gat), .Z(new_n290_));
  XOR2_X1   g089(.A(G113gat), .B(G120gat), .Z(new_n291_));
  XOR2_X1   g090(.A(new_n290_), .B(new_n291_), .Z(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n286_), .A2(KEYINPUT83), .ZN(new_n294_));
  OR3_X1    g093(.A1(new_n289_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n293_), .B1(new_n289_), .B2(new_n294_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT100), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299_));
  INV_X1    g098(.A(G155gat), .ZN(new_n300_));
  INV_X1    g099(.A(G162gat), .ZN(new_n301_));
  AND3_X1   g100(.A1(new_n300_), .A2(new_n301_), .A3(KEYINPUT85), .ZN(new_n302_));
  AOI21_X1  g101(.A(KEYINPUT85), .B1(new_n300_), .B2(new_n301_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n299_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT87), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G141gat), .A2(G148gat), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT2), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT3), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n309_), .B1(G141gat), .B2(G148gat), .ZN(new_n310_));
  INV_X1    g109(.A(G141gat), .ZN(new_n311_));
  INV_X1    g110(.A(G148gat), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n311_), .A2(new_n312_), .A3(KEYINPUT3), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n308_), .B1(new_n310_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n306_), .A2(KEYINPUT84), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT84), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n316_), .A2(G141gat), .A3(G148gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n317_), .A3(new_n307_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n314_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT87), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n320_), .B(new_n299_), .C1(new_n302_), .C2(new_n303_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n305_), .A2(new_n319_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n315_), .A2(new_n317_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n323_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n299_), .A2(KEYINPUT1), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT86), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  OAI22_X1  g126(.A1(new_n302_), .A2(new_n303_), .B1(KEYINPUT1), .B2(new_n299_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n324_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n322_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT88), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT88), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n322_), .A2(new_n332_), .A3(new_n329_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n331_), .A2(KEYINPUT29), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(G204gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(KEYINPUT92), .A3(G197gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(G197gat), .ZN(new_n337_));
  INV_X1    g136(.A(G197gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(G204gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  OAI211_X1 g139(.A(KEYINPUT21), .B(new_n336_), .C1(new_n340_), .C2(KEYINPUT92), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT21), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n337_), .A2(new_n339_), .A3(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G211gat), .B(G218gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n341_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n340_), .A2(KEYINPUT21), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n346_), .A2(new_n344_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(G233gat), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n350_), .A2(KEYINPUT91), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(KEYINPUT91), .ZN(new_n352_));
  NOR2_X1   g151(.A1(KEYINPUT90), .A2(G228gat), .ZN(new_n353_));
  AND2_X1   g152(.A1(KEYINPUT90), .A2(G228gat), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n351_), .B(new_n352_), .C1(new_n353_), .C2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n349_), .A2(new_n356_), .ZN(new_n357_));
  AOI22_X1  g156(.A1(KEYINPUT87), .A2(new_n304_), .B1(new_n314_), .B2(new_n318_), .ZN(new_n358_));
  OR2_X1    g157(.A1(new_n299_), .A2(KEYINPUT1), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n325_), .A2(KEYINPUT86), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n326_), .B1(new_n299_), .B2(KEYINPUT1), .ZN(new_n361_));
  OAI221_X1 g160(.A(new_n359_), .B1(new_n302_), .B2(new_n303_), .C1(new_n360_), .C2(new_n361_), .ZN(new_n362_));
  AOI22_X1  g161(.A1(new_n358_), .A2(new_n321_), .B1(new_n362_), .B2(new_n324_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT29), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT93), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n345_), .A2(new_n365_), .A3(new_n347_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n365_), .B1(new_n345_), .B2(new_n347_), .ZN(new_n367_));
  OAI22_X1  g166(.A1(new_n363_), .A2(new_n364_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  AOI22_X1  g167(.A1(new_n334_), .A2(new_n357_), .B1(new_n368_), .B2(new_n356_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G78gat), .B(G106gat), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT94), .B1(new_n369_), .B2(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n366_), .A2(new_n367_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n364_), .B1(new_n322_), .B2(new_n329_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n356_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n322_), .A2(new_n332_), .A3(new_n329_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n332_), .B1(new_n322_), .B2(new_n329_), .ZN(new_n377_));
  NOR3_X1   g176(.A1(new_n376_), .A2(new_n377_), .A3(new_n364_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n357_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n375_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT94), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n380_), .A2(new_n381_), .A3(new_n370_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n372_), .A2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G22gat), .B(G50gat), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT28), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n331_), .A2(new_n333_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n386_), .B1(new_n387_), .B2(new_n364_), .ZN(new_n388_));
  AOI211_X1 g187(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n331_), .C2(new_n333_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n385_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n376_), .A2(new_n377_), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT28), .B1(new_n391_), .B2(KEYINPUT29), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n387_), .A2(new_n386_), .A3(new_n364_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n392_), .A2(new_n393_), .A3(new_n384_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n375_), .B(new_n371_), .C1(new_n378_), .C2(new_n379_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n390_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n383_), .A2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(KEYINPUT89), .B1(new_n390_), .B2(new_n394_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n390_), .A2(KEYINPUT89), .A3(new_n394_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n380_), .A2(new_n370_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n395_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n397_), .B1(new_n399_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT27), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n349_), .A2(new_n266_), .A3(new_n273_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n258_), .B1(G183gat), .B2(G190gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n271_), .A2(new_n268_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n255_), .B(KEYINPUT97), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT25), .B(G183gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT26), .B(G190gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n259_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT96), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n259_), .A2(KEYINPUT96), .A3(new_n414_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n411_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  OAI211_X1 g218(.A(KEYINPUT20), .B(new_n406_), .C1(new_n419_), .C2(new_n349_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G226gat), .A2(G233gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n420_), .A2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G8gat), .B(G36gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT18), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G64gat), .B(G92gat), .ZN(new_n428_));
  XOR2_X1   g227(.A(new_n427_), .B(new_n428_), .Z(new_n429_));
  NAND2_X1  g228(.A1(new_n419_), .A2(new_n349_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT20), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n431_), .B1(new_n274_), .B2(new_n348_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n423_), .A3(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n425_), .A2(new_n429_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n429_), .B1(new_n425_), .B2(new_n433_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n405_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT4), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n331_), .A2(new_n333_), .A3(new_n292_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n330_), .A2(new_n292_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n438_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(KEYINPUT4), .B1(new_n391_), .B2(new_n292_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G225gat), .A2(G233gat), .ZN(new_n444_));
  NOR3_X1   g243(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n444_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n447_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G1gat), .B(G29gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(G85gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT0), .B(G57gat), .ZN(new_n452_));
  XOR2_X1   g251(.A(new_n451_), .B(new_n452_), .Z(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n446_), .A2(new_n449_), .A3(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n453_), .B1(new_n445_), .B2(new_n448_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n429_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n420_), .A2(new_n424_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n373_), .A2(new_n410_), .A3(new_n415_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n423_), .B1(new_n459_), .B2(new_n432_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n457_), .B1(new_n458_), .B2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(KEYINPUT27), .A3(new_n434_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n437_), .A2(new_n455_), .A3(new_n456_), .A4(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n298_), .B1(new_n404_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n437_), .A2(new_n462_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n400_), .A2(new_n402_), .ZN(new_n467_));
  OAI22_X1  g266(.A1(new_n467_), .A2(new_n398_), .B1(new_n396_), .B2(new_n383_), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n455_), .A2(new_n456_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n466_), .A2(new_n468_), .A3(new_n469_), .A4(KEYINPUT100), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n464_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT98), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n456_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT33), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT33), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n456_), .A2(new_n472_), .A3(new_n475_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n417_), .A2(new_n418_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n348_), .B1(new_n477_), .B2(new_n411_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n274_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n431_), .B1(new_n479_), .B2(new_n349_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n423_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n430_), .A2(new_n423_), .A3(new_n432_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n457_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(new_n434_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n444_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n485_), .A2(KEYINPUT99), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n439_), .A2(new_n441_), .A3(new_n447_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(new_n454_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n488_), .B1(new_n485_), .B2(KEYINPUT99), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n484_), .B1(new_n486_), .B2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n474_), .A2(new_n476_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n455_), .A2(new_n456_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n429_), .A2(KEYINPUT32), .ZN(new_n493_));
  NOR3_X1   g292(.A1(new_n481_), .A2(new_n482_), .A3(new_n493_), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n458_), .A2(new_n460_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n494_), .B1(new_n495_), .B2(new_n493_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n492_), .A2(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n468_), .B1(new_n491_), .B2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n297_), .B1(new_n471_), .B2(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n297_), .A2(new_n492_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(new_n404_), .A3(new_n466_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n251_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n502_));
  AND2_X1   g301(.A1(G230gat), .A2(G233gat), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT65), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT9), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT9), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(KEYINPUT65), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n505_), .A2(new_n507_), .A3(G85gat), .A4(G92gat), .ZN(new_n508_));
  INV_X1    g307(.A(G85gat), .ZN(new_n509_));
  INV_X1    g308(.A(G92gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G85gat), .A2(G92gat), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n511_), .A2(new_n504_), .A3(KEYINPUT9), .A4(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G99gat), .A2(G106gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT6), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT6), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n516_), .A2(G99gat), .A3(G106gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n508_), .A2(new_n513_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(G106gat), .ZN(new_n520_));
  OR2_X1    g319(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT64), .ZN(new_n522_));
  NAND2_X1  g321(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n521_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n522_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n520_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n519_), .A2(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT7), .ZN(new_n529_));
  INV_X1    g328(.A(G99gat), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(new_n530_), .A3(new_n520_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n518_), .A2(new_n528_), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT8), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n511_), .A2(new_n512_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n532_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n533_), .B1(new_n532_), .B2(new_n534_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n527_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G71gat), .B(G78gat), .ZN(new_n539_));
  INV_X1    g338(.A(G64gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(G57gat), .ZN(new_n541_));
  INV_X1    g340(.A(G57gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(G64gat), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n539_), .A2(KEYINPUT11), .A3(new_n541_), .A4(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n541_), .A2(new_n543_), .A3(KEYINPUT11), .ZN(new_n545_));
  INV_X1    g344(.A(G78gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(G71gat), .ZN(new_n547_));
  INV_X1    g346(.A(G71gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(G78gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n545_), .A2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(KEYINPUT11), .B1(new_n541_), .B2(new_n543_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n544_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT66), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT66), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n544_), .B(new_n555_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n538_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(KEYINPUT67), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n538_), .A2(new_n557_), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n561_), .A2(KEYINPUT67), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n503_), .B(new_n560_), .C1(new_n562_), .C2(new_n559_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT12), .ZN(new_n564_));
  INV_X1    g363(.A(new_n556_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT11), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n542_), .A2(G64gat), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n540_), .A2(G57gat), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n566_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n569_), .A2(new_n545_), .A3(new_n550_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n555_), .B1(new_n570_), .B2(new_n544_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n565_), .A2(new_n571_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n515_), .A2(new_n517_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n531_), .A2(new_n528_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n534_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(KEYINPUT8), .ZN(new_n576_));
  AOI22_X1  g375(.A1(new_n576_), .A2(new_n535_), .B1(new_n526_), .B2(new_n519_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n564_), .B1(new_n572_), .B2(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n503_), .B1(new_n572_), .B2(new_n577_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT68), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n570_), .A2(KEYINPUT12), .A3(new_n544_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n580_), .B1(new_n577_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n581_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n538_), .A2(KEYINPUT68), .A3(new_n583_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n578_), .A2(new_n579_), .A3(new_n582_), .A4(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n563_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G120gat), .B(G148gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT5), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G176gat), .B(G204gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT69), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n586_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n563_), .A2(new_n585_), .A3(new_n590_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n593_), .A2(KEYINPUT70), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT13), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT70), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n586_), .A2(new_n597_), .A3(new_n592_), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n595_), .A2(new_n596_), .A3(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n596_), .B1(new_n595_), .B2(new_n598_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G127gat), .B(G155gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT16), .ZN(new_n603_));
  XOR2_X1   g402(.A(G183gat), .B(G211gat), .Z(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT17), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT78), .Z(new_n609_));
  XNOR2_X1  g408(.A(new_n229_), .B(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n607_), .B1(new_n610_), .B2(new_n557_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n611_), .B1(new_n610_), .B2(new_n557_), .ZN(new_n612_));
  AOI211_X1 g411(.A(new_n606_), .B(new_n605_), .C1(new_n610_), .C2(new_n553_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n613_), .B1(new_n553_), .B2(new_n610_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G190gat), .B(G218gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT73), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT74), .ZN(new_n619_));
  XOR2_X1   g418(.A(G134gat), .B(G162gat), .Z(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT36), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n235_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT35), .ZN(new_n625_));
  NAND2_X1  g424(.A1(G232gat), .A2(G233gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT34), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  AOI22_X1  g427(.A1(new_n577_), .A2(new_n624_), .B1(new_n625_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT72), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n220_), .A2(new_n630_), .A3(new_n538_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n630_), .B1(new_n220_), .B2(new_n538_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n629_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n628_), .A2(new_n625_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  OAI221_X1 g434(.A(new_n629_), .B1(new_n625_), .B2(new_n628_), .C1(new_n631_), .C2(new_n632_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n623_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(KEYINPUT75), .B(KEYINPUT36), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n621_), .A2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n635_), .A2(new_n636_), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT76), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n635_), .A2(new_n636_), .A3(KEYINPUT76), .A4(new_n639_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n637_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(KEYINPUT77), .A2(KEYINPUT37), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT77), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT37), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n644_), .A2(new_n645_), .A3(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n642_), .A2(new_n643_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n637_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n601_), .A2(new_n616_), .A3(new_n649_), .A4(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n502_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(new_n222_), .A3(new_n492_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT38), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT101), .ZN(new_n661_));
  AOI211_X1 g460(.A(new_n615_), .B(new_n644_), .C1(new_n499_), .C2(new_n501_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n601_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n663_), .A2(new_n251_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n222_), .B1(new_n666_), .B2(new_n492_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n667_), .B1(new_n659_), .B2(new_n658_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n661_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT102), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT102), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n661_), .A2(new_n671_), .A3(new_n668_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(G1324gat));
  OAI21_X1  g472(.A(G8gat), .B1(new_n665_), .B2(new_n466_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT39), .ZN(new_n676_));
  OAI21_X1  g475(.A(KEYINPUT103), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n675_), .A2(new_n678_), .A3(new_n676_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n674_), .A2(new_n680_), .A3(KEYINPUT39), .ZN(new_n681_));
  OAI21_X1  g480(.A(KEYINPUT104), .B1(new_n674_), .B2(KEYINPUT39), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n677_), .A2(new_n679_), .A3(new_n681_), .A4(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n657_), .A2(new_n223_), .A3(new_n465_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT40), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n683_), .A2(KEYINPUT40), .A3(new_n684_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1325gat));
  OAI21_X1  g488(.A(G15gat), .B1(new_n665_), .B2(new_n297_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT41), .Z(new_n691_));
  INV_X1    g490(.A(new_n297_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n657_), .A2(new_n279_), .A3(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1326gat));
  OAI21_X1  g493(.A(G22gat), .B1(new_n665_), .B2(new_n404_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT42), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n404_), .A2(G22gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n696_), .B1(new_n656_), .B2(new_n697_), .ZN(G1327gat));
  AND4_X1   g497(.A1(new_n502_), .A2(new_n615_), .A3(new_n644_), .A4(new_n601_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n492_), .A2(new_n211_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT105), .Z(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n664_), .A2(new_n615_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n499_), .A2(new_n501_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n653_), .A2(new_n649_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT43), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n704_), .A2(new_n708_), .A3(new_n705_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n703_), .B1(new_n707_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n710_), .B(new_n711_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n712_), .A2(new_n492_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n702_), .B1(new_n713_), .B2(new_n211_), .ZN(G1328gat));
  OR2_X1    g513(.A1(new_n710_), .A2(KEYINPUT44), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n710_), .A2(KEYINPUT44), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n715_), .A2(new_n465_), .A3(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(G36gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n699_), .A2(new_n209_), .A3(new_n465_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT45), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n718_), .B(new_n720_), .C1(KEYINPUT106), .C2(KEYINPUT46), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1329gat));
  NAND3_X1  g524(.A1(new_n712_), .A2(G43gat), .A3(new_n692_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n699_), .A2(new_n692_), .ZN(new_n727_));
  XOR2_X1   g526(.A(KEYINPUT107), .B(G43gat), .Z(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n726_), .A2(new_n729_), .A3(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n726_), .B2(new_n729_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1330gat));
  AOI21_X1  g532(.A(G50gat), .B1(new_n699_), .B2(new_n468_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n468_), .A2(G50gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n712_), .B2(new_n735_), .ZN(G1331gat));
  NOR2_X1   g535(.A1(new_n601_), .A2(new_n250_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n662_), .A2(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT109), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(G57gat), .B1(new_n740_), .B2(new_n469_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n704_), .A2(new_n737_), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n742_), .A2(new_n615_), .A3(new_n705_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n743_), .A2(new_n542_), .A3(new_n492_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n741_), .A2(new_n744_), .ZN(G1332gat));
  NAND3_X1  g544(.A1(new_n743_), .A2(new_n540_), .A3(new_n465_), .ZN(new_n746_));
  OAI21_X1  g545(.A(G64gat), .B1(new_n740_), .B2(new_n466_), .ZN(new_n747_));
  XOR2_X1   g546(.A(KEYINPUT110), .B(KEYINPUT48), .Z(new_n748_));
  AND2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n747_), .A2(new_n748_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(G1333gat));
  NAND3_X1  g550(.A1(new_n743_), .A2(new_n548_), .A3(new_n692_), .ZN(new_n752_));
  OAI21_X1  g551(.A(G71gat), .B1(new_n740_), .B2(new_n297_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n753_), .A2(KEYINPUT49), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n753_), .A2(KEYINPUT49), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n752_), .B1(new_n754_), .B2(new_n755_), .ZN(G1334gat));
  NAND3_X1  g555(.A1(new_n743_), .A2(new_n546_), .A3(new_n468_), .ZN(new_n757_));
  OAI21_X1  g556(.A(G78gat), .B1(new_n740_), .B2(new_n404_), .ZN(new_n758_));
  XOR2_X1   g557(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n759_));
  AND2_X1   g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n758_), .A2(new_n759_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n757_), .B1(new_n760_), .B2(new_n761_), .ZN(G1335gat));
  NAND2_X1  g561(.A1(new_n737_), .A2(new_n615_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n763_), .B1(new_n707_), .B2(new_n709_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(G85gat), .B1(new_n765_), .B2(new_n469_), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n742_), .A2(new_n616_), .A3(new_n652_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n767_), .A2(new_n509_), .A3(new_n492_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1336gat));
  OAI21_X1  g568(.A(G92gat), .B1(new_n765_), .B2(new_n466_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n767_), .A2(new_n510_), .A3(new_n465_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(G1337gat));
  OAI21_X1  g571(.A(G99gat), .B1(new_n765_), .B2(new_n297_), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n767_), .B(new_n692_), .C1(new_n524_), .C2(new_n525_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g575(.A1(new_n767_), .A2(new_n520_), .A3(new_n468_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT113), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n601_), .A2(new_n250_), .A3(new_n616_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n708_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n705_), .ZN(new_n781_));
  AOI211_X1 g580(.A(KEYINPUT43), .B(new_n781_), .C1(new_n499_), .C2(new_n501_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n468_), .B(new_n779_), .C1(new_n780_), .C2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(G106gat), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n778_), .B1(new_n784_), .B2(KEYINPUT52), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786_));
  AOI211_X1 g585(.A(KEYINPUT113), .B(new_n786_), .C1(new_n783_), .C2(G106gat), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n785_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n789_), .B1(new_n784_), .B2(KEYINPUT52), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n783_), .A2(KEYINPUT112), .A3(new_n786_), .A4(G106gat), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n777_), .B1(new_n788_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT53), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n795_), .B(new_n777_), .C1(new_n788_), .C2(new_n792_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(G1339gat));
  NOR4_X1   g596(.A1(new_n297_), .A2(new_n468_), .A3(new_n465_), .A4(new_n469_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT59), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT56), .ZN(new_n801_));
  INV_X1    g600(.A(new_n561_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n802_), .A2(new_n582_), .A3(new_n578_), .A4(new_n584_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n503_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n585_), .A2(KEYINPUT55), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n585_), .A2(KEYINPUT55), .ZN(new_n806_));
  OAI211_X1 g605(.A(KEYINPUT114), .B(new_n804_), .C1(new_n805_), .C2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n592_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n576_), .A2(new_n535_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n581_), .B1(new_n809_), .B2(new_n527_), .ZN(new_n810_));
  AOI22_X1  g609(.A1(new_n564_), .A2(new_n558_), .B1(new_n810_), .B2(KEYINPUT68), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(new_n582_), .A4(new_n579_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n585_), .A2(KEYINPUT55), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT114), .B1(new_n815_), .B2(new_n804_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n801_), .B1(new_n808_), .B2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n804_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT114), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n820_), .A2(KEYINPUT56), .A3(new_n592_), .A4(new_n807_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n817_), .A2(new_n821_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n231_), .A2(new_n238_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n230_), .A2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n243_), .B1(new_n237_), .B2(new_n232_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT115), .B1(new_n249_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n829_));
  AOI211_X1 g628(.A(new_n829_), .B(new_n826_), .C1(new_n247_), .C2(new_n248_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n594_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n822_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT58), .ZN(new_n834_));
  AOI22_X1  g633(.A1(new_n833_), .A2(new_n834_), .B1(new_n649_), .B2(new_n653_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n822_), .A2(KEYINPUT58), .A3(new_n832_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n836_), .A2(KEYINPUT116), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT116), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n831_), .B1(new_n817_), .B2(new_n821_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n838_), .B1(new_n839_), .B2(KEYINPUT58), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n835_), .B1(new_n837_), .B2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n250_), .A2(new_n594_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n817_), .B2(new_n821_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n595_), .A2(new_n598_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n828_), .A2(new_n830_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n652_), .B1(new_n843_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n841_), .A2(KEYINPUT119), .A3(new_n849_), .ZN(new_n850_));
  OAI211_X1 g649(.A(KEYINPUT57), .B(new_n652_), .C1(new_n843_), .C2(new_n846_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(KEYINPUT119), .B1(new_n841_), .B2(new_n849_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n615_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n705_), .A2(new_n615_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT54), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n855_), .A2(new_n856_), .A3(new_n251_), .A4(new_n601_), .ZN(new_n857_));
  OAI21_X1  g656(.A(KEYINPUT54), .B1(new_n654_), .B2(new_n250_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n800_), .B1(new_n854_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n849_), .A2(new_n851_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n864_));
  AND4_X1   g663(.A1(new_n650_), .A2(new_n651_), .A3(new_n645_), .A4(new_n648_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n648_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n866_));
  OAI22_X1  g665(.A1(new_n839_), .A2(KEYINPUT58), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n836_), .A2(KEYINPUT116), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n839_), .A2(new_n838_), .A3(KEYINPUT58), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n867_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n863_), .B1(new_n864_), .B2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n841_), .A2(KEYINPUT117), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n616_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n859_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n862_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n849_), .A2(new_n851_), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n835_), .B(new_n864_), .C1(new_n837_), .C2(new_n840_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n870_), .A2(new_n864_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n615_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n880_), .A2(KEYINPUT118), .A3(new_n859_), .ZN(new_n881_));
  AND3_X1   g680(.A1(new_n875_), .A2(new_n881_), .A3(new_n798_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n861_), .B1(new_n882_), .B2(new_n799_), .ZN(new_n883_));
  OAI21_X1  g682(.A(G113gat), .B1(new_n883_), .B2(new_n251_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n875_), .A2(new_n881_), .A3(new_n798_), .ZN(new_n885_));
  OR3_X1    g684(.A1(new_n885_), .A2(G113gat), .A3(new_n251_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n886_), .ZN(G1340gat));
  OAI21_X1  g686(.A(G120gat), .B1(new_n883_), .B2(new_n601_), .ZN(new_n888_));
  INV_X1    g687(.A(G120gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n889_), .B1(new_n601_), .B2(KEYINPUT60), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n882_), .B(new_n890_), .C1(KEYINPUT60), .C2(new_n889_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n888_), .A2(new_n891_), .ZN(G1341gat));
  INV_X1    g691(.A(G127gat), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n615_), .A2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  AOI211_X1 g694(.A(new_n860_), .B(new_n895_), .C1(new_n885_), .C2(KEYINPUT59), .ZN(new_n896_));
  AOI21_X1  g695(.A(G127gat), .B1(new_n882_), .B2(new_n616_), .ZN(new_n897_));
  OAI21_X1  g696(.A(KEYINPUT120), .B1(new_n896_), .B2(new_n897_), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n861_), .B(new_n894_), .C1(new_n882_), .C2(new_n799_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n893_), .B1(new_n885_), .B2(new_n615_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n899_), .A2(new_n900_), .A3(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n898_), .A2(new_n902_), .ZN(G1342gat));
  OAI21_X1  g702(.A(G134gat), .B1(new_n883_), .B2(new_n781_), .ZN(new_n904_));
  OR3_X1    g703(.A1(new_n885_), .A2(G134gat), .A3(new_n652_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1343gat));
  NAND3_X1  g705(.A1(new_n872_), .A2(new_n877_), .A3(new_n876_), .ZN(new_n907_));
  AOI211_X1 g706(.A(new_n862_), .B(new_n874_), .C1(new_n907_), .C2(new_n615_), .ZN(new_n908_));
  AOI21_X1  g707(.A(KEYINPUT118), .B1(new_n880_), .B2(new_n859_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n692_), .A2(new_n465_), .A3(new_n469_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n910_), .A2(new_n468_), .A3(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(KEYINPUT121), .B(G141gat), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n913_), .A2(new_n250_), .A3(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n914_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n916_), .B1(new_n912_), .B2(new_n251_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n915_), .A2(new_n917_), .ZN(G1344gat));
  NAND3_X1  g717(.A1(new_n913_), .A2(new_n312_), .A3(new_n663_), .ZN(new_n919_));
  OAI21_X1  g718(.A(G148gat), .B1(new_n912_), .B2(new_n601_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(G1345gat));
  XNOR2_X1  g720(.A(KEYINPUT61), .B(G155gat), .ZN(new_n922_));
  OR3_X1    g721(.A1(new_n912_), .A2(new_n615_), .A3(new_n922_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n922_), .B1(new_n912_), .B2(new_n615_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1346gat));
  NAND2_X1  g724(.A1(new_n705_), .A2(G162gat), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(KEYINPUT122), .ZN(new_n927_));
  NAND4_X1  g726(.A1(new_n910_), .A2(new_n468_), .A3(new_n644_), .A4(new_n911_), .ZN(new_n928_));
  AOI22_X1  g727(.A1(new_n913_), .A2(new_n927_), .B1(new_n928_), .B2(new_n301_), .ZN(G1347gat));
  NAND2_X1  g728(.A1(new_n854_), .A2(new_n859_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n500_), .A2(new_n465_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n932_), .A2(new_n468_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n933_), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n931_), .A2(new_n251_), .A3(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n936_));
  INV_X1    g735(.A(G169gat), .ZN(new_n937_));
  OR3_X1    g736(.A1(new_n935_), .A2(new_n936_), .A3(new_n937_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n936_), .B1(new_n935_), .B2(new_n937_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n935_), .A2(new_n271_), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n938_), .A2(new_n939_), .A3(new_n940_), .ZN(G1348gat));
  NOR2_X1   g740(.A1(new_n931_), .A2(new_n934_), .ZN(new_n942_));
  AOI21_X1  g741(.A(G176gat), .B1(new_n942_), .B2(new_n663_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT123), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n910_), .A2(new_n944_), .A3(new_n404_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n875_), .A2(new_n881_), .ZN(new_n946_));
  OAI21_X1  g745(.A(KEYINPUT123), .B1(new_n946_), .B2(new_n468_), .ZN(new_n947_));
  INV_X1    g746(.A(new_n932_), .ZN(new_n948_));
  AND3_X1   g747(.A1(new_n945_), .A2(new_n947_), .A3(new_n948_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n601_), .A2(new_n268_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n943_), .B1(new_n949_), .B2(new_n950_), .ZN(G1349gat));
  NAND4_X1  g750(.A1(new_n945_), .A2(new_n947_), .A3(new_n616_), .A4(new_n948_), .ZN(new_n952_));
  INV_X1    g751(.A(new_n264_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n615_), .A2(new_n412_), .ZN(new_n954_));
  AOI22_X1  g753(.A1(new_n952_), .A2(new_n953_), .B1(new_n942_), .B2(new_n954_), .ZN(G1350gat));
  NAND3_X1  g754(.A1(new_n942_), .A2(new_n413_), .A3(new_n644_), .ZN(new_n956_));
  NOR3_X1   g755(.A1(new_n931_), .A2(new_n781_), .A3(new_n934_), .ZN(new_n957_));
  INV_X1    g756(.A(G190gat), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n956_), .B1(new_n957_), .B2(new_n958_), .ZN(G1351gat));
  NOR3_X1   g758(.A1(new_n692_), .A2(new_n466_), .A3(new_n492_), .ZN(new_n960_));
  NAND4_X1  g759(.A1(new_n910_), .A2(new_n250_), .A3(new_n468_), .A4(new_n960_), .ZN(new_n961_));
  OAI21_X1  g760(.A(KEYINPUT124), .B1(new_n961_), .B2(new_n338_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n961_), .A2(new_n338_), .ZN(new_n963_));
  AND4_X1   g762(.A1(new_n468_), .A2(new_n875_), .A3(new_n881_), .A4(new_n960_), .ZN(new_n964_));
  INV_X1    g763(.A(KEYINPUT124), .ZN(new_n965_));
  NAND4_X1  g764(.A1(new_n964_), .A2(new_n965_), .A3(G197gat), .A4(new_n250_), .ZN(new_n966_));
  AND3_X1   g765(.A1(new_n962_), .A2(new_n963_), .A3(new_n966_), .ZN(G1352gat));
  NAND2_X1  g766(.A1(new_n964_), .A2(new_n663_), .ZN(new_n968_));
  XNOR2_X1  g767(.A(KEYINPUT125), .B(G204gat), .ZN(new_n969_));
  INV_X1    g768(.A(new_n969_), .ZN(new_n970_));
  XNOR2_X1  g769(.A(new_n968_), .B(new_n970_), .ZN(G1353gat));
  AOI21_X1  g770(.A(new_n615_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n964_), .A2(new_n972_), .ZN(new_n973_));
  NOR2_X1   g772(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n974_));
  XNOR2_X1  g773(.A(new_n974_), .B(KEYINPUT126), .ZN(new_n975_));
  XNOR2_X1  g774(.A(new_n973_), .B(new_n975_), .ZN(G1354gat));
  INV_X1    g775(.A(new_n964_), .ZN(new_n977_));
  OAI21_X1  g776(.A(G218gat), .B1(new_n977_), .B2(new_n781_), .ZN(new_n978_));
  OR2_X1    g777(.A1(new_n652_), .A2(G218gat), .ZN(new_n979_));
  OAI21_X1  g778(.A(new_n978_), .B1(new_n977_), .B2(new_n979_), .ZN(G1355gat));
endmodule


