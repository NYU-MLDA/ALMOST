//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 0 1 1 0 1 0 1 1 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 0 0 0 0 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n911_,
    new_n913_, new_n914_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_;
  NOR2_X1   g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT84), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT1), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n208_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n209_), .B(KEYINPUT3), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n211_), .B(KEYINPUT2), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n212_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT85), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G127gat), .B(G134gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G113gat), .B(G120gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(KEYINPUT82), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n212_), .A2(new_n216_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT85), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n219_), .A2(new_n223_), .A3(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n226_), .A2(KEYINPUT4), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n217_), .A2(new_n222_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(KEYINPUT4), .A3(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n227_), .B1(KEYINPUT95), .B2(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n226_), .A2(new_n228_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT95), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(new_n232_), .A3(KEYINPUT4), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n230_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G225gat), .A2(G233gat), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(G1gat), .B(G29gat), .Z(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G57gat), .B(G85gat), .ZN(new_n241_));
  XOR2_X1   g040(.A(new_n240_), .B(new_n241_), .Z(new_n242_));
  NOR2_X1   g041(.A1(new_n231_), .A2(new_n236_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n237_), .A2(new_n242_), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n242_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n235_), .B1(new_n230_), .B2(new_n233_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n246_), .B1(new_n247_), .B2(new_n243_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n245_), .A2(KEYINPUT99), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT99), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n237_), .A2(new_n250_), .A3(new_n242_), .A4(new_n244_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT22), .B(G169gat), .ZN(new_n253_));
  INV_X1    g052(.A(G176gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(new_n255_), .B(KEYINPUT81), .Z(new_n256_));
  NOR2_X1   g055(.A1(G183gat), .A2(G190gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT23), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G183gat), .A2(G190gat), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n257_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n261_));
  AOI22_X1  g060(.A1(new_n260_), .A2(new_n261_), .B1(G169gat), .B2(G176gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n256_), .A2(new_n262_), .ZN(new_n263_));
  OR2_X1    g062(.A1(G169gat), .A2(G176gat), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n264_), .A2(KEYINPUT24), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n259_), .A2(KEYINPUT23), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n258_), .A2(G183gat), .A3(G190gat), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n265_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT25), .B(G183gat), .ZN(new_n269_));
  INV_X1    g068(.A(G190gat), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT26), .B1(new_n270_), .B2(KEYINPUT80), .ZN(new_n271_));
  OR2_X1    g070(.A1(new_n270_), .A2(KEYINPUT26), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n269_), .B(new_n271_), .C1(new_n272_), .C2(KEYINPUT80), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G169gat), .A2(G176gat), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n264_), .A2(KEYINPUT24), .A3(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n268_), .A2(new_n273_), .A3(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n263_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G227gat), .A2(G233gat), .ZN(new_n278_));
  INV_X1    g077(.A(G15gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT30), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n277_), .B(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(G71gat), .B(G99gat), .Z(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(G43gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n282_), .B(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n223_), .B(KEYINPUT31), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT83), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n285_), .A2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n286_), .A2(KEYINPUT83), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n285_), .B1(new_n290_), .B2(new_n288_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n252_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT91), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G211gat), .B(G218gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT86), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G197gat), .B(G204gat), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT21), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT87), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n295_), .B(KEYINPUT86), .Z(new_n302_));
  XNOR2_X1  g101(.A(new_n297_), .B(KEYINPUT21), .ZN(new_n303_));
  AOI22_X1  g102(.A1(new_n300_), .A2(new_n301_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  AND3_X1   g103(.A1(new_n302_), .A2(new_n303_), .A3(new_n301_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G228gat), .A2(G233gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT29), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n219_), .A2(new_n225_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n309_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n217_), .A2(new_n310_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n308_), .B1(new_n306_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT90), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G78gat), .B(G106gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n317_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n312_), .B(new_n314_), .C1(KEYINPUT90), .C2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G22gat), .B(G50gat), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT28), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n311_), .A2(new_n324_), .A3(new_n310_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n324_), .B1(new_n311_), .B2(new_n310_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n323_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n311_), .A2(new_n310_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT28), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n330_), .A2(new_n325_), .A3(new_n322_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n294_), .B1(new_n321_), .B2(new_n332_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n328_), .A2(new_n331_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n334_), .A2(KEYINPUT91), .A3(new_n318_), .A4(new_n320_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n317_), .A2(KEYINPUT88), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n315_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n337_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n317_), .A2(KEYINPUT88), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n312_), .A2(new_n339_), .A3(new_n314_), .A4(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT89), .B1(new_n334_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT89), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n332_), .A2(new_n344_), .A3(new_n338_), .A4(new_n341_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n336_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT27), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n277_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT26), .B(G190gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n269_), .A2(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT92), .B1(new_n351_), .B2(new_n275_), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n266_), .A2(new_n267_), .ZN(new_n353_));
  NOR3_X1   g152(.A1(new_n352_), .A2(new_n265_), .A3(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n351_), .A2(KEYINPUT92), .A3(new_n275_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n253_), .B(KEYINPUT93), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n254_), .ZN(new_n357_));
  AOI22_X1  g156(.A1(new_n354_), .A2(new_n355_), .B1(new_n357_), .B2(new_n262_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n306_), .A2(new_n358_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n349_), .A2(new_n359_), .A3(KEYINPUT20), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT19), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n360_), .A2(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n306_), .A2(new_n358_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT20), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n306_), .A2(new_n263_), .A3(new_n276_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n367_), .A2(new_n363_), .A3(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n364_), .A2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G8gat), .B(G36gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT18), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G64gat), .B(G92gat), .ZN(new_n373_));
  XOR2_X1   g172(.A(new_n372_), .B(new_n373_), .Z(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n348_), .B1(new_n370_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT94), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n360_), .A2(new_n377_), .A3(new_n363_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n363_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n349_), .A2(new_n359_), .A3(KEYINPUT20), .A4(new_n363_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT94), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n378_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(new_n374_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n376_), .A2(new_n383_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n378_), .B(new_n375_), .C1(new_n379_), .C2(new_n381_), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n384_), .B1(new_n386_), .B2(KEYINPUT27), .ZN(new_n387_));
  NOR3_X1   g186(.A1(new_n293_), .A2(new_n347_), .A3(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n374_), .A2(KEYINPUT32), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n389_), .B1(new_n364_), .B2(new_n369_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n390_), .B1(new_n389_), .B2(new_n382_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n249_), .A2(new_n251_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT33), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n248_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT98), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n395_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n230_), .A2(new_n233_), .A3(KEYINPUT98), .A4(new_n235_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n226_), .A2(new_n228_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n242_), .B1(new_n398_), .B2(new_n235_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT97), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n396_), .A2(new_n397_), .A3(new_n400_), .ZN(new_n401_));
  OAI211_X1 g200(.A(KEYINPUT33), .B(new_n246_), .C1(new_n247_), .C2(new_n243_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n386_), .A2(new_n394_), .A3(new_n401_), .A4(new_n402_), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n392_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n252_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n383_), .A2(new_n385_), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n406_), .A2(new_n348_), .B1(new_n376_), .B2(new_n383_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n347_), .A2(new_n407_), .ZN(new_n408_));
  OAI22_X1  g207(.A1(new_n404_), .A2(new_n347_), .B1(new_n405_), .B2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n292_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n388_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G29gat), .B(G36gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G43gat), .B(G50gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT15), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G1gat), .B(G8gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT75), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G15gat), .B(G22gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G1gat), .A2(G8gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT14), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n418_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n417_), .A2(new_n421_), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n416_), .A2(KEYINPUT75), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n416_), .A2(KEYINPUT75), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n423_), .A2(new_n420_), .A3(new_n418_), .A4(new_n424_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n422_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n415_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n422_), .A2(new_n425_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n414_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G229gat), .A2(G233gat), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n427_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT78), .ZN(new_n432_));
  INV_X1    g231(.A(new_n414_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n422_), .A2(new_n433_), .A3(new_n425_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n429_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n430_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n432_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  AOI211_X1 g236(.A(KEYINPUT78), .B(new_n430_), .C1(new_n429_), .C2(new_n434_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n431_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G113gat), .B(G141gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G169gat), .B(G197gat), .ZN(new_n441_));
  XOR2_X1   g240(.A(new_n440_), .B(new_n441_), .Z(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n439_), .A2(KEYINPUT79), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(KEYINPUT79), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n445_), .B(new_n431_), .C1(new_n437_), .C2(new_n438_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT13), .ZN(new_n449_));
  INV_X1    g248(.A(G230gat), .ZN(new_n450_));
  INV_X1    g249(.A(G233gat), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G85gat), .B(G92gat), .ZN(new_n453_));
  INV_X1    g252(.A(G92gat), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n453_), .B1(KEYINPUT9), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(G85gat), .ZN(new_n456_));
  OR2_X1    g255(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n456_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  XOR2_X1   g258(.A(KEYINPUT64), .B(KEYINPUT9), .Z(new_n460_));
  OAI21_X1  g259(.A(new_n455_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G99gat), .A2(G106gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT6), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT6), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n464_), .A2(G99gat), .A3(G106gat), .ZN(new_n465_));
  AND3_X1   g264(.A1(new_n463_), .A2(new_n465_), .A3(KEYINPUT66), .ZN(new_n466_));
  AOI21_X1  g265(.A(KEYINPUT66), .B1(new_n463_), .B2(new_n465_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  XOR2_X1   g267(.A(KEYINPUT10), .B(G99gat), .Z(new_n469_));
  INV_X1    g268(.A(G106gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n461_), .A2(new_n468_), .A3(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT8), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n463_), .A2(new_n465_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT68), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT68), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n463_), .A2(new_n465_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(G99gat), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT67), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n478_), .B(new_n470_), .C1(new_n479_), .C2(KEYINPUT7), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT7), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n481_), .B(KEYINPUT67), .C1(G99gat), .C2(G106gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n475_), .A2(new_n477_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n453_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n473_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n453_), .A2(KEYINPUT8), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n488_), .B1(new_n468_), .B2(new_n483_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n472_), .B1(new_n486_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT69), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  OAI211_X1 g291(.A(KEYINPUT69), .B(new_n472_), .C1(new_n486_), .C2(new_n489_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G57gat), .B(G64gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT11), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT70), .ZN(new_n496_));
  OR2_X1    g295(.A1(new_n494_), .A2(KEYINPUT11), .ZN(new_n497_));
  XOR2_X1   g296(.A(G71gat), .B(G78gat), .Z(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n496_), .B(new_n499_), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n492_), .A2(new_n493_), .A3(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n500_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n452_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(G120gat), .B(G148gat), .Z(new_n504_));
  XNOR2_X1  g303(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G176gat), .B(G204gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n497_), .A2(new_n498_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n496_), .B(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n511_), .A2(KEYINPUT12), .A3(new_n490_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n512_), .B1(new_n502_), .B2(KEYINPUT12), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n492_), .A2(new_n493_), .A3(new_n500_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n514_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n503_), .B(new_n509_), .C1(new_n513_), .C2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n493_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT66), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n474_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n463_), .A2(new_n465_), .A3(KEYINPUT66), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(new_n521_), .A3(new_n483_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(new_n487_), .ZN(new_n523_));
  AOI22_X1  g322(.A1(new_n474_), .A2(KEYINPUT68), .B1(new_n480_), .B2(new_n482_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n453_), .B1(new_n524_), .B2(new_n477_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n523_), .B1(new_n525_), .B2(new_n473_), .ZN(new_n526_));
  AOI21_X1  g325(.A(KEYINPUT69), .B1(new_n526_), .B2(new_n472_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n518_), .A2(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n452_), .B1(new_n528_), .B2(new_n500_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n511_), .B1(new_n518_), .B2(new_n527_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT12), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n529_), .A2(new_n532_), .A3(new_n512_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n509_), .B1(new_n533_), .B2(new_n503_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n449_), .B1(new_n517_), .B2(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n503_), .B1(new_n513_), .B2(new_n515_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(new_n508_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n537_), .A2(KEYINPUT13), .A3(new_n516_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n535_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT72), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G190gat), .B(G218gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT74), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G134gat), .B(G162gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT36), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n544_), .A2(new_n545_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G232gat), .A2(G233gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT34), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT35), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n490_), .A2(new_n415_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT73), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n492_), .A2(new_n414_), .A3(new_n493_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n550_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n549_), .B(KEYINPUT35), .Z(new_n555_));
  NAND3_X1  g354(.A1(new_n553_), .A2(new_n551_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n546_), .B(new_n547_), .C1(new_n554_), .C2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT73), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n551_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n553_), .ZN(new_n561_));
  OAI211_X1 g360(.A(KEYINPUT35), .B(new_n549_), .C1(new_n560_), .C2(new_n561_), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n562_), .A2(new_n545_), .A3(new_n544_), .A4(new_n556_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n558_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT37), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n558_), .A2(new_n563_), .A3(KEYINPUT37), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(G231gat), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n570_), .A2(new_n451_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n426_), .A2(new_n571_), .ZN(new_n572_));
  NOR3_X1   g371(.A1(new_n428_), .A2(new_n570_), .A3(new_n451_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n511_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n426_), .A2(new_n571_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n428_), .B1(new_n570_), .B2(new_n451_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n500_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G127gat), .B(G155gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G183gat), .B(G211gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT17), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n574_), .A2(new_n577_), .A3(new_n583_), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n582_), .A2(KEYINPUT17), .ZN(new_n585_));
  AOI22_X1  g384(.A1(new_n574_), .A2(new_n577_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(KEYINPUT77), .B1(new_n584_), .B2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n574_), .A2(new_n577_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n585_), .A2(new_n583_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT77), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n574_), .A2(new_n577_), .A3(new_n583_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n590_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n587_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n569_), .A2(new_n595_), .ZN(new_n596_));
  OR4_X1    g395(.A1(new_n411_), .A2(new_n448_), .A3(new_n540_), .A4(new_n596_), .ZN(new_n597_));
  NOR3_X1   g396(.A1(new_n597_), .A2(G1gat), .A3(new_n252_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT38), .Z(new_n599_));
  AND3_X1   g398(.A1(new_n252_), .A2(new_n347_), .A3(new_n407_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n347_), .B1(new_n392_), .B2(new_n403_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n410_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n387_), .A2(new_n347_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(new_n252_), .A3(new_n292_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(KEYINPUT100), .B1(new_n605_), .B2(new_n564_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT100), .ZN(new_n607_));
  INV_X1    g406(.A(new_n564_), .ZN(new_n608_));
  AOI211_X1 g407(.A(new_n607_), .B(new_n608_), .C1(new_n602_), .C2(new_n604_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n606_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n539_), .A2(new_n448_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n613_), .A2(new_n594_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n611_), .A2(new_n405_), .A3(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(G1gat), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n599_), .A2(new_n616_), .ZN(G1324gat));
  XNOR2_X1  g416(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n387_), .B(new_n614_), .C1(new_n606_), .C2(new_n609_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(G8gat), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(KEYINPUT39), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT39), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n619_), .A2(new_n622_), .A3(G8gat), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  OR3_X1    g423(.A1(new_n597_), .A2(G8gat), .A3(new_n407_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n618_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n619_), .A2(new_n622_), .A3(G8gat), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n622_), .B1(new_n619_), .B2(G8gat), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n625_), .B(new_n618_), .C1(new_n627_), .C2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n626_), .A2(new_n630_), .ZN(G1325gat));
  INV_X1    g430(.A(new_n597_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(new_n279_), .A3(new_n292_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n611_), .A2(new_n292_), .A3(new_n614_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n634_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n635_));
  AOI21_X1  g434(.A(KEYINPUT41), .B1(new_n634_), .B2(G15gat), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n633_), .B1(new_n635_), .B2(new_n636_), .ZN(G1326gat));
  INV_X1    g436(.A(new_n347_), .ZN(new_n638_));
  OR3_X1    g437(.A1(new_n597_), .A2(G22gat), .A3(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n611_), .A2(new_n347_), .A3(new_n614_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(G22gat), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n641_), .A2(KEYINPUT42), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n641_), .A2(KEYINPUT42), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n639_), .B1(new_n642_), .B2(new_n643_), .ZN(G1327gat));
  INV_X1    g443(.A(new_n539_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n564_), .A2(new_n595_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  AOI211_X1 g446(.A(new_n448_), .B(new_n647_), .C1(new_n602_), .C2(new_n604_), .ZN(new_n648_));
  AOI21_X1  g447(.A(G29gat), .B1(new_n648_), .B2(new_n405_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n613_), .A2(new_n595_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(new_n605_), .B2(new_n568_), .ZN(new_n652_));
  AOI211_X1 g451(.A(KEYINPUT43), .B(new_n569_), .C1(new_n602_), .C2(new_n604_), .ZN(new_n653_));
  OAI211_X1 g452(.A(KEYINPUT44), .B(new_n650_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n650_), .ZN(new_n655_));
  OAI21_X1  g454(.A(KEYINPUT43), .B1(new_n411_), .B2(new_n569_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n605_), .A2(new_n651_), .A3(new_n568_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n655_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT102), .B(KEYINPUT44), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n654_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n405_), .A2(G29gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n649_), .B1(new_n661_), .B2(new_n662_), .ZN(G1328gat));
  OAI211_X1 g462(.A(new_n387_), .B(new_n654_), .C1(new_n658_), .C2(new_n659_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(G36gat), .ZN(new_n665_));
  NOR2_X1   g464(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT103), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n407_), .A2(G36gat), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n648_), .A2(new_n667_), .A3(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n647_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n605_), .A2(new_n447_), .A3(new_n670_), .A4(new_n668_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT103), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n669_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT45), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT45), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n669_), .A2(new_n672_), .A3(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n666_), .B1(new_n674_), .B2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n665_), .A2(new_n677_), .ZN(new_n678_));
  OAI21_X1  g477(.A(KEYINPUT105), .B1(KEYINPUT104), .B2(KEYINPUT46), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT106), .Z(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n678_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n665_), .A2(new_n677_), .A3(new_n680_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1329gat));
  NAND2_X1  g483(.A1(new_n292_), .A2(G43gat), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n648_), .A2(new_n292_), .ZN(new_n686_));
  OAI22_X1  g485(.A1(new_n660_), .A2(new_n685_), .B1(G43gat), .B2(new_n686_), .ZN(new_n687_));
  XOR2_X1   g486(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(G1330gat));
  AOI21_X1  g488(.A(G50gat), .B1(new_n648_), .B2(new_n347_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n347_), .A2(G50gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n661_), .B2(new_n691_), .ZN(G1331gat));
  NOR2_X1   g491(.A1(new_n594_), .A2(new_n447_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n540_), .A2(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n610_), .A2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(new_n405_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(G57gat), .ZN(new_n697_));
  NOR4_X1   g496(.A1(new_n411_), .A2(new_n447_), .A3(new_n645_), .A4(new_n596_), .ZN(new_n698_));
  INV_X1    g497(.A(G57gat), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n698_), .A2(new_n699_), .A3(new_n405_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n697_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(KEYINPUT108), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n697_), .A2(new_n703_), .A3(new_n700_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(G1332gat));
  INV_X1    g504(.A(G64gat), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n698_), .A2(new_n706_), .A3(new_n387_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT48), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n695_), .A2(new_n387_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n709_), .B2(G64gat), .ZN(new_n710_));
  AOI211_X1 g509(.A(KEYINPUT48), .B(new_n706_), .C1(new_n695_), .C2(new_n387_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n710_), .B2(new_n711_), .ZN(G1333gat));
  INV_X1    g511(.A(G71gat), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n698_), .A2(new_n713_), .A3(new_n292_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT49), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n695_), .A2(new_n292_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n716_), .B2(G71gat), .ZN(new_n717_));
  AOI211_X1 g516(.A(KEYINPUT49), .B(new_n713_), .C1(new_n695_), .C2(new_n292_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n714_), .B1(new_n717_), .B2(new_n718_), .ZN(G1334gat));
  INV_X1    g518(.A(G78gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n698_), .A2(new_n720_), .A3(new_n347_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT50), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n695_), .A2(new_n347_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n723_), .B2(G78gat), .ZN(new_n724_));
  AOI211_X1 g523(.A(KEYINPUT50), .B(new_n720_), .C1(new_n695_), .C2(new_n347_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n721_), .B1(new_n724_), .B2(new_n725_), .ZN(G1335gat));
  NAND2_X1  g525(.A1(new_n656_), .A2(new_n657_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n645_), .A2(new_n595_), .A3(new_n447_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G85gat), .B1(new_n729_), .B2(new_n252_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n411_), .A2(new_n447_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n540_), .A2(new_n646_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n733_), .A2(new_n456_), .A3(new_n405_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n730_), .A2(new_n734_), .ZN(G1336gat));
  AOI21_X1  g534(.A(G92gat), .B1(new_n733_), .B2(new_n387_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n729_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n407_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n736_), .B1(new_n737_), .B2(new_n738_), .ZN(G1337gat));
  OAI21_X1  g538(.A(G99gat), .B1(new_n729_), .B2(new_n410_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n733_), .A2(new_n292_), .A3(new_n469_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(KEYINPUT109), .B(KEYINPUT51), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n742_), .B(new_n743_), .ZN(G1338gat));
  OAI211_X1 g543(.A(new_n347_), .B(new_n728_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(G106gat), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT52), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n745_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n638_), .A2(G106gat), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n731_), .A2(new_n732_), .A3(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT110), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n731_), .A2(new_n753_), .A3(new_n732_), .A4(new_n750_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n748_), .A2(new_n749_), .A3(new_n755_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g556(.A1(new_n603_), .A2(new_n405_), .A3(new_n292_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT119), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT119), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n603_), .A2(new_n760_), .A3(new_n405_), .A4(new_n292_), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n759_), .A2(KEYINPUT121), .A3(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(KEYINPUT121), .B1(new_n759_), .B2(new_n761_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n764_));
  NOR3_X1   g563(.A1(new_n762_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n535_), .A2(new_n538_), .A3(new_n693_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT111), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT111), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n535_), .A2(new_n693_), .A3(new_n538_), .A4(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n569_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT113), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT113), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n770_), .A2(new_n774_), .A3(new_n569_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n772_), .A2(new_n773_), .A3(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n774_), .B1(new_n770_), .B2(new_n569_), .ZN(new_n777_));
  AOI211_X1 g576(.A(KEYINPUT113), .B(new_n568_), .C1(new_n767_), .C2(new_n769_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT112), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n776_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT54), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n776_), .A2(new_n779_), .A3(KEYINPUT54), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n427_), .A2(new_n429_), .A3(new_n436_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n436_), .B1(new_n429_), .B2(new_n434_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n443_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n439_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n787_), .B1(new_n788_), .B2(new_n443_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT116), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT116), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n791_), .B(new_n787_), .C1(new_n788_), .C2(new_n443_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n537_), .A2(new_n516_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n448_), .A2(new_n517_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n511_), .A2(KEYINPUT12), .A3(new_n490_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n798_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n799_), .A2(KEYINPUT55), .A3(new_n529_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n452_), .B1(new_n513_), .B2(new_n501_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT55), .B1(new_n799_), .B2(new_n529_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n800_), .B(new_n801_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n533_), .A2(new_n803_), .A3(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n508_), .B1(new_n804_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT56), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n805_), .B1(new_n513_), .B2(new_n515_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT114), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n812_), .A2(new_n806_), .A3(new_n800_), .A4(new_n801_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n813_), .A2(KEYINPUT56), .A3(new_n508_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n797_), .B1(new_n810_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n795_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n813_), .A2(KEYINPUT56), .A3(new_n508_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT56), .B1(new_n813_), .B2(new_n508_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n796_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n820_), .A2(KEYINPUT115), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n564_), .B1(new_n817_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT57), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT117), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n810_), .A2(new_n824_), .A3(new_n814_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n790_), .A2(new_n516_), .A3(new_n792_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n826_), .B1(new_n819_), .B2(KEYINPUT117), .ZN(new_n827_));
  NOR2_X1   g626(.A1(KEYINPUT118), .A2(KEYINPUT58), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n825_), .A2(new_n827_), .A3(new_n829_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n830_), .A2(new_n568_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n825_), .A2(new_n827_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n828_), .ZN(new_n833_));
  AOI22_X1  g632(.A1(new_n822_), .A2(new_n823_), .B1(new_n831_), .B2(new_n833_), .ZN(new_n834_));
  AOI22_X1  g633(.A1(new_n820_), .A2(KEYINPUT115), .B1(new_n794_), .B2(new_n793_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n815_), .A2(new_n816_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n608_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT57), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n595_), .B1(new_n834_), .B2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n765_), .B1(new_n784_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n759_), .A2(new_n761_), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n776_), .A2(new_n779_), .A3(KEYINPUT54), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT54), .B1(new_n776_), .B2(new_n779_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n833_), .A2(new_n568_), .A3(new_n830_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(new_n837_), .B2(KEYINPUT57), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n822_), .A2(new_n823_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n594_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n841_), .B1(new_n844_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n840_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(G113gat), .B1(new_n851_), .B2(new_n448_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n844_), .A2(new_n848_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n841_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  OR2_X1    g654(.A1(new_n448_), .A2(G113gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n852_), .B1(new_n855_), .B2(new_n856_), .ZN(G1340gat));
  INV_X1    g656(.A(new_n540_), .ZN(new_n858_));
  OAI21_X1  g657(.A(G120gat), .B1(new_n851_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(G120gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n645_), .B2(KEYINPUT60), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n861_), .B1(KEYINPUT60), .B2(new_n860_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n859_), .B1(new_n855_), .B2(new_n862_), .ZN(G1341gat));
  INV_X1    g662(.A(G127gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n864_), .B1(new_n855_), .B2(new_n594_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  OAI211_X1 g666(.A(KEYINPUT122), .B(new_n864_), .C1(new_n855_), .C2(new_n594_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n851_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n594_), .A2(new_n864_), .ZN(new_n870_));
  AOI22_X1  g669(.A1(new_n867_), .A2(new_n868_), .B1(new_n869_), .B2(new_n870_), .ZN(G1342gat));
  INV_X1    g670(.A(G134gat), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n569_), .A2(new_n872_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n840_), .B(new_n873_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n608_), .B(new_n854_), .C1(new_n784_), .C2(new_n839_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n872_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT123), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n874_), .A2(KEYINPUT123), .A3(new_n876_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1343gat));
  NOR2_X1   g680(.A1(new_n784_), .A2(new_n839_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n408_), .A2(new_n252_), .A3(new_n292_), .ZN(new_n883_));
  XOR2_X1   g682(.A(new_n883_), .B(KEYINPUT124), .Z(new_n884_));
  NOR2_X1   g683(.A1(new_n882_), .A2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n447_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n540_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT125), .B(G148gat), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1345gat));
  NAND2_X1  g689(.A1(new_n885_), .A2(new_n595_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT61), .B(G155gat), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(G1346gat));
  INV_X1    g692(.A(G162gat), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n885_), .A2(new_n894_), .A3(new_n608_), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n882_), .A2(new_n569_), .A3(new_n884_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n894_), .B2(new_n896_), .ZN(G1347gat));
  NOR3_X1   g696(.A1(new_n293_), .A2(new_n347_), .A3(new_n407_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n853_), .A2(new_n447_), .A3(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(G169gat), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT62), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n898_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n882_), .A2(new_n903_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n904_), .A2(new_n356_), .A3(new_n447_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n899_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n902_), .A2(new_n905_), .A3(new_n906_), .ZN(G1348gat));
  NAND3_X1  g706(.A1(new_n904_), .A2(new_n254_), .A3(new_n539_), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n882_), .A2(new_n858_), .A3(new_n903_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n254_), .B2(new_n909_), .ZN(G1349gat));
  NOR3_X1   g709(.A1(new_n882_), .A2(new_n594_), .A3(new_n903_), .ZN(new_n911_));
  MUX2_X1   g710(.A(G183gat), .B(new_n269_), .S(new_n911_), .Z(G1350gat));
  NAND3_X1  g711(.A1(new_n904_), .A2(new_n350_), .A3(new_n608_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n882_), .A2(new_n569_), .A3(new_n903_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n270_), .B2(new_n914_), .ZN(G1351gat));
  NOR4_X1   g714(.A1(new_n405_), .A2(new_n638_), .A3(new_n407_), .A4(new_n292_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n916_), .B1(new_n784_), .B2(new_n839_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT126), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  OAI211_X1 g718(.A(KEYINPUT126), .B(new_n916_), .C1(new_n784_), .C2(new_n839_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  AOI21_X1  g720(.A(G197gat), .B1(new_n921_), .B2(new_n447_), .ZN(new_n922_));
  INV_X1    g721(.A(G197gat), .ZN(new_n923_));
  AOI211_X1 g722(.A(new_n923_), .B(new_n448_), .C1(new_n919_), .C2(new_n920_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n922_), .A2(new_n924_), .ZN(G1352gat));
  AOI21_X1  g724(.A(KEYINPUT126), .B1(new_n853_), .B2(new_n916_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n920_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n540_), .B1(new_n926_), .B2(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(G204gat), .ZN(new_n929_));
  INV_X1    g728(.A(G204gat), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n921_), .A2(new_n930_), .A3(new_n540_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n929_), .A2(new_n931_), .ZN(G1353gat));
  NOR2_X1   g731(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n933_));
  INV_X1    g732(.A(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n595_), .A2(new_n935_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n936_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n934_), .B1(new_n921_), .B2(new_n937_), .ZN(new_n938_));
  AOI211_X1 g737(.A(new_n933_), .B(new_n936_), .C1(new_n919_), .C2(new_n920_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1354gat));
  INV_X1    g739(.A(G218gat), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n921_), .A2(new_n941_), .A3(new_n608_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n569_), .B1(new_n919_), .B2(new_n920_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n942_), .B1(new_n941_), .B2(new_n943_), .ZN(G1355gat));
endmodule


