//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 1 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 0 0 0 1 1 0 0 0 0 0 0 1 0 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n875_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n902_, new_n904_, new_n905_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_;
  INV_X1    g000(.A(KEYINPUT104), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT85), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(KEYINPUT85), .A2(KEYINPUT23), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT86), .ZN(new_n209_));
  INV_X1    g008(.A(new_n206_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(new_n204_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT86), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n205_), .A2(new_n212_), .A3(new_n206_), .A4(new_n207_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n209_), .A2(new_n211_), .A3(new_n213_), .ZN(new_n214_));
  AND2_X1   g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT24), .ZN(new_n217_));
  NOR3_X1   g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n218_), .A2(KEYINPUT84), .ZN(new_n219_));
  NAND2_X1  g018(.A1(KEYINPUT83), .A2(G190gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT26), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(KEYINPUT83), .A2(KEYINPUT26), .A3(G190gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT25), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(G183gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT82), .B(G183gat), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n224_), .B(new_n226_), .C1(new_n227_), .C2(new_n225_), .ZN(new_n228_));
  INV_X1    g027(.A(G169gat), .ZN(new_n229_));
  INV_X1    g028(.A(G176gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n231_), .A2(KEYINPUT24), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT84), .B1(new_n218_), .B2(new_n232_), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n214_), .A2(new_n219_), .A3(new_n228_), .A4(new_n233_), .ZN(new_n234_));
  AND2_X1   g033(.A1(KEYINPUT85), .A2(KEYINPUT23), .ZN(new_n235_));
  NOR2_X1   g034(.A1(KEYINPUT85), .A2(KEYINPUT23), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n210_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n206_), .A2(KEYINPUT23), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G190gat), .ZN(new_n240_));
  INV_X1    g039(.A(G183gat), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n241_), .A2(KEYINPUT82), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(KEYINPUT82), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n240_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n215_), .B1(new_n239_), .B2(new_n244_), .ZN(new_n245_));
  AND2_X1   g044(.A1(KEYINPUT87), .A2(G169gat), .ZN(new_n246_));
  NOR2_X1   g045(.A1(KEYINPUT87), .A2(G169gat), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT22), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT88), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT88), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n250_), .B(KEYINPUT22), .C1(new_n246_), .C2(new_n247_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT22), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n252_), .A2(KEYINPUT89), .A3(G169gat), .ZN(new_n253_));
  AOI21_X1  g052(.A(KEYINPUT89), .B1(new_n252_), .B2(G169gat), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n249_), .A2(new_n230_), .A3(new_n251_), .A4(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n245_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(G204gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(G197gat), .ZN(new_n259_));
  INV_X1    g058(.A(G197gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(G204gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT21), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT21), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n259_), .A2(new_n261_), .A3(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G211gat), .B(G218gat), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n263_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n266_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n268_), .A2(KEYINPUT21), .A3(new_n262_), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n234_), .A2(new_n257_), .A3(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT20), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT96), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n241_), .A2(new_n240_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n214_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n215_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT22), .B(G169gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n230_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n275_), .A2(new_n276_), .A3(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(KEYINPUT97), .B(KEYINPUT24), .Z(new_n280_));
  OR2_X1    g079(.A1(new_n280_), .A2(new_n231_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT25), .B(G183gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT26), .B(G190gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n280_), .A2(new_n276_), .A3(new_n231_), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n281_), .A2(new_n239_), .A3(new_n284_), .A4(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n279_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n270_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT96), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n271_), .A2(new_n290_), .A3(KEYINPUT20), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n273_), .A2(new_n289_), .A3(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G226gat), .A2(G233gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT19), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n279_), .A2(new_n270_), .A3(new_n286_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n234_), .A2(new_n257_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n288_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n294_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n299_), .A2(KEYINPUT20), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n296_), .A2(new_n298_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G8gat), .B(G36gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(G92gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT18), .B(G64gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT32), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n295_), .A2(new_n302_), .A3(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(KEYINPUT102), .B(KEYINPUT20), .Z(new_n310_));
  NAND3_X1  g109(.A1(new_n296_), .A2(new_n298_), .A3(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n294_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT103), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n273_), .A2(new_n299_), .A3(new_n289_), .A4(new_n291_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT103), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n311_), .A2(new_n315_), .A3(new_n294_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n313_), .A2(new_n314_), .A3(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n317_), .A2(KEYINPUT32), .A3(new_n307_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT92), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G141gat), .A2(G148gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT2), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT2), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n322_), .A2(G141gat), .A3(G148gat), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT3), .ZN(new_n325_));
  INV_X1    g124(.A(G141gat), .ZN(new_n326_));
  INV_X1    g125(.A(G148gat), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n325_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n319_), .B1(new_n324_), .B2(new_n330_), .ZN(new_n331_));
  AND2_X1   g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332_));
  NOR2_X1   g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n321_), .A2(new_n323_), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n335_), .A2(KEYINPUT92), .A3(new_n329_), .A4(new_n328_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n331_), .A2(new_n334_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT1), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n334_), .A2(new_n338_), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n332_), .A2(KEYINPUT1), .B1(new_n326_), .B2(new_n327_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(new_n340_), .A3(new_n320_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n337_), .A2(KEYINPUT98), .A3(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G127gat), .B(G134gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G113gat), .B(G120gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n342_), .A2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(KEYINPUT98), .B1(new_n337_), .B2(new_n341_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n337_), .A2(new_n341_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT98), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(new_n351_), .A3(new_n345_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT4), .B1(new_n349_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n337_), .A2(new_n341_), .ZN(new_n357_));
  NOR3_X1   g156(.A1(new_n357_), .A2(KEYINPUT4), .A3(new_n345_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n354_), .A2(new_n356_), .A3(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G57gat), .B(G85gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G1gat), .B(G29gat), .ZN(new_n364_));
  XOR2_X1   g163(.A(new_n363_), .B(new_n364_), .Z(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT100), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n350_), .A2(new_n351_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n368_), .A2(new_n342_), .A3(new_n346_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(new_n352_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n367_), .B1(new_n370_), .B2(new_n355_), .ZN(new_n371_));
  AOI211_X1 g170(.A(KEYINPUT100), .B(new_n356_), .C1(new_n369_), .C2(new_n352_), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n360_), .B(new_n366_), .C1(new_n371_), .C2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n355_), .B1(new_n349_), .B2(new_n353_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT100), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n370_), .A2(new_n367_), .A3(new_n355_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n366_), .B1(new_n378_), .B2(new_n360_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n309_), .B(new_n318_), .C1(new_n374_), .C2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT33), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n373_), .A2(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n307_), .B1(new_n295_), .B2(new_n302_), .ZN(new_n383_));
  AOI211_X1 g182(.A(new_n306_), .B(new_n301_), .C1(new_n292_), .C2(new_n294_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n354_), .A2(KEYINPUT101), .A3(new_n355_), .A4(new_n359_), .ZN(new_n386_));
  AOI211_X1 g185(.A(new_n356_), .B(new_n358_), .C1(new_n370_), .C2(KEYINPUT4), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT101), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n388_), .B1(new_n370_), .B2(new_n356_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n365_), .B(new_n386_), .C1(new_n387_), .C2(new_n389_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n378_), .A2(KEYINPUT33), .A3(new_n360_), .A4(new_n366_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n382_), .A2(new_n385_), .A3(new_n390_), .A4(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n380_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT95), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n396_), .B1(new_n337_), .B2(new_n341_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n397_), .A2(new_n270_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(KEYINPUT93), .A2(G228gat), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(KEYINPUT93), .A2(G228gat), .ZN(new_n401_));
  OAI21_X1  g200(.A(G233gat), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n394_), .B1(new_n398_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n402_), .ZN(new_n404_));
  OAI211_X1 g203(.A(KEYINPUT95), .B(new_n404_), .C1(new_n397_), .C2(new_n270_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  AOI211_X1 g205(.A(new_n404_), .B(new_n270_), .C1(new_n350_), .C2(KEYINPUT29), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G78gat), .B(G106gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  OR3_X1    g210(.A1(new_n350_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT28), .B1(new_n350_), .B2(KEYINPUT29), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G22gat), .B(G50gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n414_), .B(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n410_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n406_), .A2(new_n418_), .A3(new_n408_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n411_), .A2(new_n417_), .A3(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n414_), .B(new_n415_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n418_), .B1(new_n406_), .B2(new_n408_), .ZN(new_n422_));
  AOI211_X1 g221(.A(new_n410_), .B(new_n407_), .C1(new_n403_), .C2(new_n405_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n421_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n420_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n202_), .B1(new_n393_), .B2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n371_), .A2(new_n372_), .ZN(new_n428_));
  AOI211_X1 g227(.A(new_n355_), .B(new_n358_), .C1(new_n370_), .C2(KEYINPUT4), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n365_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  AND4_X1   g229(.A1(new_n430_), .A2(new_n420_), .A3(new_n424_), .A4(new_n373_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT105), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT27), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n433_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n317_), .A2(new_n306_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n295_), .A2(new_n307_), .A3(new_n302_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n435_), .A2(KEYINPUT27), .A3(new_n436_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n431_), .A2(new_n432_), .A3(new_n434_), .A4(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n434_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n430_), .A2(new_n420_), .A3(new_n424_), .A4(new_n373_), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT105), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n438_), .A2(new_n441_), .ZN(new_n442_));
  AOI211_X1 g241(.A(KEYINPUT104), .B(new_n425_), .C1(new_n380_), .C2(new_n392_), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n427_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n297_), .B(KEYINPUT30), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(new_n346_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G15gat), .B(G43gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G227gat), .A2(G233gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n446_), .B(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G71gat), .B(G99gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT90), .B(KEYINPUT31), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  XOR2_X1   g252(.A(new_n450_), .B(new_n453_), .Z(new_n454_));
  INV_X1    g253(.A(KEYINPUT91), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT106), .B1(new_n444_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n439_), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n454_), .A2(new_n426_), .A3(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n374_), .A2(new_n379_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n393_), .A2(new_n426_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT104), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n393_), .A2(new_n202_), .A3(new_n426_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n463_), .A2(new_n464_), .A3(new_n441_), .A4(new_n438_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n454_), .B(KEYINPUT91), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT106), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n457_), .A2(new_n461_), .A3(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G127gat), .B(G155gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(G211gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT16), .B(G183gat), .ZN(new_n473_));
  XOR2_X1   g272(.A(new_n472_), .B(new_n473_), .Z(new_n474_));
  INV_X1    g273(.A(KEYINPUT17), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT76), .B(G15gat), .ZN(new_n477_));
  INV_X1    g276(.A(G22gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(KEYINPUT77), .B(G8gat), .ZN(new_n480_));
  INV_X1    g279(.A(G1gat), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT14), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n479_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(G8gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT78), .B(G1gat), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n484_), .B(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G231gat), .A2(G233gat), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n488_), .B(KEYINPUT79), .Z(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n484_), .B(new_n485_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n489_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(G57gat), .B(G64gat), .Z(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n495_), .A2(KEYINPUT11), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n495_), .A2(KEYINPUT11), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G71gat), .B(G78gat), .ZN(new_n498_));
  OR3_X1    g297(.A1(new_n496_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n495_), .A2(new_n498_), .A3(KEYINPUT11), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n490_), .A2(new_n493_), .A3(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n502_), .B1(new_n490_), .B2(new_n493_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n476_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n505_), .A2(KEYINPUT80), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(KEYINPUT80), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n474_), .A2(new_n475_), .ZN(new_n508_));
  NOR3_X1   g307(.A1(new_n503_), .A2(new_n504_), .A3(new_n476_), .ZN(new_n509_));
  AOI22_X1  g308(.A1(new_n506_), .A2(new_n507_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G99gat), .A2(G106gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT69), .ZN(new_n513_));
  XNOR2_X1  g312(.A(KEYINPUT68), .B(KEYINPUT6), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT69), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n512_), .B(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n514_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT7), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT67), .ZN(new_n521_));
  NOR2_X1   g320(.A1(G99gat), .A2(G106gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n515_), .A2(new_n519_), .A3(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G85gat), .B(G92gat), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT70), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT70), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n524_), .A2(new_n529_), .A3(new_n526_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n528_), .A2(KEYINPUT8), .A3(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n512_), .B(KEYINPUT6), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n523_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT8), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(new_n534_), .A3(new_n526_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n531_), .A2(new_n535_), .ZN(new_n536_));
  OR2_X1    g335(.A1(KEYINPUT66), .A2(G85gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(KEYINPUT66), .A2(G85gat), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n537_), .B1(KEYINPUT9), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(G92gat), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n540_), .A2(new_n532_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(KEYINPUT10), .B(G99gat), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n542_), .A2(G106gat), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n543_), .A2(KEYINPUT65), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n526_), .A2(KEYINPUT9), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(KEYINPUT65), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n541_), .A2(new_n544_), .A3(new_n545_), .A4(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n536_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G43gat), .B(G50gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(G36gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT75), .B(G29gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT15), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n548_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n547_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n555_), .B1(new_n531_), .B2(new_n535_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(new_n552_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G232gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT34), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n554_), .B(new_n557_), .C1(KEYINPUT35), .C2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(KEYINPUT35), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n563_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT36), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G190gat), .B(G218gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G134gat), .B(G162gat), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n567_), .B(new_n568_), .Z(new_n569_));
  AOI22_X1  g368(.A1(new_n564_), .A2(new_n565_), .B1(new_n566_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT37), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n569_), .B(KEYINPUT36), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n564_), .A2(new_n565_), .A3(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n571_), .A2(new_n572_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n575_), .ZN(new_n577_));
  OAI21_X1  g376(.A(KEYINPUT37), .B1(new_n577_), .B2(new_n570_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  NOR3_X1   g378(.A1(new_n470_), .A2(new_n511_), .A3(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n548_), .A2(new_n502_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT71), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n582_), .B1(new_n556_), .B2(new_n501_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n581_), .A2(new_n583_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G230gat), .A2(G233gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT64), .ZN(new_n587_));
  NOR3_X1   g386(.A1(new_n584_), .A2(new_n585_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n587_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT12), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n590_), .B1(new_n556_), .B2(new_n501_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n581_), .A2(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n548_), .A2(new_n590_), .A3(new_n502_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n589_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G176gat), .B(G204gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G120gat), .B(G148gat), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n597_), .B(new_n598_), .Z(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  OR3_X1    g399(.A1(new_n588_), .A2(new_n594_), .A3(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n600_), .B1(new_n588_), .B2(new_n594_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n601_), .A2(KEYINPUT13), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(KEYINPUT13), .B1(new_n601_), .B2(new_n602_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n491_), .A2(new_n552_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n487_), .A2(new_n553_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G229gat), .A2(G233gat), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n552_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n487_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n608_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n611_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G113gat), .B(G141gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(new_n260_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(KEYINPUT81), .B(G169gat), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n619_), .B(new_n620_), .Z(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n612_), .A2(new_n617_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n622_), .B1(new_n612_), .B2(new_n617_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n607_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n580_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n460_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(new_n481_), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT38), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n571_), .A2(new_n575_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n469_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT107), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n469_), .A2(KEYINPUT107), .A3(new_n635_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n638_), .A2(new_n627_), .A3(new_n510_), .A4(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G1gat), .B1(new_n640_), .B2(new_n460_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n631_), .A2(new_n632_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n633_), .A2(new_n641_), .A3(new_n642_), .ZN(G1324gat));
  XNOR2_X1  g442(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n644_));
  INV_X1    g443(.A(new_n639_), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT107), .B1(new_n469_), .B2(new_n635_), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n645_), .A2(new_n646_), .A3(new_n511_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n647_), .A2(KEYINPUT108), .A3(new_n627_), .A4(new_n439_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT108), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n649_), .B1(new_n640_), .B2(new_n458_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n648_), .A2(new_n650_), .A3(G8gat), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(KEYINPUT39), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT39), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n648_), .A2(new_n650_), .A3(new_n653_), .A4(G8gat), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n629_), .A2(new_n480_), .A3(new_n439_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n644_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n644_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n656_), .ZN(new_n659_));
  AOI211_X1 g458(.A(new_n658_), .B(new_n659_), .C1(new_n652_), .C2(new_n654_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n657_), .A2(new_n660_), .ZN(G1325gat));
  OR3_X1    g460(.A1(new_n628_), .A2(G15gat), .A3(new_n466_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n647_), .A2(new_n627_), .A3(new_n456_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n663_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT41), .B1(new_n663_), .B2(G15gat), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n662_), .B1(new_n665_), .B2(new_n666_), .ZN(G1326gat));
  NAND3_X1  g466(.A1(new_n629_), .A2(new_n478_), .A3(new_n425_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n647_), .A2(new_n627_), .A3(new_n425_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n669_), .A2(new_n670_), .A3(G22gat), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n670_), .B1(new_n669_), .B2(G22gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n668_), .B1(new_n672_), .B2(new_n673_), .ZN(G1327gat));
  NAND2_X1  g473(.A1(new_n469_), .A2(new_n579_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n675_), .A2(KEYINPUT43), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n677_), .B1(new_n469_), .B2(new_n579_), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n676_), .A2(new_n678_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n607_), .A2(new_n626_), .A3(new_n510_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n679_), .A2(KEYINPUT44), .A3(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n680_), .B1(new_n676_), .B2(new_n678_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  AND4_X1   g483(.A1(G29gat), .A2(new_n681_), .A3(new_n630_), .A4(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n470_), .A2(new_n635_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n686_), .A2(new_n680_), .ZN(new_n687_));
  AOI21_X1  g486(.A(G29gat), .B1(new_n687_), .B2(new_n630_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n685_), .A2(new_n688_), .ZN(G1328gat));
  NAND3_X1  g488(.A1(new_n681_), .A2(new_n439_), .A3(new_n684_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(G36gat), .ZN(new_n691_));
  INV_X1    g490(.A(G36gat), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n439_), .B(KEYINPUT110), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n687_), .A2(new_n692_), .A3(new_n693_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT45), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n691_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT46), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n696_), .B(new_n697_), .ZN(G1329gat));
  NAND3_X1  g497(.A1(new_n681_), .A2(new_n454_), .A3(new_n684_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n466_), .A2(G43gat), .ZN(new_n700_));
  AOI22_X1  g499(.A1(new_n699_), .A2(G43gat), .B1(new_n687_), .B2(new_n700_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g501(.A1(new_n681_), .A2(new_n425_), .A3(new_n684_), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n703_), .A2(KEYINPUT111), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(KEYINPUT111), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(G50gat), .A3(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(G50gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n687_), .A2(new_n707_), .A3(new_n425_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(G1331gat));
  INV_X1    g508(.A(new_n626_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n606_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n580_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT112), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n460_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n580_), .A2(KEYINPUT112), .A3(new_n711_), .ZN(new_n715_));
  AOI21_X1  g514(.A(G57gat), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n638_), .A2(new_n510_), .A3(new_n639_), .A4(new_n711_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n630_), .A2(G57gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n716_), .B1(new_n718_), .B2(new_n719_), .ZN(G1332gat));
  INV_X1    g519(.A(new_n693_), .ZN(new_n721_));
  OR3_X1    g520(.A1(new_n712_), .A2(G64gat), .A3(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n718_), .A2(new_n693_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT48), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n723_), .A2(new_n724_), .A3(G64gat), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n724_), .B1(new_n723_), .B2(G64gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n722_), .B1(new_n726_), .B2(new_n727_), .ZN(G1333gat));
  OR3_X1    g527(.A1(new_n712_), .A2(G71gat), .A3(new_n466_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n718_), .A2(new_n456_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT49), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n731_), .A3(G71gat), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n731_), .B1(new_n730_), .B2(G71gat), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n729_), .B1(new_n733_), .B2(new_n734_), .ZN(G1334gat));
  OR3_X1    g534(.A1(new_n712_), .A2(G78gat), .A3(new_n426_), .ZN(new_n736_));
  OAI21_X1  g535(.A(G78gat), .B1(new_n717_), .B2(new_n426_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(KEYINPUT113), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT50), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT113), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n740_), .B(G78gat), .C1(new_n717_), .C2(new_n426_), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n738_), .A2(new_n739_), .A3(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n739_), .B1(new_n738_), .B2(new_n741_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n736_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT114), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT114), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n736_), .B(new_n746_), .C1(new_n742_), .C2(new_n743_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(G1335gat));
  NOR3_X1   g547(.A1(new_n606_), .A2(new_n710_), .A3(new_n510_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n686_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(G85gat), .B1(new_n751_), .B2(new_n630_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n679_), .A2(new_n749_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n460_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n752_), .B1(new_n753_), .B2(new_n754_), .ZN(G1336gat));
  AOI21_X1  g554(.A(G92gat), .B1(new_n751_), .B2(new_n439_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n693_), .A2(G92gat), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n753_), .B2(new_n757_), .ZN(G1337gat));
  NAND3_X1  g557(.A1(new_n679_), .A2(new_n456_), .A3(new_n749_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n542_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n454_), .A2(new_n760_), .ZN(new_n761_));
  AOI22_X1  g560(.A1(new_n759_), .A2(G99gat), .B1(new_n751_), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT115), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n763_), .A2(KEYINPUT51), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n762_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(KEYINPUT51), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n765_), .B(new_n766_), .Z(G1338gat));
  OR3_X1    g566(.A1(new_n750_), .A2(G106gat), .A3(new_n426_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n679_), .A2(new_n425_), .A3(new_n749_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n769_), .A2(new_n770_), .A3(G106gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n769_), .B2(G106gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g573(.A1(new_n615_), .A2(new_n611_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT119), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n776_), .A3(new_n621_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n616_), .B1(new_n608_), .B2(new_n614_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT119), .B1(new_n778_), .B2(new_n622_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n610_), .A2(new_n616_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n777_), .A2(new_n779_), .A3(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT120), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT120), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n777_), .A2(new_n779_), .A3(new_n783_), .A4(new_n780_), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n782_), .A2(new_n623_), .A3(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n601_), .A2(new_n602_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n592_), .A2(new_n589_), .A3(new_n593_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n594_), .B1(KEYINPUT55), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n592_), .A2(new_n593_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n790_), .A2(KEYINPUT55), .A3(new_n587_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  OAI211_X1 g591(.A(KEYINPUT56), .B(new_n600_), .C1(new_n789_), .C2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n788_), .A2(KEYINPUT55), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n790_), .A2(new_n587_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n791_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT56), .B1(new_n799_), .B2(new_n600_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n710_), .B1(new_n795_), .B2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n600_), .B1(new_n789_), .B2(new_n792_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT56), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(KEYINPUT118), .A3(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n601_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n787_), .B1(new_n801_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n635_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n601_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n793_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT121), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n810_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n802_), .A2(new_n803_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n814_), .A2(KEYINPUT121), .A3(new_n793_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n813_), .A2(new_n815_), .A3(new_n785_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT58), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n813_), .A2(new_n815_), .A3(KEYINPUT58), .A4(new_n785_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n579_), .A3(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n806_), .A2(KEYINPUT57), .A3(new_n635_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n809_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n511_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT117), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n510_), .A2(KEYINPUT116), .A3(new_n626_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT116), .B1(new_n510_), .B2(new_n626_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n605_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n829_), .A2(new_n603_), .A3(new_n576_), .A4(new_n578_), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n824_), .B(new_n825_), .C1(new_n828_), .C2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n827_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n510_), .A2(KEYINPUT116), .A3(new_n626_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n579_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(KEYINPUT117), .A2(KEYINPUT54), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n824_), .A2(new_n825_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n834_), .A2(new_n835_), .A3(new_n836_), .A4(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n831_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT122), .B1(new_n823_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT122), .ZN(new_n842_));
  AOI211_X1 g641(.A(new_n842_), .B(new_n839_), .C1(new_n822_), .C2(new_n511_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n841_), .A2(new_n843_), .A3(new_n460_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n459_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT59), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n823_), .A2(new_n840_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT59), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n847_), .A2(new_n848_), .A3(new_n630_), .A4(new_n459_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n846_), .A2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(G113gat), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n626_), .A2(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n844_), .A2(new_n710_), .A3(new_n459_), .ZN(new_n853_));
  AOI22_X1  g652(.A1(new_n850_), .A2(new_n852_), .B1(new_n851_), .B2(new_n853_), .ZN(G1340gat));
  NOR2_X1   g653(.A1(new_n606_), .A2(G120gat), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n844_), .B(new_n459_), .C1(KEYINPUT60), .C2(new_n855_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n846_), .A2(new_n607_), .A3(new_n856_), .A4(new_n849_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(G120gat), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n856_), .A2(KEYINPUT60), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(G1341gat));
  NAND2_X1  g659(.A1(new_n510_), .A2(G127gat), .ZN(new_n861_));
  XOR2_X1   g660(.A(new_n861_), .B(KEYINPUT123), .Z(new_n862_));
  INV_X1    g661(.A(G127gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n844_), .A2(new_n510_), .A3(new_n459_), .ZN(new_n864_));
  AOI22_X1  g663(.A1(new_n850_), .A2(new_n862_), .B1(new_n863_), .B2(new_n864_), .ZN(G1342gat));
  INV_X1    g664(.A(new_n579_), .ZN(new_n866_));
  INV_X1    g665(.A(G134gat), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n844_), .A2(new_n634_), .A3(new_n459_), .ZN(new_n869_));
  AOI22_X1  g668(.A1(new_n850_), .A2(new_n868_), .B1(new_n867_), .B2(new_n869_), .ZN(G1343gat));
  NOR2_X1   g669(.A1(new_n456_), .A2(new_n426_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n844_), .A2(new_n721_), .A3(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n872_), .A2(new_n626_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(new_n326_), .ZN(G1344gat));
  NOR2_X1   g673(.A1(new_n872_), .A2(new_n606_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(new_n327_), .ZN(G1345gat));
  AND2_X1   g675(.A1(new_n844_), .A2(new_n721_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n877_), .A2(new_n510_), .A3(new_n871_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(KEYINPUT61), .B(G155gat), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(G1346gat));
  INV_X1    g679(.A(G162gat), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n872_), .A2(new_n881_), .A3(new_n866_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n877_), .A2(new_n634_), .A3(new_n871_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n881_), .B2(new_n883_), .ZN(G1347gat));
  NOR2_X1   g683(.A1(new_n721_), .A2(new_n630_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n885_), .A2(new_n456_), .A3(new_n426_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n847_), .A2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n229_), .B1(new_n889_), .B2(new_n710_), .ZN(new_n890_));
  OR2_X1    g689(.A1(new_n890_), .A2(KEYINPUT62), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n889_), .A2(new_n710_), .A3(new_n277_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(KEYINPUT62), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n891_), .A2(new_n892_), .A3(new_n893_), .ZN(G1348gat));
  OAI21_X1  g693(.A(new_n230_), .B1(new_n888_), .B2(new_n606_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n841_), .A2(new_n843_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n896_), .A2(G176gat), .A3(new_n607_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n895_), .B1(new_n897_), .B2(new_n886_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(KEYINPUT124), .ZN(G1349gat));
  NOR3_X1   g698(.A1(new_n888_), .A2(new_n511_), .A3(new_n282_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n896_), .A2(new_n510_), .A3(new_n887_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n227_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n900_), .B1(new_n901_), .B2(new_n902_), .ZN(G1350gat));
  OAI21_X1  g702(.A(G190gat), .B1(new_n888_), .B2(new_n866_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n634_), .A2(new_n283_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n888_), .B2(new_n905_), .ZN(G1351gat));
  NAND2_X1  g705(.A1(new_n847_), .A2(new_n842_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n823_), .A2(KEYINPUT122), .A3(new_n840_), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n907_), .A2(new_n908_), .A3(new_n871_), .A4(new_n885_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT125), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n896_), .A2(KEYINPUT125), .A3(new_n871_), .A4(new_n885_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n626_), .B1(new_n911_), .B2(new_n912_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(new_n260_), .ZN(G1352gat));
  AOI21_X1  g713(.A(new_n606_), .B1(new_n911_), .B2(new_n912_), .ZN(new_n915_));
  AND2_X1   g714(.A1(new_n258_), .A2(KEYINPUT126), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n258_), .A2(KEYINPUT126), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n915_), .B1(new_n916_), .B2(new_n917_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n918_), .B1(new_n915_), .B2(new_n916_), .ZN(G1353gat));
  NAND2_X1  g718(.A1(new_n911_), .A2(new_n912_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(KEYINPUT127), .ZN(new_n922_));
  NAND2_X1  g721(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n923_));
  AND4_X1   g722(.A1(new_n510_), .A2(new_n920_), .A3(new_n922_), .A4(new_n923_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n511_), .B1(new_n911_), .B2(new_n912_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n922_), .B1(new_n925_), .B2(new_n923_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n924_), .A2(new_n926_), .ZN(G1354gat));
  AOI21_X1  g726(.A(G218gat), .B1(new_n920_), .B2(new_n634_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n866_), .B1(new_n911_), .B2(new_n912_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n928_), .B1(G218gat), .B2(new_n929_), .ZN(G1355gat));
endmodule


