//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1 1 0 1 0 0 0 0 0 1 1 1 1 0 0 0 1 1 0 0 0 0 1 0 0 0 0 1 0 0 1 0 1 0 0 1 1 0 1 1 0 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n837_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n877_, new_n878_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n903_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  OAI21_X1  g002(.A(new_n203_), .B1(G183gat), .B2(G190gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n205_));
  OR3_X1    g004(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT24), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n203_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT81), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G169gat), .ZN(new_n214_));
  INV_X1    g013(.A(G176gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT24), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n216_), .A2(new_n208_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT26), .B(G190gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT80), .ZN(new_n219_));
  INV_X1    g018(.A(G183gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n219_), .B1(new_n220_), .B2(KEYINPUT25), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT25), .B(G183gat), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n218_), .B(new_n221_), .C1(new_n222_), .C2(new_n219_), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n217_), .B(new_n223_), .C1(new_n211_), .C2(KEYINPUT81), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n207_), .B1(new_n213_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(G204gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT88), .B1(new_n226_), .B2(G197gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT88), .ZN(new_n228_));
  INV_X1    g027(.A(G197gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(new_n229_), .A3(G204gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n226_), .A2(G197gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n227_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n232_), .A2(KEYINPUT21), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G211gat), .B(G218gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n229_), .A2(G204gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(new_n231_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n236_), .A2(KEYINPUT87), .A3(KEYINPUT21), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(KEYINPUT21), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT87), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n233_), .A2(new_n234_), .A3(new_n237_), .A4(new_n240_), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n232_), .A2(KEYINPUT89), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n232_), .A2(KEYINPUT89), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT21), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n234_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n242_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n241_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n225_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G226gat), .A2(G233gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n211_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT93), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n208_), .B1(new_n216_), .B2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n254_), .B1(new_n253_), .B2(new_n216_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT92), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n222_), .B(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n218_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n252_), .B(new_n255_), .C1(new_n257_), .C2(new_n258_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n259_), .A2(new_n246_), .A3(new_n241_), .A4(new_n207_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n248_), .A2(KEYINPUT20), .A3(new_n251_), .A4(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT95), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n260_), .A2(KEYINPUT20), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n264_), .A2(KEYINPUT95), .A3(new_n251_), .A4(new_n248_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G8gat), .B(G36gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT18), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G64gat), .B(G92gat), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n268_), .B(new_n269_), .Z(new_n270_));
  OR2_X1    g069(.A1(new_n213_), .A2(new_n224_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n271_), .A2(new_n246_), .A3(new_n241_), .A4(new_n207_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT20), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n259_), .A2(new_n207_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n273_), .B1(new_n274_), .B2(new_n247_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n251_), .B1(new_n272_), .B2(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n276_), .A2(KEYINPUT94), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT94), .ZN(new_n278_));
  AOI211_X1 g077(.A(new_n278_), .B(new_n251_), .C1(new_n272_), .C2(new_n275_), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n266_), .B(new_n270_), .C1(new_n277_), .C2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT27), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n272_), .A2(new_n275_), .A3(new_n251_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n248_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n260_), .A2(KEYINPUT20), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n282_), .B1(new_n285_), .B2(new_n251_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n270_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n281_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n280_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n280_), .A2(KEYINPUT96), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n276_), .B(KEYINPUT94), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT96), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n291_), .A2(new_n292_), .A3(new_n270_), .A4(new_n266_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n277_), .A2(new_n279_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n266_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n287_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n290_), .A2(new_n293_), .A3(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n289_), .B1(new_n297_), .B2(new_n281_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G227gat), .A2(G233gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT83), .ZN(new_n300_));
  XOR2_X1   g099(.A(G71gat), .B(G99gat), .Z(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n225_), .B(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(G127gat), .B(G134gat), .Z(new_n304_));
  XOR2_X1   g103(.A(G113gat), .B(G120gat), .Z(new_n305_));
  XOR2_X1   g104(.A(new_n304_), .B(new_n305_), .Z(new_n306_));
  XNOR2_X1  g105(.A(new_n303_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G15gat), .B(G43gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT82), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT30), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT31), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n307_), .B(new_n311_), .Z(new_n312_));
  NAND2_X1  g111(.A1(G225gat), .A2(G233gat), .ZN(new_n313_));
  INV_X1    g112(.A(new_n306_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G141gat), .A2(G148gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(G141gat), .A2(G148gat), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n316_), .A2(KEYINPUT84), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(KEYINPUT84), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n315_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320_));
  NOR2_X1   g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n320_), .B1(new_n321_), .B2(KEYINPUT1), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n322_), .A2(KEYINPUT85), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n320_), .A2(KEYINPUT1), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n324_), .B1(new_n322_), .B2(KEYINPUT85), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n319_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n316_), .B(KEYINPUT3), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n315_), .B(KEYINPUT2), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT86), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT86), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n328_), .A2(new_n332_), .A3(new_n329_), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n321_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(new_n320_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n314_), .B(new_n327_), .C1(new_n334_), .C2(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n336_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n306_), .B1(new_n338_), .B2(new_n326_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(KEYINPUT4), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT4), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n341_), .B(new_n306_), .C1(new_n338_), .C2(new_n326_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n313_), .B1(new_n340_), .B2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G1gat), .B(G29gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(G85gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT0), .B(G57gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n345_), .B(new_n346_), .Z(new_n347_));
  INV_X1    g146(.A(new_n313_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n348_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n349_));
  OR3_X1    g148(.A1(new_n343_), .A2(new_n347_), .A3(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n347_), .B1(new_n343_), .B2(new_n349_), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n350_), .A2(KEYINPUT99), .A3(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(KEYINPUT99), .B1(new_n350_), .B2(new_n351_), .ZN(new_n353_));
  NOR3_X1   g152(.A1(new_n312_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n338_), .A2(new_n326_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT29), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n247_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G228gat), .A2(G233gat), .ZN(new_n358_));
  INV_X1    g157(.A(G78gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(G106gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n357_), .B(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT90), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT28), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n366_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NOR4_X1   g167(.A1(new_n338_), .A2(new_n326_), .A3(KEYINPUT28), .A4(KEYINPUT29), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G22gat), .B(G50gat), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n368_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n371_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n373_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n364_), .A2(new_n365_), .A3(new_n372_), .A4(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n372_), .A2(new_n365_), .A3(new_n374_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n357_), .B(new_n362_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n365_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n375_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n298_), .A2(new_n354_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n350_), .A2(new_n351_), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n270_), .A2(KEYINPUT32), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n286_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n291_), .A2(new_n266_), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n382_), .B(new_n384_), .C1(new_n385_), .C2(new_n383_), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n351_), .A2(KEYINPUT97), .A3(KEYINPUT33), .ZN(new_n387_));
  AOI21_X1  g186(.A(KEYINPUT33), .B1(new_n351_), .B2(KEYINPUT97), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n337_), .A2(new_n348_), .A3(new_n339_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n347_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n389_), .A2(KEYINPUT98), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n340_), .A2(new_n342_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n391_), .B1(new_n348_), .B2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(KEYINPUT98), .B1(new_n389_), .B2(new_n390_), .ZN(new_n394_));
  OAI22_X1  g193(.A1(new_n387_), .A2(new_n388_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n386_), .B1(new_n395_), .B2(new_n297_), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n352_), .A2(new_n380_), .A3(new_n353_), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n396_), .A2(new_n380_), .B1(new_n298_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n312_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n381_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G113gat), .B(G141gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G169gat), .B(G197gat), .ZN(new_n402_));
  XOR2_X1   g201(.A(new_n401_), .B(new_n402_), .Z(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G229gat), .A2(G233gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G29gat), .B(G36gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT74), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT75), .ZN(new_n408_));
  OR2_X1    g207(.A1(new_n406_), .A2(KEYINPUT74), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT75), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n406_), .A2(KEYINPUT74), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n409_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G43gat), .B(G50gat), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n408_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n413_), .B1(new_n408_), .B2(new_n412_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G15gat), .B(G22gat), .ZN(new_n418_));
  INV_X1    g217(.A(G1gat), .ZN(new_n419_));
  INV_X1    g218(.A(G8gat), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT14), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n418_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G1gat), .B(G8gat), .ZN(new_n423_));
  XOR2_X1   g222(.A(new_n422_), .B(new_n423_), .Z(new_n424_));
  NOR2_X1   g223(.A1(new_n417_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n417_), .A2(new_n424_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n405_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n405_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT15), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n430_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n416_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n432_), .A2(KEYINPUT15), .A3(new_n414_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n424_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n429_), .A2(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n404_), .B1(new_n428_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n432_), .A2(new_n414_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(new_n424_), .ZN(new_n438_));
  OAI221_X1 g237(.A(new_n403_), .B1(new_n429_), .B2(new_n434_), .C1(new_n438_), .C2(new_n405_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n436_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G230gat), .A2(G233gat), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT66), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  OAI211_X1 g245(.A(KEYINPUT66), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G99gat), .A2(G106gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT6), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT6), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n451_), .A2(G99gat), .A3(G106gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  OR2_X1    g252(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n454_));
  INV_X1    g253(.A(G99gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n454_), .A2(new_n455_), .A3(new_n361_), .A4(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n448_), .A2(new_n453_), .A3(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT68), .ZN(new_n459_));
  AND2_X1   g258(.A1(G85gat), .A2(G92gat), .ZN(new_n460_));
  NOR2_X1   g259(.A1(G85gat), .A2(G92gat), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n459_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(G85gat), .ZN(new_n463_));
  INV_X1    g262(.A(G92gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G85gat), .A2(G92gat), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(KEYINPUT68), .A3(new_n466_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n462_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n458_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT8), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT65), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n451_), .B1(G99gat), .B2(G106gat), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n449_), .A2(KEYINPUT6), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n471_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n450_), .A2(new_n452_), .A3(KEYINPUT65), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n474_), .A2(new_n475_), .A3(new_n448_), .A4(new_n457_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT8), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n462_), .A2(new_n467_), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n470_), .A2(new_n479_), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n450_), .A2(new_n452_), .A3(KEYINPUT65), .ZN(new_n481_));
  AOI21_X1  g280(.A(KEYINPUT65), .B1(new_n450_), .B2(new_n452_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT10), .B(G99gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT64), .B(G106gat), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n465_), .A2(KEYINPUT9), .A3(new_n466_), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n466_), .A2(KEYINPUT9), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n483_), .A2(new_n486_), .A3(new_n489_), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n480_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G57gat), .B(G64gat), .ZN(new_n492_));
  OR2_X1    g291(.A1(new_n492_), .A2(KEYINPUT11), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(KEYINPUT11), .ZN(new_n494_));
  XOR2_X1   g293(.A(G71gat), .B(G78gat), .Z(new_n495_));
  NAND3_X1  g294(.A1(new_n493_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n496_));
  OR2_X1    g295(.A1(new_n494_), .A2(new_n495_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n491_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n480_), .A2(new_n490_), .A3(new_n498_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n443_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT69), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT69), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n504_), .B(new_n443_), .C1(new_n499_), .C2(new_n501_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n498_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT12), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT71), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n483_), .A2(KEYINPUT70), .A3(new_n486_), .A4(new_n489_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT70), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n474_), .A2(new_n475_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n487_), .B(new_n488_), .C1(new_n484_), .C2(new_n485_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n512_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n511_), .A2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n510_), .B1(new_n516_), .B2(new_n480_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n511_), .A2(new_n515_), .ZN(new_n518_));
  AOI22_X1  g317(.A1(new_n469_), .A2(KEYINPUT8), .B1(new_n476_), .B2(new_n478_), .ZN(new_n519_));
  NOR3_X1   g318(.A1(new_n518_), .A2(new_n519_), .A3(KEYINPUT71), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n509_), .B1(new_n517_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n480_), .A2(new_n490_), .ZN(new_n522_));
  AOI21_X1  g321(.A(KEYINPUT12), .B1(new_n522_), .B2(new_n507_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n500_), .A2(new_n442_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n521_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n506_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G120gat), .B(G148gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT5), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G176gat), .B(G204gat), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n529_), .B(new_n530_), .Z(new_n531_));
  NAND2_X1  g330(.A1(new_n527_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n531_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n506_), .A2(new_n526_), .A3(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT13), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n532_), .B(new_n534_), .C1(KEYINPUT72), .C2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT73), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT73), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n537_), .A2(new_n542_), .A3(new_n539_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n441_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT77), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT76), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G232gat), .A2(G233gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT34), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT35), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n516_), .A2(new_n510_), .A3(new_n480_), .ZN(new_n550_));
  OAI21_X1  g349(.A(KEYINPUT71), .B1(new_n518_), .B2(new_n519_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n431_), .A2(new_n433_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n548_), .A2(KEYINPUT76), .A3(KEYINPUT35), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n548_), .A2(KEYINPUT35), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n553_), .B(new_n554_), .C1(new_n437_), .C2(new_n522_), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n546_), .B(new_n549_), .C1(new_n552_), .C2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n555_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n431_), .A2(new_n433_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n550_), .A2(new_n551_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n549_), .A2(new_n546_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n557_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G190gat), .B(G218gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G134gat), .B(G162gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n565_), .B(KEYINPUT36), .Z(new_n566_));
  AND3_X1   g365(.A1(new_n556_), .A2(new_n562_), .A3(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n565_), .A2(KEYINPUT36), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n569_), .B1(new_n556_), .B2(new_n562_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n545_), .B1(new_n567_), .B2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n556_), .A2(new_n562_), .A3(new_n566_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT77), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT78), .B(KEYINPUT37), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n571_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT37), .B1(new_n567_), .B2(new_n570_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n424_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(new_n498_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT79), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G127gat), .B(G155gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT16), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G183gat), .B(G211gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT17), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n582_), .B(new_n587_), .ZN(new_n588_));
  OR3_X1    g387(.A1(new_n581_), .A2(KEYINPUT17), .A3(new_n586_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n578_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n400_), .A2(new_n544_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n352_), .A2(new_n353_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n593_), .A2(new_n419_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT38), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT100), .Z(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(new_n597_), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n600_), .B(KEYINPUT101), .Z(new_n601_));
  NAND2_X1  g400(.A1(new_n571_), .A2(new_n573_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n400_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n590_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n544_), .A2(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(G1gat), .B1(new_n607_), .B2(new_n594_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n599_), .A2(new_n601_), .A3(new_n608_), .ZN(G1324gat));
  INV_X1    g408(.A(new_n298_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n593_), .A2(new_n420_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT39), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n606_), .A2(new_n610_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n612_), .B1(new_n613_), .B2(G8gat), .ZN(new_n614_));
  AOI211_X1 g413(.A(KEYINPUT39), .B(new_n420_), .C1(new_n606_), .C2(new_n610_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n611_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT40), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(G1325gat));
  OR3_X1    g417(.A1(new_n592_), .A2(G15gat), .A3(new_n312_), .ZN(new_n619_));
  OAI21_X1  g418(.A(G15gat), .B1(new_n607_), .B2(new_n312_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT41), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n620_), .A2(new_n621_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n619_), .B1(new_n622_), .B2(new_n623_), .ZN(G1326gat));
  XOR2_X1   g423(.A(new_n380_), .B(KEYINPUT102), .Z(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  OR3_X1    g425(.A1(new_n592_), .A2(G22gat), .A3(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(G22gat), .B1(new_n607_), .B2(new_n626_), .ZN(new_n628_));
  XOR2_X1   g427(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n629_));
  AND2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n628_), .A2(new_n629_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n627_), .B1(new_n630_), .B2(new_n631_), .ZN(G1327gat));
  AND2_X1   g431(.A1(new_n544_), .A2(new_n590_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT43), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n396_), .A2(new_n380_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n298_), .A2(new_n397_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n399_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n381_), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n634_), .B(new_n578_), .C1(new_n637_), .C2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n634_), .B1(new_n400_), .B2(new_n578_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n633_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT44), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  OAI211_X1 g443(.A(KEYINPUT44), .B(new_n633_), .C1(new_n640_), .C2(new_n641_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n646_), .A2(new_n595_), .ZN(new_n647_));
  INV_X1    g446(.A(G29gat), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n604_), .A2(new_n602_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n400_), .A2(new_n544_), .A3(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n594_), .A2(G29gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT104), .ZN(new_n652_));
  OAI22_X1  g451(.A1(new_n647_), .A2(new_n648_), .B1(new_n650_), .B2(new_n652_), .ZN(G1328gat));
  OR2_X1    g452(.A1(new_n298_), .A2(G36gat), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n650_), .A2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT45), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n644_), .A2(new_n610_), .A3(new_n645_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n656_), .B1(new_n657_), .B2(G36gat), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT46), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n658_), .A2(KEYINPUT105), .A3(new_n659_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n659_), .A2(KEYINPUT105), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n659_), .A2(KEYINPUT105), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n658_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n660_), .A2(new_n663_), .ZN(G1329gat));
  NAND3_X1  g463(.A1(new_n646_), .A2(G43gat), .A3(new_n399_), .ZN(new_n665_));
  INV_X1    g464(.A(G43gat), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n666_), .B1(new_n650_), .B2(new_n312_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n665_), .A2(new_n667_), .A3(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n665_), .B2(new_n667_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1330gat));
  OR3_X1    g470(.A1(new_n650_), .A2(G50gat), .A3(new_n626_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT107), .ZN(new_n673_));
  INV_X1    g472(.A(new_n380_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n646_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(G50gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n673_), .B1(new_n646_), .B2(new_n674_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n672_), .B1(new_n676_), .B2(new_n677_), .ZN(G1331gat));
  NAND2_X1  g477(.A1(new_n541_), .A2(new_n543_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n679_), .A2(new_n590_), .A3(new_n440_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n603_), .A2(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G57gat), .B1(new_n681_), .B2(new_n594_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n679_), .A2(new_n440_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n683_), .A2(new_n591_), .A3(new_n400_), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n594_), .A2(G57gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n682_), .B1(new_n684_), .B2(new_n685_), .ZN(G1332gat));
  INV_X1    g485(.A(new_n684_), .ZN(new_n687_));
  INV_X1    g486(.A(G64gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(new_n688_), .A3(new_n610_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT48), .ZN(new_n690_));
  INV_X1    g489(.A(new_n681_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(new_n610_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n690_), .B1(new_n692_), .B2(G64gat), .ZN(new_n693_));
  AOI211_X1 g492(.A(KEYINPUT48), .B(new_n688_), .C1(new_n691_), .C2(new_n610_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n689_), .B1(new_n693_), .B2(new_n694_), .ZN(G1333gat));
  OAI21_X1  g494(.A(G71gat), .B1(new_n681_), .B2(new_n312_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n696_), .A2(KEYINPUT49), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n696_), .A2(KEYINPUT49), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n312_), .A2(G71gat), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT108), .Z(new_n700_));
  OAI22_X1  g499(.A1(new_n697_), .A2(new_n698_), .B1(new_n684_), .B2(new_n700_), .ZN(G1334gat));
  NAND3_X1  g500(.A1(new_n687_), .A2(new_n359_), .A3(new_n625_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n691_), .A2(new_n625_), .ZN(new_n703_));
  XOR2_X1   g502(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n704_));
  AND3_X1   g503(.A1(new_n703_), .A2(G78gat), .A3(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n703_), .B2(G78gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n702_), .B1(new_n705_), .B2(new_n706_), .ZN(G1335gat));
  OR2_X1    g506(.A1(new_n640_), .A2(new_n641_), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n679_), .A2(new_n604_), .A3(new_n440_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(G85gat), .B1(new_n710_), .B2(new_n594_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n683_), .A2(new_n400_), .A3(new_n649_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n595_), .A2(new_n463_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n711_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT110), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n714_), .B(new_n715_), .ZN(G1336gat));
  OAI21_X1  g515(.A(G92gat), .B1(new_n710_), .B2(new_n298_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n610_), .A2(new_n464_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n717_), .B1(new_n712_), .B2(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT111), .ZN(G1337gat));
  NOR3_X1   g519(.A1(new_n712_), .A2(new_n484_), .A3(new_n312_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT112), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n710_), .A2(new_n312_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(new_n455_), .B2(new_n723_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT51), .ZN(G1338gat));
  OR3_X1    g524(.A1(new_n712_), .A2(new_n485_), .A3(new_n380_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n708_), .A2(new_n674_), .A3(new_n709_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT52), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n727_), .A2(new_n728_), .A3(G106gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n727_), .B2(G106gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n726_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT53), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT53), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n733_), .B(new_n726_), .C1(new_n729_), .C2(new_n730_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(G1339gat));
  AOI21_X1  g534(.A(new_n440_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n591_), .A2(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n591_), .A2(new_n736_), .A3(new_n738_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT114), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT55), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n521_), .A2(new_n524_), .A3(new_n500_), .ZN(new_n745_));
  AOI22_X1  g544(.A1(new_n744_), .A2(new_n526_), .B1(new_n745_), .B2(new_n443_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n521_), .A2(KEYINPUT55), .A3(new_n524_), .A4(new_n525_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n533_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n743_), .B1(new_n748_), .B2(KEYINPUT56), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n745_), .A2(new_n443_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n526_), .A2(new_n744_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(new_n751_), .A3(new_n747_), .ZN(new_n752_));
  AOI21_X1  g551(.A(KEYINPUT56), .B1(new_n752_), .B2(new_n531_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT114), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n752_), .A2(KEYINPUT56), .A3(new_n531_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n749_), .A2(new_n754_), .A3(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n405_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n427_), .A2(new_n757_), .ZN(new_n758_));
  OAI221_X1 g557(.A(new_n404_), .B1(new_n758_), .B2(new_n434_), .C1(new_n438_), .C2(new_n757_), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n534_), .A2(new_n439_), .A3(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT58), .B1(new_n756_), .B2(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT115), .B1(new_n761_), .B2(new_n577_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n755_), .B1(new_n753_), .B2(KEYINPUT114), .ZN(new_n763_));
  AOI211_X1 g562(.A(new_n743_), .B(KEYINPUT56), .C1(new_n752_), .C2(new_n531_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n760_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT58), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT115), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n767_), .A2(new_n768_), .A3(new_n578_), .ZN(new_n769_));
  OAI211_X1 g568(.A(KEYINPUT58), .B(new_n760_), .C1(new_n763_), .C2(new_n764_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n762_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n440_), .A2(new_n534_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n753_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n773_), .B2(new_n755_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n759_), .A2(new_n439_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n775_), .B1(new_n532_), .B2(new_n534_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n602_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT57), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  OAI211_X1 g578(.A(KEYINPUT57), .B(new_n602_), .C1(new_n774_), .C2(new_n776_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n771_), .A2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT117), .B1(new_n782_), .B2(new_n590_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT117), .ZN(new_n784_));
  AOI211_X1 g583(.A(new_n784_), .B(new_n604_), .C1(new_n771_), .C2(new_n781_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n742_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n610_), .A2(new_n674_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n787_), .A2(new_n595_), .A3(new_n399_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n788_), .A2(KEYINPUT59), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n786_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT116), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n779_), .A2(new_n780_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n770_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n577_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n794_), .B2(new_n768_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n792_), .B1(new_n795_), .B2(new_n762_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n742_), .B1(new_n796_), .B2(new_n604_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n788_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n791_), .B1(new_n799_), .B2(KEYINPUT59), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT59), .ZN(new_n801_));
  AOI211_X1 g600(.A(KEYINPUT116), .B(new_n801_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n790_), .B(new_n440_), .C1(new_n800_), .C2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(G113gat), .ZN(new_n804_));
  OR3_X1    g603(.A1(new_n799_), .A2(G113gat), .A3(new_n441_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(G1340gat));
  INV_X1    g605(.A(new_n679_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n790_), .B(new_n807_), .C1(new_n800_), .C2(new_n802_), .ZN(new_n808_));
  XOR2_X1   g607(.A(KEYINPUT118), .B(G120gat), .Z(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n799_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n809_), .B1(new_n679_), .B2(KEYINPUT60), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n812_), .B(new_n813_), .C1(KEYINPUT60), .C2(new_n809_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n811_), .A2(new_n814_), .ZN(G1341gat));
  AOI21_X1  g614(.A(G127gat), .B1(new_n812_), .B2(new_n604_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n800_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n802_), .ZN(new_n818_));
  AOI22_X1  g617(.A1(new_n817_), .A2(new_n818_), .B1(new_n786_), .B2(new_n789_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n590_), .A2(KEYINPUT119), .ZN(new_n820_));
  MUX2_X1   g619(.A(KEYINPUT119), .B(new_n820_), .S(G127gat), .Z(new_n821_));
  AOI21_X1  g620(.A(new_n816_), .B1(new_n819_), .B2(new_n821_), .ZN(G1342gat));
  INV_X1    g621(.A(G134gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n799_), .B2(new_n602_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT120), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT120), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n826_), .B(new_n823_), .C1(new_n799_), .C2(new_n602_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n577_), .A2(new_n823_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n819_), .B2(new_n829_), .ZN(G1343gat));
  AOI22_X1  g629(.A1(new_n782_), .A2(new_n590_), .B1(new_n741_), .B2(new_n740_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n595_), .A2(new_n674_), .A3(new_n312_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n831_), .A2(new_n610_), .A3(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n440_), .ZN(new_n834_));
  XOR2_X1   g633(.A(KEYINPUT121), .B(G141gat), .Z(new_n835_));
  XNOR2_X1  g634(.A(new_n834_), .B(new_n835_), .ZN(G1344gat));
  NAND2_X1  g635(.A1(new_n833_), .A2(new_n807_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g637(.A1(new_n833_), .A2(new_n604_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(KEYINPUT61), .B(G155gat), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n839_), .B(new_n840_), .ZN(G1346gat));
  INV_X1    g640(.A(G162gat), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n833_), .A2(new_n842_), .A3(new_n571_), .A4(new_n573_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n833_), .A2(new_n578_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n843_), .B1(new_n845_), .B2(new_n842_), .ZN(G1347gat));
  AND2_X1   g645(.A1(new_n740_), .A2(new_n741_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n784_), .B1(new_n796_), .B2(new_n604_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n782_), .A2(KEYINPUT117), .A3(new_n590_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n847_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n610_), .A2(new_n354_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(KEYINPUT122), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n852_), .A2(new_n625_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n850_), .A2(new_n854_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT22), .B(G169gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(new_n440_), .A3(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n786_), .A2(new_n440_), .A3(new_n853_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n214_), .B1(KEYINPUT123), .B2(KEYINPUT62), .ZN(new_n859_));
  NOR2_X1   g658(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n858_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n857_), .B1(new_n861_), .B2(new_n862_), .ZN(G1348gat));
  INV_X1    g662(.A(KEYINPUT124), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n850_), .A2(new_n679_), .A3(new_n854_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(G176gat), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n786_), .A2(new_n807_), .A3(new_n853_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(KEYINPUT124), .A3(new_n215_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n831_), .A2(new_n674_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n852_), .A2(new_n679_), .A3(new_n215_), .ZN(new_n870_));
  AOI22_X1  g669(.A1(new_n866_), .A2(new_n868_), .B1(new_n869_), .B2(new_n870_), .ZN(G1349gat));
  AND2_X1   g670(.A1(new_n604_), .A2(new_n257_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n852_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n869_), .A2(new_n604_), .A3(new_n873_), .ZN(new_n874_));
  AOI22_X1  g673(.A1(new_n855_), .A2(new_n872_), .B1(new_n874_), .B2(new_n220_), .ZN(G1350gat));
  NAND4_X1  g674(.A1(new_n855_), .A2(new_n571_), .A3(new_n573_), .A4(new_n218_), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n850_), .A2(new_n577_), .A3(new_n854_), .ZN(new_n877_));
  INV_X1    g676(.A(G190gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n876_), .B1(new_n877_), .B2(new_n878_), .ZN(G1351gat));
  NAND3_X1  g678(.A1(new_n610_), .A2(new_n397_), .A3(new_n312_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n831_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n440_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n807_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(KEYINPUT125), .B2(G204gat), .ZN(new_n885_));
  XOR2_X1   g684(.A(KEYINPUT125), .B(G204gat), .Z(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n884_), .B2(new_n886_), .ZN(G1353gat));
  NAND2_X1  g686(.A1(new_n881_), .A2(new_n604_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT127), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n888_), .A2(KEYINPUT127), .A3(new_n889_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT126), .ZN(new_n894_));
  XOR2_X1   g693(.A(KEYINPUT63), .B(G211gat), .Z(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n894_), .B1(new_n888_), .B2(new_n896_), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n881_), .A2(KEYINPUT126), .A3(new_n604_), .A4(new_n895_), .ZN(new_n898_));
  AOI22_X1  g697(.A1(new_n892_), .A2(new_n893_), .B1(new_n897_), .B2(new_n898_), .ZN(G1354gat));
  INV_X1    g698(.A(G218gat), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n881_), .A2(new_n900_), .A3(new_n571_), .A4(new_n573_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n881_), .A2(new_n578_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n901_), .B1(new_n903_), .B2(new_n900_), .ZN(G1355gat));
endmodule


