//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 0 1 0 0 0 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 0 1 1 1 0 1 0 0 0 1 1 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n979_,
    new_n980_, new_n981_, new_n982_, new_n983_, new_n984_, new_n985_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n992_, new_n993_,
    new_n994_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_,
    new_n1001_, new_n1002_, new_n1003_, new_n1005_, new_n1006_, new_n1007_,
    new_n1009_, new_n1011_, new_n1012_, new_n1014_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1030_,
    new_n1031_, new_n1033_, new_n1034_, new_n1036_, new_n1037_, new_n1039_,
    new_n1040_, new_n1042_, new_n1044_, new_n1045_, new_n1046_, new_n1047_,
    new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT73), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n207_), .A2(KEYINPUT73), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n206_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(G1gat), .B(G8gat), .Z(new_n212_));
  INV_X1    g011(.A(KEYINPUT73), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n214_), .A2(new_n205_), .A3(new_n202_), .A4(new_n208_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n211_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G29gat), .B(G36gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  XOR2_X1   g017(.A(G43gat), .B(G50gat), .Z(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G43gat), .B(G50gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n217_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT70), .B(KEYINPUT15), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n220_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n220_), .A2(new_n222_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n223_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n216_), .A2(new_n224_), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT76), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G229gat), .A2(G233gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT76), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n216_), .A2(new_n231_), .A3(new_n224_), .A4(new_n227_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n211_), .A2(new_n215_), .A3(new_n225_), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n229_), .A2(new_n230_), .A3(new_n232_), .A4(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT77), .ZN(new_n235_));
  INV_X1    g034(.A(new_n233_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n236_), .B1(new_n228_), .B2(KEYINPUT76), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT77), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n237_), .A2(new_n238_), .A3(new_n230_), .A4(new_n232_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n230_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n225_), .B1(new_n211_), .B2(new_n215_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n240_), .B1(new_n236_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT75), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n225_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n216_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(new_n233_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n247_), .A2(KEYINPUT75), .A3(new_n240_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n244_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n235_), .A2(new_n239_), .A3(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G113gat), .B(G141gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G169gat), .B(G197gat), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n251_), .B(new_n252_), .Z(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n250_), .A2(new_n254_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n235_), .A2(new_n249_), .A3(new_n239_), .A4(new_n253_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT81), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G71gat), .B(G99gat), .ZN(new_n260_));
  INV_X1    g059(.A(G43gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT30), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G227gat), .A2(G233gat), .ZN(new_n264_));
  INV_X1    g063(.A(G15gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n263_), .B(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT80), .B(KEYINPUT23), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G183gat), .A2(G190gat), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n268_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(G183gat), .A2(G190gat), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n276_));
  INV_X1    g075(.A(G169gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n275_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(G183gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT25), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT25), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(G183gat), .ZN(new_n284_));
  INV_X1    g083(.A(G190gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT26), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT26), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(G190gat), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n282_), .A2(new_n284_), .A3(new_n286_), .A4(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT78), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT25), .B(G183gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT78), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n291_), .A2(new_n292_), .A3(new_n286_), .A4(new_n288_), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n290_), .A2(new_n293_), .ZN(new_n294_));
  AND2_X1   g093(.A1(KEYINPUT80), .A2(KEYINPUT23), .ZN(new_n295_));
  NOR2_X1   g094(.A1(KEYINPUT80), .A2(KEYINPUT23), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n270_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT23), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n271_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT24), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT79), .ZN(new_n302_));
  NOR3_X1   g101(.A1(new_n302_), .A2(G169gat), .A3(G176gat), .ZN(new_n303_));
  INV_X1    g102(.A(G176gat), .ZN(new_n304_));
  AOI21_X1  g103(.A(KEYINPUT79), .B1(new_n277_), .B2(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n301_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n277_), .A2(new_n304_), .A3(KEYINPUT79), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n302_), .B1(G169gat), .B2(G176gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n307_), .A2(new_n308_), .A3(KEYINPUT24), .A4(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n300_), .A2(new_n306_), .A3(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n280_), .B1(new_n294_), .B2(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n259_), .B1(new_n267_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n266_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n263_), .B(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n278_), .B1(new_n272_), .B2(new_n274_), .ZN(new_n316_));
  AND3_X1   g115(.A1(new_n300_), .A2(new_n306_), .A3(new_n310_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n290_), .A2(new_n293_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n316_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n315_), .A2(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT31), .B1(new_n313_), .B2(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(G127gat), .B(G134gat), .Z(new_n322_));
  XOR2_X1   g121(.A(G113gat), .B(G120gat), .Z(new_n323_));
  XOR2_X1   g122(.A(new_n322_), .B(new_n323_), .Z(new_n324_));
  AOI21_X1  g123(.A(KEYINPUT81), .B1(new_n315_), .B2(new_n319_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT31), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n267_), .A2(new_n312_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n325_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n321_), .A2(new_n324_), .A3(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n324_), .B1(new_n321_), .B2(new_n328_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(G228gat), .ZN(new_n333_));
  INV_X1    g132(.A(G233gat), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT29), .ZN(new_n336_));
  NOR2_X1   g135(.A1(G155gat), .A2(G162gat), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G155gat), .A2(G162gat), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n338_), .A2(KEYINPUT87), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT87), .ZN(new_n341_));
  AND2_X1   g140(.A1(G155gat), .A2(G162gat), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n341_), .B1(new_n342_), .B2(new_n337_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n340_), .A2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT86), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT86), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n347_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT3), .ZN(new_n349_));
  INV_X1    g148(.A(G141gat), .ZN(new_n350_));
  INV_X1    g149(.A(G148gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n349_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n346_), .A2(new_n348_), .A3(new_n352_), .A4(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(KEYINPUT82), .A2(G141gat), .A3(G148gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT82), .B1(G141gat), .B2(G148gat), .ZN(new_n357_));
  NOR3_X1   g156(.A1(new_n356_), .A2(new_n357_), .A3(KEYINPUT2), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n344_), .B1(new_n354_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT88), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n344_), .B(KEYINPUT88), .C1(new_n354_), .C2(new_n358_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT84), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n364_), .B1(new_n339_), .B2(KEYINPUT1), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT1), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n366_), .A2(KEYINPUT84), .A3(G155gat), .A4(G162gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n339_), .A2(KEYINPUT1), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n365_), .A2(new_n367_), .A3(new_n368_), .A4(new_n338_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n356_), .A2(new_n357_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n350_), .A2(new_n351_), .A3(KEYINPUT83), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT83), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n372_), .B1(G141gat), .B2(G148gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n369_), .A2(new_n370_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT85), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT85), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n369_), .A2(new_n377_), .A3(new_n370_), .A4(new_n374_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n336_), .B1(new_n363_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(G218gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(G211gat), .ZN(new_n382_));
  INV_X1    g181(.A(G211gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(G218gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT21), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G197gat), .B(G204gat), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n385_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(G197gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(G204gat), .ZN(new_n390_));
  INV_X1    g189(.A(G204gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(G197gat), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n390_), .A2(new_n392_), .A3(KEYINPUT90), .ZN(new_n393_));
  OR3_X1    g192(.A1(new_n391_), .A2(KEYINPUT90), .A3(G197gat), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n393_), .A2(new_n394_), .A3(KEYINPUT21), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n388_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n385_), .A2(KEYINPUT91), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n390_), .A2(new_n392_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT91), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n382_), .A2(new_n384_), .A3(new_n399_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n397_), .A2(KEYINPUT21), .A3(new_n398_), .A4(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n396_), .A2(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n402_), .A2(KEYINPUT92), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT92), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n404_), .B1(new_n396_), .B2(new_n401_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n335_), .B1(new_n380_), .B2(new_n406_), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n361_), .A2(new_n362_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n408_));
  OAI221_X1 g207(.A(new_n402_), .B1(new_n333_), .B2(new_n334_), .C1(new_n408_), .C2(new_n336_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G78gat), .B(G106gat), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT94), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n407_), .A2(new_n409_), .A3(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n412_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n352_), .A2(new_n353_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n357_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT2), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n417_), .A2(new_n418_), .A3(new_n355_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n416_), .A2(new_n419_), .A3(new_n348_), .A4(new_n346_), .ZN(new_n420_));
  AOI21_X1  g219(.A(KEYINPUT88), .B1(new_n420_), .B2(new_n344_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n362_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n379_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT28), .B1(new_n423_), .B2(KEYINPUT29), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT89), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT28), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n408_), .A2(new_n426_), .A3(new_n336_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n424_), .A2(new_n425_), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n425_), .B1(new_n424_), .B2(new_n427_), .ZN(new_n430_));
  XOR2_X1   g229(.A(G22gat), .B(G50gat), .Z(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NOR3_X1   g231(.A1(new_n429_), .A2(new_n430_), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n427_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n426_), .B1(new_n408_), .B2(new_n336_), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT89), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n431_), .B1(new_n436_), .B2(new_n428_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n415_), .B1(new_n433_), .B2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n432_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n407_), .A2(new_n409_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n410_), .A2(KEYINPUT93), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n436_), .A2(new_n431_), .A3(new_n428_), .ZN(new_n443_));
  XOR2_X1   g242(.A(new_n410_), .B(KEYINPUT93), .Z(new_n444_));
  NAND3_X1  g243(.A1(new_n407_), .A2(new_n409_), .A3(new_n444_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n439_), .A2(new_n442_), .A3(new_n443_), .A4(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n438_), .A2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G1gat), .B(G29gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(G85gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT0), .B(G57gat), .ZN(new_n450_));
  XOR2_X1   g249(.A(new_n449_), .B(new_n450_), .Z(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G225gat), .A2(G233gat), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT4), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n324_), .A2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n454_), .B1(new_n408_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT100), .ZN(new_n458_));
  INV_X1    g257(.A(new_n324_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n423_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n458_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n324_), .A2(KEYINPUT100), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n408_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n460_), .A2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n457_), .B1(new_n464_), .B2(KEYINPUT4), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n454_), .B1(new_n460_), .B2(new_n463_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n452_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT102), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n464_), .A2(new_n453_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n455_), .B1(new_n460_), .B2(new_n463_), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n469_), .B(new_n451_), .C1(new_n470_), .C2(new_n457_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n467_), .A2(new_n468_), .A3(new_n471_), .ZN(new_n472_));
  OAI211_X1 g271(.A(KEYINPUT102), .B(new_n452_), .C1(new_n465_), .C2(new_n466_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n447_), .A2(new_n474_), .ZN(new_n475_));
  XOR2_X1   g274(.A(G8gat), .B(G36gat), .Z(new_n476_));
  XNOR2_X1  g275(.A(G64gat), .B(G92gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G226gat), .A2(G233gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT19), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT97), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n400_), .A2(KEYINPUT21), .A3(new_n398_), .ZN(new_n484_));
  AOI22_X1  g283(.A1(new_n484_), .A2(new_n397_), .B1(new_n388_), .B2(new_n395_), .ZN(new_n485_));
  NOR3_X1   g284(.A1(new_n319_), .A2(new_n483_), .A3(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(KEYINPUT97), .B1(new_n312_), .B2(new_n402_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT96), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT22), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n490_), .A2(G169gat), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n277_), .A2(KEYINPUT22), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n489_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n277_), .A2(KEYINPUT22), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n490_), .A2(G169gat), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n494_), .A2(new_n495_), .A3(KEYINPUT96), .ZN(new_n496_));
  AOI21_X1  g295(.A(G176gat), .B1(new_n493_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n309_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n273_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n499_));
  NOR3_X1   g298(.A1(new_n497_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n286_), .A2(new_n288_), .A3(KEYINPUT95), .ZN(new_n501_));
  AOI21_X1  g300(.A(KEYINPUT95), .B1(new_n286_), .B2(new_n288_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n282_), .A2(new_n284_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n501_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n271_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n268_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n301_), .A2(new_n277_), .A3(new_n304_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n310_), .A2(new_n505_), .A3(new_n506_), .A4(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n504_), .A2(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n500_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n405_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n485_), .A2(new_n404_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT20), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n482_), .B1(new_n488_), .B2(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n402_), .B1(new_n500_), .B2(new_n509_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n303_), .A2(new_n305_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n498_), .A2(new_n301_), .ZN(new_n518_));
  AOI22_X1  g317(.A1(new_n517_), .A2(new_n518_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n318_), .A2(new_n519_), .A3(new_n306_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n520_), .A2(new_n485_), .A3(new_n280_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n516_), .A2(KEYINPUT20), .A3(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n522_), .A2(new_n482_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n480_), .B1(new_n515_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n522_), .A2(new_n482_), .ZN(new_n526_));
  AND3_X1   g325(.A1(new_n494_), .A2(new_n495_), .A3(KEYINPUT96), .ZN(new_n527_));
  AOI21_X1  g326(.A(KEYINPUT96), .B1(new_n494_), .B2(new_n495_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n304_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n300_), .A2(new_n274_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(new_n530_), .A3(new_n309_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT95), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n287_), .A2(G190gat), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n285_), .A2(KEYINPUT26), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n532_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n286_), .A2(new_n288_), .A3(KEYINPUT95), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n535_), .A2(new_n291_), .A3(new_n536_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n537_), .A2(new_n310_), .A3(new_n272_), .A4(new_n507_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n485_), .A2(new_n531_), .A3(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT98), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT98), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n485_), .A2(new_n531_), .A3(new_n538_), .A4(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT20), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n482_), .A2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n540_), .A2(new_n542_), .A3(new_n544_), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n526_), .B(new_n480_), .C1(new_n488_), .C2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT27), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n525_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT103), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n526_), .B1(new_n488_), .B2(new_n545_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n480_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(new_n546_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT27), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n550_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  AOI211_X1 g355(.A(KEYINPUT103), .B(KEYINPUT27), .C1(new_n553_), .C2(new_n546_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n549_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n475_), .A2(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n483_), .B1(new_n319_), .B2(new_n485_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n312_), .A2(KEYINPUT97), .A3(new_n402_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n562_), .A2(KEYINPUT20), .A3(new_n513_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n523_), .B1(new_n563_), .B2(new_n482_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n480_), .A2(KEYINPUT32), .ZN(new_n565_));
  OAI21_X1  g364(.A(KEYINPUT101), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT101), .ZN(new_n567_));
  INV_X1    g366(.A(new_n565_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n482_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n543_), .B1(new_n406_), .B2(new_n510_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n569_), .B1(new_n570_), .B2(new_n562_), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n567_), .B(new_n568_), .C1(new_n571_), .C2(new_n523_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n566_), .A2(new_n572_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n542_), .A2(new_n544_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n562_), .A2(new_n540_), .A3(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n575_), .A2(new_n526_), .A3(new_n565_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n573_), .A2(new_n472_), .A3(new_n473_), .A4(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n465_), .A2(new_n466_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n578_), .A2(KEYINPUT33), .A3(new_n451_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n554_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT33), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n471_), .A2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n451_), .B1(new_n464_), .B2(new_n454_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n453_), .B1(new_n408_), .B2(new_n456_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n583_), .B1(new_n470_), .B2(new_n584_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n579_), .A2(new_n580_), .A3(new_n582_), .A4(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n447_), .B1(new_n577_), .B2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n332_), .B1(new_n559_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n447_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n331_), .A2(new_n474_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n546_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n480_), .B1(new_n575_), .B2(new_n526_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n555_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT103), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n554_), .A2(new_n550_), .A3(new_n555_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(KEYINPUT104), .B1(new_n596_), .B2(new_n549_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT104), .ZN(new_n598_));
  AOI211_X1 g397(.A(new_n598_), .B(new_n548_), .C1(new_n594_), .C2(new_n595_), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n589_), .B(new_n590_), .C1(new_n597_), .C2(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n258_), .B1(new_n588_), .B2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G230gat), .A2(G233gat), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G99gat), .A2(G106gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT6), .ZN(new_n604_));
  OAI21_X1  g403(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT7), .ZN(new_n606_));
  INV_X1    g405(.A(G99gat), .ZN(new_n607_));
  INV_X1    g406(.A(G106gat), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n606_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n604_), .A2(new_n605_), .A3(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT8), .ZN(new_n611_));
  INV_X1    g410(.A(G85gat), .ZN(new_n612_));
  INV_X1    g411(.A(G92gat), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G85gat), .A2(G92gat), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n610_), .A2(new_n611_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT6), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n603_), .B(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n609_), .A2(new_n605_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n616_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT8), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n617_), .A2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G57gat), .B(G64gat), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(KEYINPUT11), .ZN(new_n625_));
  XOR2_X1   g424(.A(G71gat), .B(G78gat), .Z(new_n626_));
  OR2_X1    g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n624_), .A2(KEYINPUT11), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n625_), .A2(new_n626_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n627_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT9), .ZN(new_n631_));
  AOI21_X1  g430(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT64), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n632_), .A2(new_n633_), .ZN(new_n635_));
  OAI221_X1 g434(.A(new_n614_), .B1(new_n631_), .B2(new_n615_), .C1(new_n634_), .C2(new_n635_), .ZN(new_n636_));
  XOR2_X1   g435(.A(KEYINPUT10), .B(G99gat), .Z(new_n637_));
  AOI21_X1  g436(.A(new_n619_), .B1(new_n608_), .B2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n623_), .A2(new_n630_), .A3(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(KEYINPUT12), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n630_), .B1(new_n623_), .B2(new_n639_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n611_), .B1(new_n610_), .B2(new_n616_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n621_), .A2(KEYINPUT8), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n639_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n630_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT12), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n646_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n602_), .B1(new_n643_), .B2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(KEYINPUT67), .ZN(new_n652_));
  INV_X1    g451(.A(new_n602_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n646_), .A2(new_n647_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n654_), .A2(KEYINPUT12), .A3(new_n640_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n653_), .B1(new_n655_), .B2(new_n649_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT67), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n640_), .A2(KEYINPUT65), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT66), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n654_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n642_), .A2(KEYINPUT66), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n640_), .A2(KEYINPUT65), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n659_), .A2(new_n661_), .A3(new_n662_), .A4(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(new_n653_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n652_), .A2(new_n658_), .A3(new_n665_), .ZN(new_n666_));
  XOR2_X1   g465(.A(KEYINPUT68), .B(KEYINPUT5), .Z(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT69), .ZN(new_n668_));
  XNOR2_X1  g467(.A(G120gat), .B(G148gat), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n668_), .B(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(G176gat), .B(G204gat), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n670_), .B(new_n671_), .Z(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n666_), .A2(new_n673_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n652_), .A2(new_n665_), .A3(new_n658_), .A4(new_n672_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT13), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n674_), .A2(KEYINPUT13), .A3(new_n675_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(G231gat), .A2(G233gat), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n630_), .B(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n216_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n683_), .B(new_n684_), .ZN(new_n685_));
  XOR2_X1   g484(.A(G127gat), .B(G155gat), .Z(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT16), .ZN(new_n687_));
  XNOR2_X1  g486(.A(G183gat), .B(G211gat), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT17), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n685_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT74), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n692_), .B(new_n693_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n689_), .A2(new_n690_), .ZN(new_n695_));
  OR3_X1    g494(.A1(new_n685_), .A2(new_n691_), .A3(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(G190gat), .B(G218gat), .ZN(new_n698_));
  XNOR2_X1  g497(.A(G134gat), .B(G162gat), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n698_), .B(new_n699_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT36), .Z(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n623_), .A2(new_n225_), .A3(new_n639_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(G232gat), .A2(G233gat), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT34), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT35), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n703_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n227_), .A2(new_n224_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n710_), .B1(new_n623_), .B2(new_n639_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n706_), .A2(new_n707_), .ZN(new_n712_));
  OR3_X1    g511(.A1(new_n709_), .A2(new_n711_), .A3(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n712_), .B1(new_n709_), .B2(new_n711_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n702_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n700_), .A2(KEYINPUT36), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n713_), .A2(new_n717_), .A3(new_n714_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n716_), .B1(KEYINPUT71), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n718_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT71), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(KEYINPUT37), .B1(new_n719_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n716_), .A2(KEYINPUT72), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT72), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n715_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT37), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n724_), .A2(new_n726_), .A3(new_n727_), .A4(new_n718_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n697_), .B1(new_n723_), .B2(new_n728_), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n601_), .A2(new_n681_), .A3(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n474_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n203_), .A3(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT38), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n697_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n724_), .A2(new_n718_), .A3(new_n726_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n588_), .B2(new_n600_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT105), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n739_), .B1(new_n680_), .B2(new_n258_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n681_), .A2(KEYINPUT105), .A3(new_n257_), .ZN(new_n741_));
  AND4_X1   g540(.A1(new_n735_), .A2(new_n738_), .A3(new_n740_), .A4(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n203_), .B1(new_n742_), .B2(new_n731_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n734_), .A2(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n744_), .B1(new_n733_), .B2(new_n732_), .ZN(G1324gat));
  NOR2_X1   g544(.A1(new_n597_), .A2(new_n599_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n730_), .A2(new_n204_), .A3(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT39), .ZN(new_n748_));
  OAI21_X1  g547(.A(G8gat), .B1(new_n748_), .B2(KEYINPUT106), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n742_), .B2(new_n746_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n750_), .A2(KEYINPUT106), .A3(new_n748_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(KEYINPUT106), .B2(new_n748_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n747_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT40), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n753_), .B(new_n754_), .ZN(G1325gat));
  AOI21_X1  g554(.A(new_n265_), .B1(new_n742_), .B2(new_n331_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT41), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n730_), .A2(new_n265_), .A3(new_n331_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1326gat));
  INV_X1    g558(.A(G22gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(new_n742_), .B2(new_n447_), .ZN(new_n761_));
  XOR2_X1   g560(.A(new_n761_), .B(KEYINPUT42), .Z(new_n762_));
  NAND3_X1  g561(.A1(new_n730_), .A2(new_n760_), .A3(new_n447_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1327gat));
  NOR3_X1   g563(.A1(new_n680_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n601_), .A2(new_n765_), .ZN(new_n766_));
  OR3_X1    g565(.A1(new_n766_), .A2(G29gat), .A3(new_n474_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n741_), .A2(new_n697_), .A3(new_n740_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT43), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n588_), .A2(new_n600_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n723_), .A2(new_n728_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n770_), .B1(new_n771_), .B2(new_n773_), .ZN(new_n774_));
  AOI211_X1 g573(.A(KEYINPUT43), .B(new_n772_), .C1(new_n588_), .C2(new_n600_), .ZN(new_n775_));
  OAI211_X1 g574(.A(KEYINPUT44), .B(new_n769_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n771_), .A2(new_n773_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT43), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n771_), .A2(new_n770_), .A3(new_n773_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n768_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(KEYINPUT107), .B1(new_n781_), .B2(KEYINPUT44), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n769_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT107), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT44), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n783_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n777_), .B1(new_n782_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT108), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n788_), .A3(new_n731_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(G29gat), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n788_), .B1(new_n787_), .B2(new_n731_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n767_), .B1(new_n790_), .B2(new_n791_), .ZN(G1328gat));
  XNOR2_X1  g591(.A(KEYINPUT111), .B(KEYINPUT46), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(G36gat), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n787_), .B2(new_n746_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT110), .ZN(new_n797_));
  INV_X1    g596(.A(new_n766_), .ZN(new_n798_));
  OR2_X1    g597(.A1(new_n746_), .A2(KEYINPUT109), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n746_), .A2(KEYINPUT109), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n801_), .A2(G36gat), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n797_), .B1(new_n798_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n798_), .A2(new_n802_), .A3(new_n797_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(KEYINPUT45), .A3(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT45), .ZN(new_n807_));
  INV_X1    g606(.A(new_n805_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n807_), .B1(new_n808_), .B2(new_n803_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n806_), .A2(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n794_), .B1(new_n796_), .B2(new_n810_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n806_), .A2(new_n809_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n746_), .ZN(new_n813_));
  AOI211_X1 g612(.A(new_n813_), .B(new_n777_), .C1(new_n782_), .C2(new_n786_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n812_), .B(new_n793_), .C1(new_n814_), .C2(new_n795_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n811_), .A2(new_n815_), .ZN(G1329gat));
  XNOR2_X1  g615(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n261_), .B1(new_n787_), .B2(new_n331_), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n766_), .A2(G43gat), .A3(new_n332_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n818_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n820_), .ZN(new_n822_));
  AOI211_X1 g621(.A(new_n332_), .B(new_n777_), .C1(new_n782_), .C2(new_n786_), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n822_), .B(new_n817_), .C1(new_n823_), .C2(new_n261_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n821_), .A2(new_n824_), .ZN(G1330gat));
  INV_X1    g624(.A(KEYINPUT113), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n783_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n784_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n447_), .B(new_n776_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(G50gat), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n589_), .A2(G50gat), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n798_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n826_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n832_), .ZN(new_n834_));
  AOI211_X1 g633(.A(KEYINPUT113), .B(new_n834_), .C1(new_n829_), .C2(G50gat), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n833_), .A2(new_n835_), .ZN(G1331gat));
  NOR2_X1   g635(.A1(new_n681_), .A2(new_n257_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n771_), .A2(new_n837_), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n838_), .A2(new_n697_), .A3(new_n773_), .ZN(new_n839_));
  INV_X1    g638(.A(G57gat), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n840_), .A3(new_n731_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n738_), .A2(new_n735_), .A3(new_n837_), .ZN(new_n842_));
  OR2_X1    g641(.A1(new_n842_), .A2(KEYINPUT114), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(KEYINPUT114), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n845_), .A2(new_n731_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n841_), .B1(new_n846_), .B2(new_n840_), .ZN(G1332gat));
  INV_X1    g646(.A(G64gat), .ZN(new_n848_));
  INV_X1    g647(.A(new_n801_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n839_), .A2(new_n848_), .A3(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n843_), .A2(new_n849_), .A3(new_n844_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(KEYINPUT115), .B(KEYINPUT48), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n851_), .A2(G64gat), .A3(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n851_), .B2(G64gat), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n850_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  OAI211_X1 g656(.A(KEYINPUT116), .B(new_n850_), .C1(new_n853_), .C2(new_n854_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(G1333gat));
  INV_X1    g658(.A(G71gat), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n839_), .A2(new_n860_), .A3(new_n331_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n845_), .A2(new_n331_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(G71gat), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n863_), .A2(KEYINPUT49), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n863_), .A2(KEYINPUT49), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n861_), .B1(new_n864_), .B2(new_n865_), .ZN(G1334gat));
  INV_X1    g665(.A(G78gat), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n839_), .A2(new_n867_), .A3(new_n447_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n845_), .A2(new_n447_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(G78gat), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n870_), .A2(KEYINPUT50), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n870_), .A2(KEYINPUT50), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n868_), .B1(new_n871_), .B2(new_n872_), .ZN(G1335gat));
  NOR3_X1   g672(.A1(new_n838_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n874_), .A2(new_n612_), .A3(new_n731_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n837_), .A2(new_n697_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(KEYINPUT117), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n779_), .A2(new_n780_), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n731_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n875_), .B1(new_n881_), .B2(new_n612_), .ZN(G1336gat));
  NAND3_X1  g681(.A1(new_n874_), .A2(new_n613_), .A3(new_n746_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n879_), .A2(new_n849_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n883_), .B1(new_n885_), .B2(new_n613_), .ZN(G1337gat));
  NAND3_X1  g685(.A1(new_n874_), .A2(new_n331_), .A3(new_n637_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n879_), .A2(new_n331_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n887_), .B1(new_n889_), .B2(new_n607_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g690(.A1(new_n874_), .A2(new_n608_), .A3(new_n447_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n877_), .A2(new_n878_), .A3(new_n447_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT52), .ZN(new_n894_));
  AND3_X1   g693(.A1(new_n893_), .A2(new_n894_), .A3(G106gat), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n894_), .B1(new_n893_), .B2(G106gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n892_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n729_), .A2(new_n258_), .A3(new_n678_), .A4(new_n679_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(KEYINPUT118), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n900_), .A2(KEYINPUT118), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n899_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n903_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n905_), .A2(KEYINPUT54), .A3(new_n901_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT56), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n655_), .A2(new_n653_), .A3(new_n649_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT55), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n909_), .B1(new_n651_), .B2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n655_), .A2(new_n649_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n657_), .B1(new_n912_), .B2(new_n602_), .ZN(new_n913_));
  AOI211_X1 g712(.A(KEYINPUT67), .B(new_n653_), .C1(new_n655_), .C2(new_n649_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n911_), .B1(new_n915_), .B2(new_n910_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n908_), .B1(new_n916_), .B2(new_n672_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n652_), .A2(new_n910_), .A3(new_n658_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n909_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n919_), .B1(KEYINPUT55), .B2(new_n656_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n918_), .A2(new_n920_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n921_), .A2(KEYINPUT56), .A3(new_n673_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n917_), .A2(KEYINPUT119), .A3(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n257_), .A2(new_n675_), .ZN(new_n924_));
  AOI211_X1 g723(.A(new_n908_), .B(new_n672_), .C1(new_n918_), .C2(new_n920_), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT119), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n924_), .B1(new_n925_), .B2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n923_), .A2(new_n927_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n237_), .A2(new_n240_), .A3(new_n232_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT120), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n253_), .B1(new_n247_), .B2(new_n230_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n929_), .A2(new_n930_), .A3(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n929_), .A2(new_n931_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(KEYINPUT120), .ZN(new_n934_));
  AND3_X1   g733(.A1(new_n256_), .A2(new_n932_), .A3(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n676_), .A2(new_n935_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n928_), .A2(new_n936_), .ZN(new_n937_));
  AOI21_X1  g736(.A(KEYINPUT57), .B1(new_n937_), .B2(new_n736_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n936_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n939_), .B1(new_n923_), .B2(new_n927_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT57), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n940_), .A2(new_n941_), .A3(new_n737_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n938_), .A2(new_n942_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT58), .ZN(new_n944_));
  AND4_X1   g743(.A1(new_n652_), .A2(new_n658_), .A3(new_n665_), .A4(new_n672_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n256_), .A2(new_n934_), .A3(new_n932_), .ZN(new_n946_));
  OAI21_X1  g745(.A(KEYINPUT121), .B1(new_n945_), .B2(new_n946_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT121), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n935_), .A2(new_n948_), .A3(new_n675_), .ZN(new_n949_));
  AOI22_X1  g748(.A1(new_n917_), .A2(new_n922_), .B1(new_n947_), .B2(new_n949_), .ZN(new_n950_));
  INV_X1    g749(.A(KEYINPUT122), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n944_), .B1(new_n950_), .B2(new_n951_), .ZN(new_n952_));
  AOI21_X1  g751(.A(KEYINPUT56), .B1(new_n921_), .B2(new_n673_), .ZN(new_n953_));
  AND3_X1   g752(.A1(new_n935_), .A2(new_n948_), .A3(new_n675_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n948_), .B1(new_n935_), .B2(new_n675_), .ZN(new_n955_));
  OAI22_X1  g754(.A1(new_n953_), .A2(new_n925_), .B1(new_n954_), .B2(new_n955_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n956_), .A2(KEYINPUT122), .ZN(new_n957_));
  OAI211_X1 g756(.A(KEYINPUT123), .B(new_n773_), .C1(new_n952_), .C2(new_n957_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n950_), .A2(KEYINPUT58), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n958_), .A2(new_n959_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n950_), .A2(new_n951_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n956_), .A2(KEYINPUT122), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n961_), .A2(new_n962_), .A3(new_n944_), .ZN(new_n963_));
  AOI21_X1  g762(.A(KEYINPUT123), .B1(new_n963_), .B2(new_n773_), .ZN(new_n964_));
  OAI21_X1  g763(.A(new_n943_), .B1(new_n960_), .B2(new_n964_), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n907_), .B1(new_n965_), .B2(new_n697_), .ZN(new_n966_));
  NOR2_X1   g765(.A1(new_n746_), .A2(new_n447_), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n967_), .A2(new_n731_), .A3(new_n331_), .ZN(new_n968_));
  NOR2_X1   g767(.A1(new_n966_), .A2(new_n968_), .ZN(new_n969_));
  INV_X1    g768(.A(G113gat), .ZN(new_n970_));
  NAND3_X1  g769(.A1(new_n969_), .A2(new_n970_), .A3(new_n257_), .ZN(new_n971_));
  INV_X1    g770(.A(new_n968_), .ZN(new_n972_));
  OAI21_X1  g771(.A(new_n773_), .B1(new_n952_), .B2(new_n957_), .ZN(new_n973_));
  INV_X1    g772(.A(KEYINPUT123), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n973_), .A2(new_n974_), .ZN(new_n975_));
  NAND3_X1  g774(.A1(new_n975_), .A2(new_n959_), .A3(new_n958_), .ZN(new_n976_));
  AOI21_X1  g775(.A(new_n735_), .B1(new_n976_), .B2(new_n943_), .ZN(new_n977_));
  OAI211_X1 g776(.A(KEYINPUT124), .B(new_n972_), .C1(new_n977_), .C2(new_n907_), .ZN(new_n978_));
  INV_X1    g777(.A(KEYINPUT59), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n978_), .A2(new_n979_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n965_), .A2(new_n697_), .ZN(new_n981_));
  INV_X1    g780(.A(new_n907_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n981_), .A2(new_n982_), .ZN(new_n983_));
  NAND4_X1  g782(.A1(new_n983_), .A2(KEYINPUT124), .A3(KEYINPUT59), .A4(new_n972_), .ZN(new_n984_));
  AOI21_X1  g783(.A(new_n258_), .B1(new_n980_), .B2(new_n984_), .ZN(new_n985_));
  OAI21_X1  g784(.A(new_n971_), .B1(new_n985_), .B2(new_n970_), .ZN(G1340gat));
  INV_X1    g785(.A(G120gat), .ZN(new_n987_));
  OAI21_X1  g786(.A(new_n987_), .B1(new_n681_), .B2(KEYINPUT60), .ZN(new_n988_));
  OAI211_X1 g787(.A(new_n969_), .B(new_n988_), .C1(KEYINPUT60), .C2(new_n987_), .ZN(new_n989_));
  AOI21_X1  g788(.A(new_n681_), .B1(new_n980_), .B2(new_n984_), .ZN(new_n990_));
  OAI21_X1  g789(.A(new_n989_), .B1(new_n990_), .B2(new_n987_), .ZN(G1341gat));
  INV_X1    g790(.A(G127gat), .ZN(new_n992_));
  NAND3_X1  g791(.A1(new_n969_), .A2(new_n992_), .A3(new_n735_), .ZN(new_n993_));
  AOI21_X1  g792(.A(new_n697_), .B1(new_n980_), .B2(new_n984_), .ZN(new_n994_));
  OAI21_X1  g793(.A(new_n993_), .B1(new_n994_), .B2(new_n992_), .ZN(G1342gat));
  NAND2_X1  g794(.A1(new_n773_), .A2(G134gat), .ZN(new_n996_));
  AOI21_X1  g795(.A(new_n996_), .B1(new_n980_), .B2(new_n984_), .ZN(new_n997_));
  NOR3_X1   g796(.A1(new_n966_), .A2(new_n736_), .A3(new_n968_), .ZN(new_n998_));
  NOR3_X1   g797(.A1(new_n998_), .A2(KEYINPUT125), .A3(G134gat), .ZN(new_n999_));
  INV_X1    g798(.A(KEYINPUT125), .ZN(new_n1000_));
  NAND3_X1  g799(.A1(new_n983_), .A2(new_n737_), .A3(new_n972_), .ZN(new_n1001_));
  INV_X1    g800(.A(G134gat), .ZN(new_n1002_));
  AOI21_X1  g801(.A(new_n1000_), .B1(new_n1001_), .B2(new_n1002_), .ZN(new_n1003_));
  NOR3_X1   g802(.A1(new_n997_), .A2(new_n999_), .A3(new_n1003_), .ZN(G1343gat));
  NOR2_X1   g803(.A1(new_n966_), .A2(new_n331_), .ZN(new_n1005_));
  NOR3_X1   g804(.A1(new_n849_), .A2(new_n474_), .A3(new_n589_), .ZN(new_n1006_));
  NAND3_X1  g805(.A1(new_n1005_), .A2(new_n257_), .A3(new_n1006_), .ZN(new_n1007_));
  XNOR2_X1  g806(.A(new_n1007_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g807(.A1(new_n1005_), .A2(new_n680_), .A3(new_n1006_), .ZN(new_n1009_));
  XNOR2_X1  g808(.A(new_n1009_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g809(.A1(new_n1005_), .A2(new_n735_), .A3(new_n1006_), .ZN(new_n1011_));
  XNOR2_X1  g810(.A(KEYINPUT61), .B(G155gat), .ZN(new_n1012_));
  XNOR2_X1  g811(.A(new_n1011_), .B(new_n1012_), .ZN(G1346gat));
  AND4_X1   g812(.A1(G162gat), .A2(new_n1005_), .A3(new_n773_), .A4(new_n1006_), .ZN(new_n1014_));
  NAND4_X1  g813(.A1(new_n983_), .A2(new_n332_), .A3(new_n737_), .A4(new_n1006_), .ZN(new_n1015_));
  INV_X1    g814(.A(G162gat), .ZN(new_n1016_));
  NAND2_X1  g815(.A1(new_n1015_), .A2(new_n1016_), .ZN(new_n1017_));
  INV_X1    g816(.A(KEYINPUT126), .ZN(new_n1018_));
  NAND2_X1  g817(.A1(new_n1017_), .A2(new_n1018_), .ZN(new_n1019_));
  NAND3_X1  g818(.A1(new_n1015_), .A2(KEYINPUT126), .A3(new_n1016_), .ZN(new_n1020_));
  AOI21_X1  g819(.A(new_n1014_), .B1(new_n1019_), .B2(new_n1020_), .ZN(G1347gat));
  NOR4_X1   g820(.A1(new_n801_), .A2(new_n731_), .A3(new_n447_), .A4(new_n332_), .ZN(new_n1022_));
  NAND3_X1  g821(.A1(new_n983_), .A2(new_n257_), .A3(new_n1022_), .ZN(new_n1023_));
  INV_X1    g822(.A(KEYINPUT62), .ZN(new_n1024_));
  AND3_X1   g823(.A1(new_n1023_), .A2(new_n1024_), .A3(G169gat), .ZN(new_n1025_));
  AND2_X1   g824(.A1(new_n983_), .A2(new_n1022_), .ZN(new_n1026_));
  OAI211_X1 g825(.A(new_n1026_), .B(new_n257_), .C1(new_n527_), .C2(new_n528_), .ZN(new_n1027_));
  AOI21_X1  g826(.A(new_n1024_), .B1(new_n1023_), .B2(G169gat), .ZN(new_n1028_));
  AOI21_X1  g827(.A(new_n1025_), .B1(new_n1027_), .B2(new_n1028_), .ZN(G1348gat));
  AND3_X1   g828(.A1(new_n1026_), .A2(G176gat), .A3(new_n680_), .ZN(new_n1030_));
  AOI21_X1  g829(.A(G176gat), .B1(new_n1026_), .B2(new_n680_), .ZN(new_n1031_));
  NOR2_X1   g830(.A1(new_n1030_), .A2(new_n1031_), .ZN(G1349gat));
  AOI21_X1  g831(.A(G183gat), .B1(new_n1026_), .B2(new_n735_), .ZN(new_n1033_));
  AND2_X1   g832(.A1(new_n1026_), .A2(new_n735_), .ZN(new_n1034_));
  AOI21_X1  g833(.A(new_n1033_), .B1(new_n503_), .B2(new_n1034_), .ZN(G1350gat));
  NAND4_X1  g834(.A1(new_n1026_), .A2(new_n535_), .A3(new_n536_), .A4(new_n737_), .ZN(new_n1036_));
  AND2_X1   g835(.A1(new_n1026_), .A2(new_n773_), .ZN(new_n1037_));
  OAI21_X1  g836(.A(new_n1036_), .B1(new_n1037_), .B2(new_n285_), .ZN(G1351gat));
  NOR2_X1   g837(.A1(new_n801_), .A2(new_n475_), .ZN(new_n1039_));
  NAND3_X1  g838(.A1(new_n1005_), .A2(new_n257_), .A3(new_n1039_), .ZN(new_n1040_));
  XNOR2_X1  g839(.A(new_n1040_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g840(.A1(new_n1005_), .A2(new_n680_), .A3(new_n1039_), .ZN(new_n1042_));
  XNOR2_X1  g841(.A(new_n1042_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g842(.A1(new_n1005_), .A2(new_n735_), .A3(new_n1039_), .ZN(new_n1044_));
  XNOR2_X1  g843(.A(KEYINPUT63), .B(G211gat), .ZN(new_n1045_));
  NOR2_X1   g844(.A1(new_n1044_), .A2(new_n1045_), .ZN(new_n1046_));
  NOR2_X1   g845(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1047_));
  AOI21_X1  g846(.A(new_n1046_), .B1(new_n1044_), .B2(new_n1047_), .ZN(G1354gat));
  AND4_X1   g847(.A1(G218gat), .A2(new_n1005_), .A3(new_n773_), .A4(new_n1039_), .ZN(new_n1049_));
  INV_X1    g848(.A(new_n1039_), .ZN(new_n1050_));
  NOR4_X1   g849(.A1(new_n966_), .A2(new_n331_), .A3(new_n736_), .A4(new_n1050_), .ZN(new_n1051_));
  INV_X1    g850(.A(KEYINPUT127), .ZN(new_n1052_));
  OR2_X1    g851(.A1(new_n1051_), .A2(new_n1052_), .ZN(new_n1053_));
  AOI21_X1  g852(.A(G218gat), .B1(new_n1051_), .B2(new_n1052_), .ZN(new_n1054_));
  AOI21_X1  g853(.A(new_n1049_), .B1(new_n1053_), .B2(new_n1054_), .ZN(G1355gat));
endmodule


