//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 0 0 0 0 0 0 0 1 0 1 0 0 1 0 0 1 1 0 0 0 1 0 0 1 0 0 0 1 0 1 0 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n856_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n893_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_;
  XNOR2_X1  g000(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G232gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G29gat), .B(G36gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G43gat), .B(G50gat), .ZN(new_n207_));
  XOR2_X1   g006(.A(new_n206_), .B(new_n207_), .Z(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n206_), .B(new_n207_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n209_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT15), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n210_), .A2(KEYINPUT15), .A3(new_n213_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT6), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT6), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(G99gat), .A3(G106gat), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT7), .ZN(new_n224_));
  INV_X1    g023(.A(G99gat), .ZN(new_n225_));
  INV_X1    g024(.A(G106gat), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .A4(KEYINPUT64), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n228_));
  OAI22_X1  g027(.A1(new_n228_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n227_), .A2(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT65), .B1(new_n223_), .B2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n220_), .A2(new_n222_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n232_), .A2(new_n233_), .A3(new_n229_), .A4(new_n227_), .ZN(new_n234_));
  INV_X1    g033(.A(G85gat), .ZN(new_n235_));
  INV_X1    g034(.A(G92gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G85gat), .A2(G92gat), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT8), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n239_), .A2(KEYINPUT66), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(KEYINPUT66), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n237_), .B(new_n238_), .C1(new_n240_), .C2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n231_), .A2(new_n234_), .A3(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n237_), .A2(new_n238_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n246_), .B1(new_n223_), .B2(new_n230_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT8), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n244_), .A2(new_n248_), .ZN(new_n249_));
  OR2_X1    g048(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(new_n226_), .A3(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n237_), .A2(KEYINPUT9), .A3(new_n238_), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n238_), .A2(KEYINPUT9), .ZN(new_n254_));
  AND4_X1   g053(.A1(new_n232_), .A2(new_n252_), .A3(new_n253_), .A4(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT69), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n218_), .B1(new_n249_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n232_), .A2(new_n229_), .A3(new_n227_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n242_), .B1(new_n259_), .B2(KEYINPUT65), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n260_), .A2(new_n234_), .B1(KEYINPUT8), .B2(new_n247_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n258_), .B1(new_n261_), .B2(new_n255_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n255_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n249_), .A2(KEYINPUT67), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(new_n214_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  OAI211_X1 g066(.A(KEYINPUT35), .B(new_n205_), .C1(new_n257_), .C2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n218_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n256_), .A2(new_n249_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT35), .ZN(new_n271_));
  AOI22_X1  g070(.A1(new_n269_), .A2(new_n270_), .B1(new_n271_), .B2(new_n204_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n204_), .A2(new_n271_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n272_), .A2(new_n266_), .A3(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G190gat), .B(G218gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT73), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G134gat), .B(G162gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT36), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n281_), .B(KEYINPUT74), .Z(new_n282_));
  NAND3_X1  g081(.A1(new_n268_), .A2(new_n275_), .A3(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n279_), .B(new_n280_), .ZN(new_n285_));
  XOR2_X1   g084(.A(new_n285_), .B(KEYINPUT75), .Z(new_n286_));
  AOI21_X1  g085(.A(new_n286_), .B1(new_n275_), .B2(new_n268_), .ZN(new_n287_));
  OAI21_X1  g086(.A(KEYINPUT37), .B1(new_n284_), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n268_), .A2(new_n275_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n285_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT37), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(new_n292_), .A3(new_n283_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n288_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G15gat), .B(G22gat), .ZN(new_n295_));
  INV_X1    g094(.A(G1gat), .ZN(new_n296_));
  INV_X1    g095(.A(G8gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT14), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n295_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G1gat), .B(G8gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G231gat), .A2(G233gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G57gat), .B(G64gat), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n304_), .A2(KEYINPUT11), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(KEYINPUT11), .ZN(new_n306_));
  XOR2_X1   g105(.A(G71gat), .B(G78gat), .Z(new_n307_));
  NAND3_X1  g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n306_), .A2(new_n307_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n303_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n303_), .A2(new_n311_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G127gat), .B(G155gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT16), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G183gat), .B(G211gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XOR2_X1   g118(.A(new_n319_), .B(KEYINPUT17), .Z(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT78), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT76), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n314_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n312_), .A2(KEYINPUT76), .A3(new_n313_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n319_), .A2(KEYINPUT17), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT77), .ZN(new_n327_));
  AOI22_X1  g126(.A1(new_n315_), .A2(new_n321_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n294_), .A2(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n329_), .B(KEYINPUT79), .Z(new_n330_));
  AOI21_X1  g129(.A(KEYINPUT67), .B1(new_n249_), .B2(new_n263_), .ZN(new_n331_));
  AOI211_X1 g130(.A(new_n258_), .B(new_n255_), .C1(new_n244_), .C2(new_n248_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n310_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n262_), .A2(new_n264_), .A3(new_n311_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G230gat), .A2(G233gat), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT68), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT12), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n334_), .A2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n270_), .A2(KEYINPUT12), .A3(new_n311_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n341_), .A2(new_n336_), .A3(new_n333_), .A4(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT68), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n335_), .A2(new_n344_), .A3(new_n337_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n339_), .A2(new_n343_), .A3(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G120gat), .B(G148gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT5), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G176gat), .B(G204gat), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n348_), .B(new_n349_), .Z(new_n350_));
  NAND2_X1  g149(.A1(new_n346_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n350_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n339_), .A2(new_n343_), .A3(new_n345_), .A4(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT13), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n351_), .A2(KEYINPUT13), .A3(new_n353_), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n216_), .A2(new_n217_), .A3(new_n301_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n301_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n214_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G229gat), .A2(G233gat), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n359_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n210_), .A2(new_n213_), .A3(new_n301_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n361_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n362_), .ZN(new_n366_));
  AOI21_X1  g165(.A(KEYINPUT80), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT80), .ZN(new_n368_));
  AOI211_X1 g167(.A(new_n368_), .B(new_n362_), .C1(new_n361_), .C2(new_n364_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n363_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G113gat), .B(G141gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G169gat), .B(G197gat), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n371_), .B(new_n372_), .Z(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n370_), .A2(new_n374_), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n363_), .B(new_n373_), .C1(new_n367_), .C2(new_n369_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT20), .ZN(new_n379_));
  NOR2_X1   g178(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n380_), .B(G169gat), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G183gat), .A2(G190gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT23), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n384_), .B1(G183gat), .B2(G190gat), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n382_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n387_), .B1(new_n386_), .B2(new_n385_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT25), .B(G183gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT26), .B(G190gat), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT24), .ZN(new_n391_));
  NOR2_X1   g190(.A1(G169gat), .A2(G176gat), .ZN(new_n392_));
  AOI22_X1  g191(.A1(new_n389_), .A2(new_n390_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n391_), .B1(G169gat), .B2(G176gat), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n393_), .B(new_n384_), .C1(new_n392_), .C2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n388_), .A2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT88), .B(G197gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(G204gat), .ZN(new_n399_));
  INV_X1    g198(.A(G204gat), .ZN(new_n400_));
  AOI21_X1  g199(.A(KEYINPUT89), .B1(new_n400_), .B2(G197gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n398_), .A2(KEYINPUT89), .A3(G204gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G211gat), .B(G218gat), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT21), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n402_), .A2(new_n403_), .A3(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(KEYINPUT21), .B1(new_n402_), .B2(new_n403_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n398_), .A2(new_n400_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n405_), .B1(G197gat), .B2(G204gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(new_n404_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n407_), .B1(new_n408_), .B2(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n379_), .B1(new_n397_), .B2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G226gat), .A2(G233gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n413_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n385_), .A2(new_n381_), .ZN(new_n420_));
  OAI22_X1  g219(.A1(new_n394_), .A2(KEYINPUT91), .B1(G169gat), .B2(G176gat), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n421_), .B1(KEYINPUT91), .B2(new_n394_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n393_), .A2(new_n384_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n420_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n418_), .B1(new_n419_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n414_), .A2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT20), .B1(new_n397_), .B2(new_n413_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT92), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n429_), .B1(new_n419_), .B2(new_n425_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n413_), .A2(KEYINPUT92), .A3(new_n424_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n428_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n427_), .B1(new_n432_), .B2(new_n417_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G8gat), .B(G36gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT18), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G64gat), .B(G92gat), .ZN(new_n436_));
  XOR2_X1   g235(.A(new_n435_), .B(new_n436_), .Z(new_n437_));
  XNOR2_X1  g236(.A(new_n433_), .B(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(G141gat), .A2(G148gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT3), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G141gat), .A2(G148gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT2), .ZN(new_n442_));
  AOI21_X1  g241(.A(KEYINPUT86), .B1(new_n440_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G155gat), .A2(G162gat), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(G155gat), .A2(G162gat), .ZN(new_n446_));
  NOR3_X1   g245(.A1(new_n443_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n440_), .A2(KEYINPUT86), .A3(new_n442_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  OR2_X1    g248(.A1(new_n444_), .A2(KEYINPUT1), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT85), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n444_), .B1(new_n446_), .B2(KEYINPUT1), .ZN(new_n452_));
  OR2_X1    g251(.A1(new_n452_), .A2(KEYINPUT84), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(KEYINPUT84), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n451_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n439_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n441_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n449_), .A2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G127gat), .B(G134gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G113gat), .B(G120gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n458_), .A2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n449_), .A2(new_n457_), .A3(new_n461_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n463_), .A2(KEYINPUT4), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT93), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G225gat), .A2(G233gat), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n461_), .B1(new_n449_), .B2(new_n457_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT4), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n467_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n465_), .A2(new_n466_), .A3(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n463_), .A2(new_n464_), .A3(new_n467_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(G1gat), .B(G29gat), .Z(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G57gat), .B(G85gat), .ZN(new_n478_));
  XOR2_X1   g277(.A(new_n477_), .B(new_n478_), .Z(new_n479_));
  NAND2_X1  g278(.A1(new_n465_), .A2(new_n470_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(KEYINPUT93), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n474_), .A2(KEYINPUT33), .A3(new_n479_), .A4(new_n481_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n481_), .A2(new_n479_), .A3(new_n472_), .A4(new_n471_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT33), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n479_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n463_), .A2(new_n464_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n465_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n467_), .B1(new_n463_), .B2(KEYINPUT4), .ZN(new_n489_));
  OAI221_X1 g288(.A(new_n486_), .B1(new_n487_), .B2(new_n467_), .C1(new_n488_), .C2(new_n489_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n438_), .A2(new_n482_), .A3(new_n485_), .A4(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n437_), .A2(KEYINPUT32), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n432_), .A2(new_n417_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT95), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n413_), .B1(new_n494_), .B2(new_n424_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n495_), .B1(new_n494_), .B2(new_n424_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(new_n414_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(new_n418_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n492_), .B1(new_n493_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n433_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n499_), .B1(new_n500_), .B2(new_n492_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n466_), .B1(new_n465_), .B2(new_n470_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n486_), .B1(new_n473_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(new_n483_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n501_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n491_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT82), .B(G15gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G227gat), .A2(G233gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n397_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n509_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n388_), .A2(new_n396_), .A3(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G71gat), .B(G99gat), .ZN(new_n513_));
  INV_X1    g312(.A(G43gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT30), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT31), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n515_), .B(KEYINPUT30), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT31), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n510_), .A2(new_n512_), .A3(new_n518_), .A4(new_n521_), .ZN(new_n522_));
  AND3_X1   g321(.A1(new_n388_), .A2(new_n396_), .A3(new_n511_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n511_), .B1(new_n388_), .B2(new_n396_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n519_), .A2(new_n520_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n517_), .A2(KEYINPUT31), .ZN(new_n526_));
  OAI22_X1  g325(.A1(new_n523_), .A2(new_n524_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT83), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n522_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n528_), .B1(new_n522_), .B2(new_n527_), .ZN(new_n530_));
  NOR3_X1   g329(.A1(new_n529_), .A2(new_n530_), .A3(new_n461_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n518_), .A2(new_n521_), .ZN(new_n532_));
  NOR3_X1   g331(.A1(new_n532_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n533_));
  AOI22_X1  g332(.A1(new_n510_), .A2(new_n512_), .B1(new_n518_), .B2(new_n521_), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT83), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n522_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n462_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n531_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G228gat), .A2(G233gat), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n539_), .B(G78gat), .Z(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(new_n226_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(G22gat), .B(G50gat), .Z(new_n543_));
  OAI21_X1  g342(.A(new_n543_), .B1(new_n458_), .B2(KEYINPUT29), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT29), .ZN(new_n545_));
  INV_X1    g344(.A(new_n543_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n449_), .A2(new_n457_), .A3(new_n545_), .A4(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n542_), .B1(new_n544_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n545_), .B1(new_n449_), .B2(new_n457_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n551_));
  OR3_X1    g350(.A1(new_n550_), .A2(new_n419_), .A3(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n551_), .B1(new_n550_), .B2(new_n419_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n544_), .A2(new_n542_), .A3(new_n547_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n549_), .A2(new_n552_), .A3(new_n553_), .A4(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n552_), .A2(new_n553_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n554_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n556_), .B1(new_n557_), .B2(new_n548_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n555_), .A2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n538_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n506_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n437_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n433_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT97), .B(KEYINPUT27), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n433_), .A2(new_n562_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT27), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n493_), .A2(new_n498_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(new_n562_), .ZN(new_n569_));
  AOI22_X1  g368(.A1(new_n563_), .A2(new_n564_), .B1(new_n567_), .B2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n504_), .A2(KEYINPUT96), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n559_), .B1(new_n531_), .B2(new_n537_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n461_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n535_), .A2(new_n462_), .A3(new_n536_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n573_), .A2(new_n574_), .A3(new_n555_), .A4(new_n558_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n572_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT96), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n503_), .A2(new_n577_), .A3(new_n483_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n570_), .A2(new_n571_), .A3(new_n576_), .A4(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n378_), .B1(new_n561_), .B2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n330_), .A2(new_n358_), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n571_), .A2(new_n578_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n581_), .A2(G1gat), .A3(new_n583_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n291_), .A2(new_n283_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(new_n561_), .B2(new_n579_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n356_), .A2(new_n357_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n328_), .ZN(new_n588_));
  NOR3_X1   g387(.A1(new_n587_), .A2(new_n378_), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n586_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n296_), .B1(new_n591_), .B2(new_n582_), .ZN(new_n592_));
  OAI21_X1  g391(.A(KEYINPUT38), .B1(new_n584_), .B2(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n593_), .B1(KEYINPUT38), .B2(new_n584_), .ZN(G1324gat));
  INV_X1    g393(.A(new_n570_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n591_), .A2(KEYINPUT98), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT98), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n597_), .B1(new_n590_), .B2(new_n570_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n596_), .A2(G8gat), .A3(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(KEYINPUT99), .A2(KEYINPUT39), .ZN(new_n600_));
  AND2_X1   g399(.A1(KEYINPUT99), .A2(KEYINPUT39), .ZN(new_n601_));
  OR3_X1    g400(.A1(new_n599_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n599_), .A2(new_n600_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n581_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n604_), .A2(new_n297_), .A3(new_n595_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n606_));
  AND4_X1   g405(.A1(new_n602_), .A2(new_n603_), .A3(new_n605_), .A4(new_n606_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n603_), .A2(new_n605_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n606_), .B1(new_n608_), .B2(new_n602_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n607_), .A2(new_n609_), .ZN(G1325gat));
  INV_X1    g409(.A(G15gat), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n611_), .B1(new_n591_), .B2(new_n538_), .ZN(new_n612_));
  XOR2_X1   g411(.A(KEYINPUT101), .B(KEYINPUT41), .Z(new_n613_));
  OR2_X1    g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n604_), .A2(new_n611_), .A3(new_n538_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n613_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n614_), .A2(new_n615_), .A3(new_n616_), .ZN(G1326gat));
  INV_X1    g416(.A(new_n559_), .ZN(new_n618_));
  OAI21_X1  g417(.A(G22gat), .B1(new_n590_), .B2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT42), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n618_), .A2(G22gat), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n620_), .B1(new_n581_), .B2(new_n621_), .ZN(G1327gat));
  INV_X1    g421(.A(KEYINPUT103), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n500_), .A2(new_n437_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n564_), .B1(new_n624_), .B2(new_n565_), .ZN(new_n625_));
  OAI211_X1 g424(.A(new_n569_), .B(KEYINPUT27), .C1(new_n562_), .C2(new_n433_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n575_), .ZN(new_n627_));
  AOI22_X1  g426(.A1(new_n573_), .A2(new_n574_), .B1(new_n555_), .B2(new_n558_), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n625_), .B(new_n626_), .C1(new_n627_), .C2(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n629_), .A2(new_n582_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n538_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(new_n618_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n632_), .B1(new_n491_), .B2(new_n505_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n377_), .B1(new_n630_), .B2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n358_), .A2(new_n585_), .A3(new_n588_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n623_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n585_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n587_), .A2(new_n637_), .A3(new_n328_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n580_), .A2(KEYINPUT103), .A3(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n636_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(G29gat), .B1(new_n641_), .B2(new_n582_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT44), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT43), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n561_), .A2(new_n579_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n294_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n644_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  AOI211_X1 g446(.A(KEYINPUT43), .B(new_n294_), .C1(new_n561_), .C2(new_n579_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n358_), .A2(new_n377_), .A3(new_n588_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n643_), .B1(new_n649_), .B2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n650_), .B(KEYINPUT102), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n654_), .B(KEYINPUT44), .C1(new_n647_), .C2(new_n648_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n582_), .A2(G29gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n642_), .B1(new_n657_), .B2(new_n658_), .ZN(G1328gat));
  XNOR2_X1  g458(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n653_), .A2(new_n655_), .A3(new_n595_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(G36gat), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n570_), .A2(G36gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n636_), .A2(new_n639_), .A3(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT45), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n636_), .A2(new_n639_), .A3(KEYINPUT45), .A4(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n662_), .A2(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n660_), .B1(new_n670_), .B2(KEYINPUT104), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n668_), .B1(new_n661_), .B2(G36gat), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n673_));
  INV_X1    g472(.A(new_n660_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n672_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n671_), .A2(new_n675_), .ZN(G1329gat));
  XNOR2_X1  g475(.A(KEYINPUT106), .B(G43gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n677_), .B1(new_n640_), .B2(new_n631_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n538_), .A2(G43gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n678_), .B1(new_n656_), .B2(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n680_), .B(new_n681_), .Z(G1330gat));
  AOI21_X1  g481(.A(G50gat), .B1(new_n641_), .B2(new_n559_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n559_), .A2(G50gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n657_), .B2(new_n684_), .ZN(G1331gat));
  INV_X1    g484(.A(G57gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n377_), .B1(new_n561_), .B2(new_n579_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n330_), .A2(new_n587_), .A3(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n686_), .B1(new_n688_), .B2(new_n583_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT108), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n378_), .A2(new_n328_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n358_), .A2(new_n691_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n586_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n694_), .A2(new_n686_), .A3(new_n583_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n690_), .A2(new_n695_), .ZN(G1332gat));
  NAND2_X1  g495(.A1(new_n693_), .A2(new_n595_), .ZN(new_n697_));
  XOR2_X1   g496(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n698_));
  AND3_X1   g497(.A1(new_n697_), .A2(G64gat), .A3(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n697_), .B2(G64gat), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n570_), .A2(G64gat), .ZN(new_n701_));
  OAI22_X1  g500(.A1(new_n699_), .A2(new_n700_), .B1(new_n688_), .B2(new_n701_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT110), .Z(G1333gat));
  OR3_X1    g502(.A1(new_n688_), .A2(G71gat), .A3(new_n631_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n693_), .A2(new_n538_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(G71gat), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n706_), .A2(KEYINPUT49), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(KEYINPUT49), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n704_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT111), .Z(G1334gat));
  OAI21_X1  g509(.A(G78gat), .B1(new_n694_), .B2(new_n618_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT50), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n618_), .A2(G78gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n712_), .B1(new_n688_), .B2(new_n713_), .ZN(G1335gat));
  NOR3_X1   g513(.A1(new_n358_), .A2(new_n377_), .A3(new_n328_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n715_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n716_));
  OAI21_X1  g515(.A(G85gat), .B1(new_n716_), .B2(new_n583_), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n358_), .A2(new_n637_), .A3(new_n328_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n687_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(new_n235_), .A3(new_n582_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n717_), .A2(new_n721_), .ZN(G1336gat));
  OAI21_X1  g521(.A(new_n236_), .B1(new_n719_), .B2(new_n570_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT112), .Z(new_n724_));
  NOR3_X1   g523(.A1(new_n716_), .A2(new_n236_), .A3(new_n570_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1337gat));
  OAI21_X1  g525(.A(G99gat), .B1(new_n716_), .B2(new_n631_), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n720_), .A2(new_n250_), .A3(new_n251_), .A4(new_n538_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT51), .ZN(new_n729_));
  AOI22_X1  g528(.A1(new_n727_), .A2(new_n728_), .B1(KEYINPUT113), .B2(new_n729_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(KEYINPUT113), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n730_), .B(new_n731_), .ZN(G1338gat));
  NOR2_X1   g531(.A1(new_n716_), .A2(new_n618_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n733_), .A2(new_n226_), .ZN(new_n734_));
  XOR2_X1   g533(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n720_), .A2(new_n226_), .A3(new_n559_), .ZN(new_n737_));
  OR2_X1    g536(.A1(KEYINPUT114), .A2(KEYINPUT52), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n736_), .B(new_n737_), .C1(new_n734_), .C2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n734_), .A2(new_n738_), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n743_), .A2(new_n736_), .A3(new_n737_), .A4(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1339gat));
  INV_X1    g544(.A(KEYINPUT122), .ZN(new_n746_));
  INV_X1    g545(.A(G113gat), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n378_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT59), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT54), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT116), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n691_), .B1(new_n288_), .B2(new_n293_), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n358_), .A2(new_n752_), .A3(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n752_), .B1(new_n358_), .B2(new_n753_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n358_), .A2(new_n753_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT116), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n358_), .A2(new_n752_), .A3(new_n753_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n758_), .A2(new_n759_), .A3(KEYINPUT54), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n756_), .A2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n359_), .A2(new_n361_), .A3(new_n366_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n373_), .B1(new_n365_), .B2(new_n362_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n376_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT119), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT119), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n376_), .A2(new_n764_), .A3(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n353_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT117), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n343_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT55), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n343_), .A2(new_n772_), .A3(new_n775_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n334_), .A2(new_n340_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n333_), .A2(new_n342_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n337_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT118), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  OAI211_X1 g580(.A(KEYINPUT118), .B(new_n337_), .C1(new_n777_), .C2(new_n778_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n774_), .A2(new_n776_), .A3(new_n781_), .A4(new_n782_), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n783_), .A2(KEYINPUT56), .A3(new_n350_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT56), .B1(new_n783_), .B2(new_n350_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n771_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT58), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n294_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n771_), .B(KEYINPUT58), .C1(new_n784_), .C2(new_n785_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n789_), .A2(KEYINPUT120), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT120), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n781_), .A2(new_n776_), .A3(new_n782_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n775_), .B1(new_n343_), .B2(new_n772_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n350_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT56), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n783_), .A2(KEYINPUT56), .A3(new_n350_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n770_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n791_), .B1(new_n798_), .B2(KEYINPUT58), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n788_), .B1(new_n790_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT57), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n585_), .B1(KEYINPUT121), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n377_), .A2(new_n353_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n803_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n354_), .A2(new_n769_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n802_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n801_), .A2(KEYINPUT121), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n802_), .B(new_n807_), .C1(new_n804_), .C2(new_n805_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n800_), .A2(new_n809_), .A3(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n761_), .B1(new_n811_), .B2(new_n588_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n583_), .A2(new_n595_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n627_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n750_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n809_), .A2(new_n810_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n646_), .B1(new_n798_), .B2(KEYINPUT58), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n789_), .A2(KEYINPUT120), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n798_), .A2(new_n791_), .A3(KEYINPUT58), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n817_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n588_), .B1(new_n816_), .B2(new_n820_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n756_), .A2(new_n760_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n814_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(KEYINPUT59), .A3(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n749_), .B1(new_n815_), .B2(new_n825_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n812_), .A2(new_n814_), .ZN(new_n827_));
  AOI21_X1  g626(.A(G113gat), .B1(new_n827_), .B2(new_n377_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n746_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(KEYINPUT59), .B1(new_n823_), .B2(new_n824_), .ZN(new_n830_));
  AOI211_X1 g629(.A(new_n750_), .B(new_n814_), .C1(new_n821_), .C2(new_n822_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n748_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n823_), .A2(new_n824_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n747_), .B1(new_n833_), .B2(new_n378_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n832_), .A2(KEYINPUT122), .A3(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n829_), .A2(new_n835_), .ZN(G1340gat));
  INV_X1    g635(.A(G120gat), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(new_n358_), .B2(KEYINPUT60), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n827_), .B(new_n838_), .C1(KEYINPUT60), .C2(new_n837_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n358_), .B1(new_n815_), .B2(new_n825_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n840_), .B2(new_n837_), .ZN(G1341gat));
  INV_X1    g640(.A(G127gat), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n827_), .A2(new_n842_), .A3(new_n328_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n588_), .B1(new_n815_), .B2(new_n825_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(new_n842_), .ZN(G1342gat));
  INV_X1    g644(.A(G134gat), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n827_), .A2(new_n846_), .A3(new_n585_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n294_), .B1(new_n815_), .B2(new_n825_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n847_), .B1(new_n848_), .B2(new_n846_), .ZN(G1343gat));
  NAND2_X1  g648(.A1(new_n813_), .A2(new_n628_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n823_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n377_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g654(.A1(new_n853_), .A2(new_n587_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g656(.A(KEYINPUT123), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n852_), .B2(new_n588_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n823_), .A2(KEYINPUT123), .A3(new_n328_), .A4(new_n851_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT61), .B(G155gat), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n859_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n861_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(G1346gat));
  OR3_X1    g663(.A1(new_n852_), .A2(G162gat), .A3(new_n637_), .ZN(new_n865_));
  OAI21_X1  g664(.A(G162gat), .B1(new_n852_), .B2(new_n294_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(G1347gat));
  NOR2_X1   g666(.A1(new_n582_), .A2(new_n570_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n869_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT22), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n870_), .A2(new_n871_), .A3(new_n627_), .A4(new_n377_), .ZN(new_n872_));
  INV_X1    g671(.A(G169gat), .ZN(new_n873_));
  AND3_X1   g672(.A1(new_n872_), .A2(KEYINPUT62), .A3(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n872_), .A2(KEYINPUT62), .ZN(new_n875_));
  NOR4_X1   g674(.A1(new_n812_), .A2(new_n575_), .A3(new_n378_), .A4(new_n869_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT62), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n873_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n874_), .B1(new_n875_), .B2(new_n878_), .ZN(G1348gat));
  NAND2_X1  g678(.A1(new_n870_), .A2(new_n627_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n880_), .A2(new_n358_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(KEYINPUT124), .B(G176gat), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n881_), .B(new_n882_), .ZN(G1349gat));
  INV_X1    g682(.A(new_n880_), .ZN(new_n884_));
  AOI21_X1  g683(.A(G183gat), .B1(new_n884_), .B2(new_n328_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n880_), .A2(new_n389_), .A3(new_n588_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1350gat));
  OAI21_X1  g686(.A(G190gat), .B1(new_n880_), .B2(new_n294_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n585_), .A2(new_n390_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n880_), .B2(new_n889_), .ZN(G1351gat));
  NAND2_X1  g689(.A1(new_n870_), .A2(new_n628_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n378_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(KEYINPUT125), .B(G197gat), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n892_), .B(new_n893_), .ZN(G1352gat));
  NOR2_X1   g693(.A1(new_n891_), .A2(new_n358_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(new_n400_), .ZN(G1353gat));
  NAND2_X1  g695(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n328_), .A2(new_n897_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(KEYINPUT126), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n891_), .A2(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n900_), .B(new_n901_), .ZN(G1354gat));
  INV_X1    g701(.A(G218gat), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n891_), .A2(new_n903_), .A3(new_n294_), .ZN(new_n904_));
  NOR4_X1   g703(.A1(new_n812_), .A2(new_n637_), .A3(new_n572_), .A4(new_n869_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT127), .ZN(new_n906_));
  AOI21_X1  g705(.A(G218gat), .B1(new_n905_), .B2(new_n906_), .ZN(new_n907_));
  OAI21_X1  g706(.A(KEYINPUT127), .B1(new_n891_), .B2(new_n637_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n904_), .B1(new_n907_), .B2(new_n908_), .ZN(G1355gat));
endmodule


