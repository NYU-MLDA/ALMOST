//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 1 0 0 0 1 0 1 1 1 1 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 0 1 1 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n605_,
    new_n606_, new_n607_, new_n608_, new_n609_, new_n610_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n810_, new_n811_, new_n812_, new_n814_,
    new_n815_, new_n817_, new_n818_, new_n819_, new_n821_, new_n822_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n849_, new_n850_, new_n852_,
    new_n853_, new_n854_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT87), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT1), .ZN(new_n209_));
  OAI211_X1 g008(.A(new_n204_), .B(new_n205_), .C1(new_n207_), .C2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT3), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n203_), .B(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n205_), .B(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n208_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n210_), .B1(new_n215_), .B2(new_n207_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n216_), .A2(KEYINPUT29), .ZN(new_n217_));
  XOR2_X1   g016(.A(new_n217_), .B(KEYINPUT28), .Z(new_n218_));
  XNOR2_X1  g017(.A(G22gat), .B(G50gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n218_), .B(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G211gat), .A2(G218gat), .ZN(new_n222_));
  AND2_X1   g021(.A1(G211gat), .A2(G218gat), .ZN(new_n223_));
  XOR2_X1   g022(.A(G197gat), .B(G204gat), .Z(new_n224_));
  OAI221_X1 g023(.A(KEYINPUT88), .B1(new_n222_), .B2(new_n223_), .C1(new_n224_), .C2(KEYINPUT21), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(KEYINPUT21), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n225_), .B(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n227_), .B1(KEYINPUT29), .B2(new_n216_), .ZN(new_n228_));
  AND2_X1   g027(.A1(G228gat), .A2(G233gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n230_), .A2(KEYINPUT89), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n230_), .A2(KEYINPUT89), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n221_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G78gat), .B(G106gat), .Z(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n218_), .B(new_n219_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n230_), .A2(KEYINPUT89), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  AND3_X1   g037(.A1(new_n233_), .A2(new_n235_), .A3(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n235_), .B1(new_n233_), .B2(new_n238_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G113gat), .B(G120gat), .ZN(new_n242_));
  INV_X1    g041(.A(G134gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT86), .B(G127gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G169gat), .A2(G176gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT22), .B(G169gat), .ZN(new_n249_));
  INV_X1    g048(.A(G176gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  AND2_X1   g050(.A1(G183gat), .A2(G190gat), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT23), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT84), .B(KEYINPUT23), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n254_), .B1(new_n252_), .B2(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(G183gat), .A2(G190gat), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n248_), .B(new_n251_), .C1(new_n256_), .C2(new_n257_), .ZN(new_n258_));
  OR2_X1    g057(.A1(G169gat), .A2(G176gat), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n259_), .A2(new_n248_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT24), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT25), .B(G183gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT26), .B(G190gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n261_), .A2(new_n264_), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n265_), .A2(KEYINPUT83), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(KEYINPUT83), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n252_), .A2(new_n253_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n268_), .B1(new_n255_), .B2(new_n252_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n266_), .A2(new_n267_), .A3(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n259_), .A2(KEYINPUT24), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n258_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n272_), .A2(KEYINPUT30), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n272_), .A2(KEYINPUT30), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT85), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT31), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G15gat), .B(G43gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G227gat), .A2(G233gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G71gat), .B(G99gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n275_), .A2(new_n276_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n276_), .B1(new_n275_), .B2(new_n281_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n247_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n275_), .A2(new_n281_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT31), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n287_), .A2(new_n246_), .A3(new_n282_), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n273_), .A2(new_n274_), .A3(KEYINPUT85), .ZN(new_n289_));
  AND3_X1   g088(.A1(new_n285_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n289_), .B1(new_n285_), .B2(new_n288_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n241_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n232_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n236_), .B1(new_n293_), .B2(new_n237_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n238_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n234_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n233_), .A2(new_n235_), .A3(new_n238_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n289_), .ZN(new_n299_));
  NOR3_X1   g098(.A1(new_n283_), .A2(new_n284_), .A3(new_n247_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n246_), .B1(new_n287_), .B2(new_n282_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n299_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n285_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n298_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT97), .ZN(new_n305_));
  XOR2_X1   g104(.A(KEYINPUT90), .B(KEYINPUT24), .Z(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n307_), .A2(new_n259_), .ZN(new_n308_));
  OR3_X1    g107(.A1(new_n308_), .A2(KEYINPUT91), .A3(new_n256_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n260_), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT91), .B1(new_n308_), .B2(new_n256_), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n309_), .A2(new_n264_), .A3(new_n310_), .A4(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n269_), .B1(G183gat), .B2(G190gat), .ZN(new_n313_));
  XOR2_X1   g112(.A(new_n249_), .B(KEYINPUT92), .Z(new_n314_));
  OAI211_X1 g113(.A(new_n248_), .B(new_n313_), .C1(new_n314_), .C2(G176gat), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n312_), .A2(new_n227_), .A3(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT20), .ZN(new_n317_));
  INV_X1    g116(.A(new_n227_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n272_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT93), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n272_), .A2(KEYINPUT93), .A3(new_n318_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n317_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G226gat), .A2(G233gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT19), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n323_), .A2(new_n326_), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n272_), .A2(new_n318_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n312_), .A2(new_n315_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n318_), .ZN(new_n330_));
  AND4_X1   g129(.A1(KEYINPUT20), .A2(new_n328_), .A3(new_n326_), .A4(new_n330_), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n327_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G8gat), .B(G36gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(G92gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT18), .B(G64gat), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n335_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT96), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n305_), .B1(new_n332_), .B2(new_n339_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n305_), .B(new_n339_), .C1(new_n327_), .C2(new_n331_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n328_), .A2(KEYINPUT20), .A3(new_n325_), .A4(new_n330_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n342_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n338_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n341_), .A2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT27), .B1(new_n340_), .B2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n343_), .B(new_n338_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT27), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  AOI22_X1  g149(.A1(new_n292_), .A2(new_n304_), .B1(new_n347_), .B2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n246_), .B(new_n216_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G225gat), .A2(G233gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT4), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n246_), .A2(new_n356_), .A3(new_n216_), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n354_), .B(KEYINPUT94), .Z(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n357_), .B(new_n359_), .C1(new_n352_), .C2(new_n356_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n355_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G1gat), .B(G29gat), .ZN(new_n362_));
  INV_X1    g161(.A(G85gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT0), .B(G57gat), .ZN(new_n365_));
  XOR2_X1   g164(.A(new_n364_), .B(new_n365_), .Z(new_n366_));
  NAND2_X1  g165(.A1(new_n361_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n366_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n355_), .A2(new_n360_), .A3(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT33), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n369_), .A2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT95), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n369_), .A2(new_n372_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n352_), .A2(new_n356_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n357_), .A2(new_n354_), .ZN(new_n377_));
  OAI221_X1 g176(.A(new_n366_), .B1(new_n352_), .B2(new_n358_), .C1(new_n376_), .C2(new_n377_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n348_), .A2(new_n374_), .A3(new_n375_), .A4(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n332_), .A2(KEYINPUT32), .A3(new_n344_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT32), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n343_), .B1(new_n381_), .B2(new_n338_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n380_), .A2(new_n370_), .A3(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n298_), .B1(new_n379_), .B2(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n290_), .A2(new_n291_), .ZN(new_n385_));
  AOI22_X1  g184(.A1(new_n351_), .A2(new_n371_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G57gat), .B(G64gat), .ZN(new_n387_));
  OR2_X1    g186(.A1(new_n387_), .A2(KEYINPUT11), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(KEYINPUT11), .ZN(new_n389_));
  XOR2_X1   g188(.A(G71gat), .B(G78gat), .Z(new_n390_));
  NAND3_X1  g189(.A1(new_n388_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  OR2_X1    g190(.A1(new_n389_), .A2(new_n390_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G231gat), .A2(G233gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(G8gat), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n396_), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n397_), .A2(KEYINPUT79), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G15gat), .B(G22gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(KEYINPUT79), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n398_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G1gat), .B(G8gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT80), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n401_), .A2(new_n403_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n395_), .B(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT17), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G127gat), .B(G155gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(G211gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT16), .B(G183gat), .ZN(new_n411_));
  XOR2_X1   g210(.A(new_n410_), .B(new_n411_), .Z(new_n412_));
  NOR3_X1   g211(.A1(new_n407_), .A2(new_n408_), .A3(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(KEYINPUT17), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n413_), .B1(new_n407_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n386_), .A2(new_n416_), .ZN(new_n417_));
  AND2_X1   g216(.A1(G230gat), .A2(G233gat), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT68), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT7), .ZN(new_n420_));
  INV_X1    g219(.A(G99gat), .ZN(new_n421_));
  INV_X1    g220(.A(G106gat), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n420_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G99gat), .A2(G106gat), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT6), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n423_), .A2(new_n426_), .A3(new_n427_), .A4(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(KEYINPUT67), .A2(KEYINPUT8), .ZN(new_n430_));
  XOR2_X1   g229(.A(G85gat), .B(G92gat), .Z(new_n431_));
  AND3_X1   g230(.A1(new_n429_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n430_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n435_), .B1(G85gat), .B2(G92gat), .ZN(new_n436_));
  OR2_X1    g235(.A1(KEYINPUT66), .A2(G92gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n363_), .A2(KEYINPUT65), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT65), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(G85gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(KEYINPUT66), .A2(G92gat), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n437_), .A2(new_n438_), .A3(new_n440_), .A4(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(KEYINPUT64), .B(KEYINPUT9), .Z(new_n443_));
  AOI21_X1  g242(.A(new_n436_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n426_), .A2(new_n427_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT10), .B(G99gat), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n446_), .A2(G106gat), .ZN(new_n447_));
  NOR3_X1   g246(.A1(new_n444_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n419_), .B1(new_n434_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n447_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n445_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n452_));
  INV_X1    g251(.A(new_n441_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(KEYINPUT66), .A2(G92gat), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT65), .B(G85gat), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n452_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n450_), .B(new_n451_), .C1(new_n457_), .C2(new_n436_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n458_), .B(KEYINPUT68), .C1(new_n433_), .C2(new_n432_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n449_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(new_n393_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT69), .ZN(new_n462_));
  INV_X1    g261(.A(new_n393_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n449_), .A2(new_n463_), .A3(new_n459_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT70), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n418_), .B1(new_n462_), .B2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT71), .B1(new_n432_), .B2(new_n433_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n429_), .A2(new_n431_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n430_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT71), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n429_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n470_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n467_), .A2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT72), .B1(new_n474_), .B2(new_n458_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT72), .ZN(new_n476_));
  AOI211_X1 g275(.A(new_n476_), .B(new_n448_), .C1(new_n467_), .C2(new_n473_), .ZN(new_n477_));
  OAI211_X1 g276(.A(KEYINPUT12), .B(new_n463_), .C1(new_n475_), .C2(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n418_), .B1(new_n460_), .B2(new_n393_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT73), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT12), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n464_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n480_), .B1(new_n464_), .B2(new_n481_), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n478_), .B(new_n479_), .C1(new_n482_), .C2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n466_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G120gat), .B(G148gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(G204gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT5), .B(G176gat), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n487_), .B(new_n488_), .Z(new_n489_));
  NAND2_X1  g288(.A1(new_n485_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n489_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n466_), .A2(new_n484_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT13), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G29gat), .B(G36gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G43gat), .B(G50gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT15), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n406_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G229gat), .A2(G233gat), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n404_), .A2(new_n498_), .A3(new_n405_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT82), .ZN(new_n504_));
  INV_X1    g303(.A(new_n501_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n502_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n498_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n505_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT82), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n500_), .A2(new_n509_), .A3(new_n501_), .A4(new_n502_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n504_), .A2(new_n508_), .A3(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G113gat), .B(G141gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G169gat), .B(G197gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n511_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n514_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n504_), .A2(new_n508_), .A3(new_n510_), .A4(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT35), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G232gat), .A2(G233gat), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n521_), .B(KEYINPUT34), .Z(new_n522_));
  INV_X1    g321(.A(new_n498_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n523_), .B1(new_n449_), .B2(new_n459_), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n432_), .A2(new_n433_), .A3(KEYINPUT71), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n471_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n458_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n476_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n474_), .A2(KEYINPUT72), .A3(new_n458_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n524_), .B1(new_n530_), .B2(new_n499_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT74), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n522_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n499_), .B1(new_n475_), .B2(new_n477_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n524_), .ZN(new_n535_));
  AND4_X1   g334(.A1(new_n532_), .A2(new_n534_), .A3(new_n535_), .A4(new_n522_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n520_), .B1(new_n533_), .B2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n531_), .A2(new_n532_), .A3(new_n522_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n534_), .A2(new_n532_), .A3(new_n535_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n522_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n531_), .A2(new_n520_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n538_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G190gat), .B(G218gat), .ZN(new_n544_));
  INV_X1    g343(.A(G162gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT75), .B(G134gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n548_), .B(KEYINPUT36), .Z(new_n549_));
  NAND3_X1  g348(.A1(new_n537_), .A2(new_n543_), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT77), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n548_), .A2(KEYINPUT36), .ZN(new_n552_));
  INV_X1    g351(.A(new_n543_), .ZN(new_n553_));
  AOI21_X1  g352(.A(KEYINPUT35), .B1(new_n538_), .B2(new_n541_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n552_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT77), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n537_), .A2(new_n556_), .A3(new_n543_), .A4(new_n549_), .ZN(new_n557_));
  AND3_X1   g356(.A1(new_n551_), .A2(new_n555_), .A3(new_n557_), .ZN(new_n558_));
  NOR3_X1   g357(.A1(new_n495_), .A2(new_n519_), .A3(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n417_), .A2(new_n559_), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n560_), .B(KEYINPUT100), .Z(new_n561_));
  AOI21_X1  g360(.A(new_n202_), .B1(new_n561_), .B2(new_n370_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT101), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(KEYINPUT78), .B(KEYINPUT37), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n551_), .A2(new_n555_), .A3(new_n557_), .A4(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n549_), .B(KEYINPUT76), .Z(new_n567_));
  NOR3_X1   g366(.A1(new_n553_), .A2(new_n554_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n552_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n569_), .B1(new_n537_), .B2(new_n543_), .ZN(new_n570_));
  OAI21_X1  g369(.A(KEYINPUT37), .B1(new_n568_), .B2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n566_), .A2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n572_), .A2(new_n494_), .A3(new_n415_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT81), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT98), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n575_), .B1(new_n386_), .B2(new_n519_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n292_), .A2(new_n304_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n347_), .A2(new_n350_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n577_), .A2(new_n371_), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n384_), .A2(new_n385_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n581_), .A2(KEYINPUT98), .A3(new_n518_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n574_), .B1(new_n576_), .B2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n583_), .A2(new_n202_), .A3(new_n370_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT38), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n586_), .B(KEYINPUT99), .Z(new_n587_));
  NAND2_X1  g386(.A1(new_n584_), .A2(new_n585_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT102), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n564_), .A2(new_n587_), .A3(new_n589_), .ZN(G1324gat));
  OR3_X1    g389(.A1(new_n560_), .A2(KEYINPUT103), .A3(new_n578_), .ZN(new_n591_));
  OAI21_X1  g390(.A(KEYINPUT103), .B1(new_n560_), .B2(new_n578_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n591_), .A2(G8gat), .A3(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT39), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT39), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n591_), .A2(new_n595_), .A3(new_n592_), .A4(G8gat), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n578_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n583_), .A2(new_n396_), .A3(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT40), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n597_), .A2(KEYINPUT40), .A3(new_n599_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(G1325gat));
  INV_X1    g403(.A(G15gat), .ZN(new_n605_));
  INV_X1    g404(.A(new_n385_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n605_), .B1(new_n561_), .B2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n583_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(G1326gat));
  INV_X1    g410(.A(G22gat), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n612_), .B1(new_n561_), .B2(new_n298_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT42), .Z(new_n614_));
  NAND3_X1  g413(.A1(new_n583_), .A2(new_n612_), .A3(new_n298_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(G1327gat));
  INV_X1    g415(.A(new_n558_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n617_), .A2(new_n415_), .ZN(new_n618_));
  AOI21_X1  g417(.A(KEYINPUT98), .B1(new_n581_), .B2(new_n518_), .ZN(new_n619_));
  AOI211_X1 g418(.A(new_n575_), .B(new_n519_), .C1(new_n579_), .C2(new_n580_), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n494_), .B(new_n618_), .C1(new_n619_), .C2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT107), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n576_), .A2(new_n582_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT107), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n623_), .A2(new_n624_), .A3(new_n494_), .A4(new_n618_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n622_), .A2(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(G29gat), .B1(new_n626_), .B2(new_n370_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT105), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n628_), .B1(new_n386_), .B2(new_n572_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(KEYINPUT43), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT43), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n628_), .B(new_n631_), .C1(new_n386_), .C2(new_n572_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n495_), .A2(new_n519_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n630_), .A2(new_n632_), .A3(new_n416_), .A4(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT106), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT44), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n634_), .A2(KEYINPUT106), .A3(KEYINPUT44), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n371_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n627_), .B1(new_n639_), .B2(G29gat), .ZN(G1328gat));
  NOR2_X1   g439(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n641_));
  INV_X1    g440(.A(G36gat), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n637_), .A2(new_n638_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n642_), .B1(new_n643_), .B2(new_n598_), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n622_), .A2(new_n642_), .A3(new_n598_), .A4(new_n625_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT45), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n641_), .B1(new_n644_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n638_), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT44), .B1(new_n634_), .B2(KEYINPUT106), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n598_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(G36gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n645_), .B(KEYINPUT45), .ZN(new_n653_));
  INV_X1    g452(.A(new_n641_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n652_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n648_), .A2(new_n655_), .ZN(G1329gat));
  INV_X1    g455(.A(G43gat), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n626_), .A2(new_n657_), .A3(new_n606_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n385_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n658_), .B1(new_n659_), .B2(new_n657_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT47), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  OAI211_X1 g461(.A(KEYINPUT47), .B(new_n658_), .C1(new_n659_), .C2(new_n657_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1330gat));
  OAI21_X1  g463(.A(new_n298_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n665_), .A2(KEYINPUT109), .A3(G50gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT109), .B1(new_n665_), .B2(G50gat), .ZN(new_n667_));
  INV_X1    g466(.A(new_n626_), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n241_), .A2(G50gat), .ZN(new_n669_));
  OAI22_X1  g468(.A1(new_n666_), .A2(new_n667_), .B1(new_n668_), .B2(new_n669_), .ZN(G1331gat));
  NOR2_X1   g469(.A1(new_n494_), .A2(new_n518_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n581_), .A2(new_n671_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n672_), .A2(new_n415_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n673_), .A2(new_n572_), .ZN(new_n674_));
  AOI21_X1  g473(.A(G57gat), .B1(new_n674_), .B2(new_n370_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n673_), .A2(new_n617_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n370_), .A2(G57gat), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n675_), .B1(new_n676_), .B2(new_n677_), .ZN(G1332gat));
  INV_X1    g477(.A(G64gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n679_), .B1(new_n676_), .B2(new_n598_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT48), .Z(new_n681_));
  NAND3_X1  g480(.A1(new_n674_), .A2(new_n679_), .A3(new_n598_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1333gat));
  INV_X1    g482(.A(G71gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n684_), .B1(new_n676_), .B2(new_n606_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n685_), .B(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n674_), .A2(new_n684_), .A3(new_n606_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1334gat));
  INV_X1    g488(.A(G78gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n690_), .B1(new_n676_), .B2(new_n298_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT50), .Z(new_n692_));
  NAND3_X1  g491(.A1(new_n674_), .A2(new_n690_), .A3(new_n298_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1335gat));
  AND2_X1   g493(.A1(new_n672_), .A2(new_n618_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G85gat), .B1(new_n695_), .B2(new_n370_), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n630_), .A2(new_n632_), .A3(new_n416_), .A4(new_n671_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n370_), .A2(new_n456_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n696_), .B1(new_n698_), .B2(new_n699_), .ZN(G1336gat));
  AOI21_X1  g499(.A(G92gat), .B1(new_n695_), .B2(new_n598_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n578_), .A2(new_n454_), .A3(new_n453_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n698_), .B2(new_n702_), .ZN(G1337gat));
  OAI21_X1  g502(.A(G99gat), .B1(new_n697_), .B2(new_n385_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n446_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n695_), .A2(new_n606_), .A3(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n704_), .A2(KEYINPUT111), .A3(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g507(.A1(new_n695_), .A2(new_n422_), .A3(new_n298_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT52), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n698_), .A2(new_n298_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n711_), .B2(G106gat), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n710_), .B(G106gat), .C1(new_n697_), .C2(new_n241_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n709_), .B1(new_n712_), .B2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT53), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT53), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n717_), .B(new_n709_), .C1(new_n712_), .C2(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(G1339gat));
  INV_X1    g518(.A(KEYINPUT58), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT112), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n484_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT55), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n478_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n418_), .B1(new_n462_), .B2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT55), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n484_), .A2(new_n721_), .A3(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n723_), .A2(new_n725_), .A3(new_n727_), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n728_), .A2(KEYINPUT56), .A3(new_n489_), .ZN(new_n729_));
  AOI21_X1  g528(.A(KEYINPUT56), .B1(new_n728_), .B2(new_n489_), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n729_), .A2(new_n730_), .A3(KEYINPUT114), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n501_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n500_), .A2(new_n505_), .A3(new_n502_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(new_n514_), .A3(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n517_), .A2(new_n734_), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT113), .Z(new_n736_));
  INV_X1    g535(.A(new_n492_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n728_), .A2(KEYINPUT114), .A3(KEYINPUT56), .A4(new_n489_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n720_), .B1(new_n731_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n572_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n728_), .A2(new_n489_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT56), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT114), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n728_), .A2(KEYINPUT56), .A3(new_n489_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n745_), .A2(new_n746_), .A3(new_n747_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n748_), .A2(KEYINPUT58), .A3(new_n739_), .A4(new_n738_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n741_), .A2(new_n742_), .A3(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n492_), .A2(new_n518_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n745_), .B2(new_n747_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n736_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n617_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT57), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n751_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n757_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n753_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n760_), .A2(KEYINPUT57), .A3(new_n617_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n750_), .A2(new_n756_), .A3(new_n761_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n572_), .A2(new_n494_), .A3(new_n519_), .A4(new_n415_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT54), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n763_), .A2(KEYINPUT54), .ZN(new_n765_));
  AOI22_X1  g564(.A1(new_n762_), .A2(new_n416_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n578_), .A2(new_n370_), .ZN(new_n767_));
  NOR4_X1   g566(.A1(new_n766_), .A2(new_n385_), .A3(new_n298_), .A4(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(G113gat), .B1(new_n768_), .B2(new_n518_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n762_), .A2(new_n416_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n765_), .A2(new_n764_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n298_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n767_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n772_), .A2(new_n606_), .A3(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT59), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT59), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT115), .B1(new_n768_), .B2(new_n776_), .ZN(new_n777_));
  AOI211_X1 g576(.A(new_n755_), .B(new_n558_), .C1(new_n759_), .C2(new_n758_), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT57), .B1(new_n760_), .B2(new_n617_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n415_), .B1(new_n780_), .B2(new_n750_), .ZN(new_n781_));
  XOR2_X1   g580(.A(new_n763_), .B(KEYINPUT54), .Z(new_n782_));
  OAI211_X1 g581(.A(new_n606_), .B(new_n241_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT115), .ZN(new_n784_));
  NOR4_X1   g583(.A1(new_n783_), .A2(new_n784_), .A3(KEYINPUT59), .A4(new_n767_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n775_), .B1(new_n777_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT116), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n784_), .B1(new_n774_), .B2(KEYINPUT59), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n768_), .A2(KEYINPUT115), .A3(new_n776_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n791_), .A2(KEYINPUT116), .A3(new_n775_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n788_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n518_), .A2(G113gat), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT117), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n769_), .B1(new_n793_), .B2(new_n795_), .ZN(G1340gat));
  INV_X1    g595(.A(G120gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n495_), .B1(new_n768_), .B2(new_n776_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n797_), .B1(new_n791_), .B2(new_n799_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n797_), .A2(KEYINPUT60), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT60), .B1(new_n495_), .B2(new_n797_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n774_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT118), .B1(new_n800_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT118), .ZN(new_n805_));
  INV_X1    g604(.A(new_n803_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n798_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n805_), .B(new_n806_), .C1(new_n807_), .C2(new_n797_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n804_), .A2(new_n808_), .ZN(G1341gat));
  AOI21_X1  g608(.A(G127gat), .B1(new_n768_), .B2(new_n415_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(KEYINPUT119), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n415_), .A2(G127gat), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n793_), .B2(new_n812_), .ZN(G1342gat));
  AOI21_X1  g612(.A(G134gat), .B1(new_n768_), .B2(new_n558_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n572_), .A2(new_n243_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n814_), .B1(new_n793_), .B2(new_n815_), .ZN(G1343gat));
  NOR2_X1   g615(.A1(new_n766_), .A2(new_n304_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n773_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n818_), .A2(new_n519_), .ZN(new_n819_));
  XOR2_X1   g618(.A(new_n819_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g619(.A1(new_n818_), .A2(new_n494_), .ZN(new_n821_));
  XOR2_X1   g620(.A(KEYINPUT120), .B(G148gat), .Z(new_n822_));
  XNOR2_X1  g621(.A(new_n821_), .B(new_n822_), .ZN(G1345gat));
  NOR2_X1   g622(.A1(new_n818_), .A2(new_n416_), .ZN(new_n824_));
  XOR2_X1   g623(.A(KEYINPUT61), .B(G155gat), .Z(new_n825_));
  XNOR2_X1  g624(.A(new_n824_), .B(new_n825_), .ZN(G1346gat));
  OAI21_X1  g625(.A(new_n545_), .B1(new_n818_), .B2(new_n617_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT121), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n818_), .A2(new_n545_), .A3(new_n572_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n828_), .A2(new_n829_), .ZN(G1347gat));
  NOR2_X1   g629(.A1(new_n578_), .A2(new_n370_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n832_), .A2(new_n385_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n772_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n518_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT122), .ZN(new_n837_));
  OR3_X1    g636(.A1(new_n834_), .A2(KEYINPUT122), .A3(new_n519_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(G169gat), .A3(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT62), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n837_), .A2(KEYINPUT62), .A3(G169gat), .A4(new_n838_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n841_), .B(new_n842_), .C1(new_n314_), .C2(new_n836_), .ZN(G1348gat));
  AOI21_X1  g642(.A(G176gat), .B1(new_n835_), .B2(new_n495_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n772_), .B(KEYINPUT123), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n845_), .A2(new_n385_), .A3(new_n832_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n494_), .A2(new_n250_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n844_), .B1(new_n846_), .B2(new_n847_), .ZN(G1349gat));
  AOI21_X1  g647(.A(G183gat), .B1(new_n846_), .B2(new_n415_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n834_), .A2(new_n262_), .A3(new_n416_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1350gat));
  NAND3_X1  g650(.A1(new_n835_), .A2(new_n263_), .A3(new_n558_), .ZN(new_n852_));
  OAI21_X1  g651(.A(G190gat), .B1(new_n834_), .B2(new_n572_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(KEYINPUT124), .ZN(G1351gat));
  INV_X1    g654(.A(new_n304_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n856_), .B(new_n831_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT125), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n518_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n495_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g662(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n864_));
  AOI21_X1  g663(.A(KEYINPUT125), .B1(new_n817_), .B2(new_n831_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n857_), .A2(new_n858_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n415_), .B(new_n864_), .C1(new_n865_), .C2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(KEYINPUT126), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT126), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n859_), .A2(new_n869_), .A3(new_n415_), .A4(new_n864_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n871_));
  AND3_X1   g670(.A1(new_n868_), .A2(new_n870_), .A3(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n871_), .B1(new_n868_), .B2(new_n870_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n872_), .A2(new_n873_), .ZN(G1354gat));
  INV_X1    g673(.A(KEYINPUT127), .ZN(new_n875_));
  AND3_X1   g674(.A1(new_n859_), .A2(new_n875_), .A3(new_n558_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n859_), .B2(new_n558_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n876_), .A2(new_n877_), .A3(G218gat), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n859_), .A2(G218gat), .A3(new_n742_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1355gat));
endmodule


