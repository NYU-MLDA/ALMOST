//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 1 1 0 0 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 1 1 0 1 1 0 0 1 1 0 1 1 1 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n813_, new_n814_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n833_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n857_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_;
  NAND2_X1  g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT84), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT2), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT85), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  OAI211_X1 g009(.A(new_n206_), .B(new_n210_), .C1(new_n205_), .C2(new_n202_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G155gat), .B(G162gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  AND2_X1   g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n209_), .B1(new_n215_), .B2(KEYINPUT1), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n204_), .B(new_n216_), .C1(KEYINPUT1), .C2(new_n212_), .ZN(new_n217_));
  AND2_X1   g016(.A1(new_n214_), .A2(new_n217_), .ZN(new_n218_));
  XOR2_X1   g017(.A(G113gat), .B(G120gat), .Z(new_n219_));
  XNOR2_X1  g018(.A(G127gat), .B(G134gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n219_), .B(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n218_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n214_), .A2(new_n217_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(new_n221_), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT4), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G225gat), .A2(G233gat), .ZN(new_n228_));
  XOR2_X1   g027(.A(new_n228_), .B(KEYINPUT96), .Z(new_n229_));
  INV_X1    g028(.A(KEYINPUT4), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n224_), .A2(new_n230_), .A3(new_n221_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT97), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n232_), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n227_), .A2(new_n229_), .A3(new_n233_), .A4(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n229_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n226_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G1gat), .B(G29gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(G85gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT0), .B(G57gat), .ZN(new_n241_));
  XOR2_X1   g040(.A(new_n240_), .B(new_n241_), .Z(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n238_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n235_), .A2(new_n242_), .A3(new_n237_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(KEYINPUT99), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT99), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n238_), .A2(new_n247_), .A3(new_n243_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT20), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT22), .B(G169gat), .ZN(new_n251_));
  INV_X1    g050(.A(G176gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G169gat), .A2(G176gat), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT83), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G183gat), .A2(G190gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT23), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT80), .B(G183gat), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n258_), .B1(G190gat), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n256_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n258_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(G169gat), .A2(G176gat), .ZN(new_n263_));
  XOR2_X1   g062(.A(new_n263_), .B(KEYINPUT82), .Z(new_n264_));
  INV_X1    g063(.A(KEYINPUT24), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n262_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n254_), .A2(KEYINPUT24), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n259_), .A2(KEYINPUT25), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n268_), .B1(KEYINPUT25), .B2(G183gat), .ZN(new_n269_));
  INV_X1    g068(.A(G190gat), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n269_), .B1(KEYINPUT26), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(KEYINPUT26), .ZN(new_n272_));
  XOR2_X1   g071(.A(new_n272_), .B(KEYINPUT81), .Z(new_n273_));
  OAI221_X1 g072(.A(new_n266_), .B1(new_n264_), .B2(new_n267_), .C1(new_n271_), .C2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n261_), .A2(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(G211gat), .B(G218gat), .Z(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT89), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT21), .ZN(new_n278_));
  INV_X1    g077(.A(G204gat), .ZN(new_n279_));
  AND2_X1   g078(.A1(new_n279_), .A2(G197gat), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(G197gat), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  OR3_X1    g081(.A1(new_n277_), .A2(new_n278_), .A3(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n278_), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n280_), .A2(KEYINPUT87), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n281_), .A2(KEYINPUT88), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n280_), .A2(KEYINPUT87), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n281_), .A2(KEYINPUT88), .ZN(new_n288_));
  AND4_X1   g087(.A1(new_n285_), .A2(new_n286_), .A3(new_n287_), .A4(new_n288_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n277_), .B(new_n284_), .C1(new_n289_), .C2(new_n278_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n283_), .A2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n250_), .B1(new_n275_), .B2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G226gat), .A2(G233gat), .ZN(new_n293_));
  XOR2_X1   g092(.A(new_n293_), .B(KEYINPUT19), .Z(new_n294_));
  OAI21_X1  g093(.A(new_n258_), .B1(G183gat), .B2(G190gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n255_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n267_), .B(KEYINPUT93), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n266_), .B1(new_n264_), .B2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT26), .B(G190gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT92), .ZN(new_n300_));
  XOR2_X1   g099(.A(KEYINPUT25), .B(G183gat), .Z(new_n301_));
  NOR2_X1   g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n296_), .B1(new_n298_), .B2(new_n302_), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n292_), .B(new_n294_), .C1(new_n291_), .C2(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n250_), .B1(new_n291_), .B2(new_n303_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n305_), .B1(new_n275_), .B2(new_n291_), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n294_), .B(KEYINPUT91), .Z(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G8gat), .B(G36gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT95), .ZN(new_n310_));
  XOR2_X1   g109(.A(G64gat), .B(G92gat), .Z(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n304_), .A2(new_n308_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT98), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n303_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n303_), .A2(new_n316_), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n317_), .A2(new_n290_), .A3(new_n283_), .A4(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n294_), .B1(new_n319_), .B2(new_n292_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n306_), .A2(new_n307_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  OAI211_X1 g121(.A(KEYINPUT27), .B(new_n315_), .C1(new_n322_), .C2(new_n314_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT100), .B(KEYINPUT27), .ZN(new_n324_));
  INV_X1    g123(.A(new_n315_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n314_), .B1(new_n304_), .B2(new_n308_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n324_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n323_), .A2(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(G15gat), .B(G43gat), .Z(new_n329_));
  XNOR2_X1  g128(.A(G71gat), .B(G99gat), .ZN(new_n330_));
  XOR2_X1   g129(.A(new_n329_), .B(new_n330_), .Z(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n275_), .A2(KEYINPUT30), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT30), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n261_), .A2(new_n274_), .A3(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n221_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n333_), .A2(new_n222_), .A3(new_n335_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G227gat), .A2(G233gat), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n339_), .B(KEYINPUT31), .Z(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n337_), .A2(new_n338_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n341_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n332_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n337_), .A2(new_n338_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(new_n340_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n347_), .A2(new_n331_), .A3(new_n342_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n345_), .A2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G22gat), .B(G50gat), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT29), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n218_), .A2(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n353_), .A2(KEYINPUT28), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n224_), .A2(KEYINPUT29), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT28), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n351_), .B1(new_n354_), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n353_), .A2(KEYINPUT28), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n355_), .A2(new_n356_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n359_), .A2(new_n360_), .A3(new_n350_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n358_), .A2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n291_), .B1(new_n218_), .B2(new_n352_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT86), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(G228gat), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n364_), .A2(G228gat), .ZN(new_n367_));
  OAI21_X1  g166(.A(G233gat), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n363_), .A2(new_n369_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n291_), .B(new_n368_), .C1(new_n218_), .C2(new_n352_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  XOR2_X1   g171(.A(G78gat), .B(G106gat), .Z(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n362_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT90), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n377_), .B1(new_n358_), .B2(new_n361_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n376_), .B1(new_n375_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n372_), .A2(new_n374_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  AND3_X1   g180(.A1(new_n378_), .A2(new_n372_), .A3(new_n374_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n349_), .A2(new_n381_), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n382_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n385_), .A2(new_n349_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n249_), .B(new_n328_), .C1(new_n384_), .C2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n314_), .A2(KEYINPUT32), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n304_), .A2(new_n308_), .A3(new_n388_), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n322_), .A2(new_n388_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n246_), .A2(new_n248_), .A3(new_n389_), .A4(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n325_), .A2(new_n326_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT33), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n245_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n226_), .A2(new_n229_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n227_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n243_), .B(new_n395_), .C1(new_n396_), .C2(new_n229_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n235_), .A2(KEYINPUT33), .A3(new_n242_), .A4(new_n237_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n392_), .A2(new_n394_), .A3(new_n397_), .A4(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n391_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n385_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n401_), .A2(new_n349_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n387_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT7), .ZN(new_n405_));
  INV_X1    g204(.A(G99gat), .ZN(new_n406_));
  INV_X1    g205(.A(G106gat), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n405_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  AND2_X1   g209(.A1(G99gat), .A2(G106gat), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT65), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n413_), .A2(KEYINPUT6), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT6), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n415_), .A2(KEYINPUT65), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n412_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(KEYINPUT65), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n413_), .A2(KEYINPUT6), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n419_), .A3(new_n411_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n410_), .B1(new_n417_), .B2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G85gat), .B(G92gat), .ZN(new_n422_));
  NOR3_X1   g221(.A1(new_n421_), .A2(KEYINPUT8), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT8), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n408_), .A2(new_n409_), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n418_), .A2(new_n419_), .A3(new_n411_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n411_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n425_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n422_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n424_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT67), .B1(new_n423_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT64), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT10), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n433_), .A2(G99gat), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n406_), .A2(KEYINPUT10), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n432_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n406_), .A2(KEYINPUT10), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n433_), .A2(G99gat), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(KEYINPUT64), .ZN(new_n439_));
  AOI21_X1  g238(.A(G106gat), .B1(new_n436_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT9), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n422_), .A2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n426_), .A2(new_n427_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n441_), .A2(G85gat), .A3(G92gat), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n443_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT8), .B1(new_n421_), .B2(new_n422_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT67), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n428_), .A2(new_n424_), .A3(new_n429_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n431_), .A2(new_n447_), .A3(new_n451_), .ZN(new_n452_));
  XOR2_X1   g251(.A(G71gat), .B(G78gat), .Z(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(G57gat), .ZN(new_n455_));
  INV_X1    g254(.A(G64gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G57gat), .A2(G64gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT11), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT11), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n457_), .A2(new_n461_), .A3(new_n458_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n454_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n453_), .B1(KEYINPUT11), .B2(new_n459_), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT68), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n460_), .A2(new_n462_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n453_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n464_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT68), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  AND3_X1   g269(.A1(new_n465_), .A2(new_n470_), .A3(KEYINPUT12), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n452_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G230gat), .A2(G233gat), .ZN(new_n473_));
  NOR3_X1   g272(.A1(new_n440_), .A2(new_n444_), .A3(new_n442_), .ZN(new_n474_));
  AOI22_X1  g273(.A1(new_n446_), .A2(new_n474_), .B1(new_n448_), .B2(new_n450_), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT66), .B1(new_n463_), .B2(new_n464_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT66), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n467_), .A2(new_n468_), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n475_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT12), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n481_), .B1(new_n475_), .B2(new_n479_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n472_), .A2(new_n473_), .A3(new_n480_), .A4(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n448_), .A2(new_n450_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n447_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(new_n479_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n483_), .B1(new_n473_), .B2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT5), .B(G176gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(new_n279_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G120gat), .B(G148gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n487_), .B(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT13), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G229gat), .A2(G233gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G29gat), .B(G36gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(G50gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT70), .B(G43gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(G50gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n496_), .B(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n498_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n499_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G15gat), .B(G22gat), .ZN(new_n505_));
  INV_X1    g304(.A(G1gat), .ZN(new_n506_));
  INV_X1    g305(.A(G8gat), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT14), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n505_), .A2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G1gat), .B(G8gat), .ZN(new_n510_));
  XOR2_X1   g309(.A(new_n509_), .B(new_n510_), .Z(new_n511_));
  NAND2_X1  g310(.A1(new_n504_), .A2(new_n511_), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n499_), .A2(new_n503_), .A3(KEYINPUT15), .ZN(new_n513_));
  AOI21_X1  g312(.A(KEYINPUT15), .B1(new_n499_), .B2(new_n503_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n495_), .B(new_n512_), .C1(new_n516_), .C2(new_n511_), .ZN(new_n517_));
  AOI21_X1  g316(.A(KEYINPUT78), .B1(new_n504_), .B2(new_n511_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n518_), .B1(new_n504_), .B2(new_n511_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n504_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n511_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(KEYINPUT78), .A3(new_n521_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n519_), .A2(G229gat), .A3(G233gat), .A4(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n517_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G113gat), .B(G141gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT79), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G169gat), .B(G197gat), .ZN(new_n527_));
  XOR2_X1   g326(.A(new_n526_), .B(new_n527_), .Z(new_n528_));
  NAND2_X1  g327(.A1(new_n524_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n528_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n517_), .A2(new_n523_), .A3(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n494_), .A2(new_n533_), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n404_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n452_), .A2(new_n515_), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT71), .B1(new_n485_), .B2(new_n520_), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G232gat), .A2(G233gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT34), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(KEYINPUT69), .B(KEYINPUT35), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT71), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n475_), .A2(new_n546_), .A3(new_n504_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n541_), .A2(new_n543_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n538_), .A2(new_n545_), .A3(new_n547_), .A4(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n536_), .A2(new_n547_), .A3(new_n537_), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n550_), .A2(KEYINPUT72), .A3(new_n544_), .ZN(new_n551_));
  AOI21_X1  g350(.A(KEYINPUT72), .B1(new_n550_), .B2(new_n544_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n549_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G190gat), .B(G218gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G134gat), .B(G162gat), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n554_), .B(new_n555_), .Z(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n557_), .A2(KEYINPUT36), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(KEYINPUT36), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n553_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n558_), .B(KEYINPUT73), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n549_), .B(new_n561_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G231gat), .A2(G233gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n511_), .B(new_n565_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n465_), .A2(new_n470_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n569_));
  XNOR2_X1  g368(.A(G127gat), .B(G155gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G183gat), .B(G211gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(KEYINPUT77), .B(KEYINPUT17), .Z(new_n574_));
  OR3_X1    g373(.A1(new_n568_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n566_), .B(new_n479_), .Z(new_n576_));
  XNOR2_X1  g375(.A(new_n573_), .B(KEYINPUT17), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n564_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n535_), .A2(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(G1gat), .B1(new_n581_), .B2(new_n249_), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n582_), .B(KEYINPUT101), .Z(new_n583_));
  INV_X1    g382(.A(KEYINPUT74), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n560_), .A2(new_n584_), .A3(new_n562_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT37), .ZN(new_n586_));
  INV_X1    g385(.A(new_n562_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n586_), .B1(new_n587_), .B2(KEYINPUT74), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT75), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n585_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n589_), .B1(new_n585_), .B2(new_n588_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n563_), .A2(KEYINPUT37), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n590_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n593_), .A2(new_n579_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n535_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n249_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(new_n506_), .A3(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT38), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n583_), .A2(new_n599_), .ZN(G1324gat));
  OAI21_X1  g399(.A(G8gat), .B1(new_n581_), .B2(new_n328_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT102), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n602_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n603_), .A2(KEYINPUT39), .A3(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n328_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n596_), .A2(new_n507_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT39), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n601_), .A2(new_n602_), .A3(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n605_), .A2(new_n607_), .A3(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g410(.A(new_n349_), .ZN(new_n612_));
  OAI21_X1  g411(.A(G15gat), .B1(new_n581_), .B2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT41), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n595_), .A2(G15gat), .A3(new_n612_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n614_), .A2(new_n615_), .ZN(G1326gat));
  XNOR2_X1  g415(.A(new_n385_), .B(KEYINPUT103), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(G22gat), .B1(new_n581_), .B2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT42), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n618_), .A2(G22gat), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n620_), .B1(new_n595_), .B2(new_n621_), .ZN(G1327gat));
  INV_X1    g421(.A(new_n579_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n563_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n535_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT105), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(G29gat), .B1(new_n627_), .B2(new_n597_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n404_), .A2(new_n593_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(KEYINPUT104), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT43), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n632_), .A2(KEYINPUT44), .A3(new_n579_), .A4(new_n534_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n630_), .A2(new_n631_), .ZN(new_n634_));
  AOI21_X1  g433(.A(KEYINPUT43), .B1(new_n629_), .B2(KEYINPUT104), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n579_), .B(new_n534_), .C1(new_n634_), .C2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT44), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n633_), .A2(new_n638_), .A3(G29gat), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n628_), .B1(new_n639_), .B2(new_n597_), .ZN(G1328gat));
  INV_X1    g439(.A(G36gat), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n328_), .B(KEYINPUT106), .Z(new_n642_));
  NAND3_X1  g441(.A1(new_n627_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(KEYINPUT45), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT45), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n627_), .A2(new_n645_), .A3(new_n641_), .A4(new_n642_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n633_), .A2(new_n638_), .A3(new_n606_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(G36gat), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT46), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n647_), .A2(new_n649_), .A3(KEYINPUT46), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1329gat));
  NAND2_X1  g453(.A1(new_n633_), .A2(new_n638_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n349_), .A2(G43gat), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n627_), .A2(new_n349_), .ZN(new_n657_));
  OAI22_X1  g456(.A1(new_n655_), .A2(new_n656_), .B1(new_n657_), .B2(G43gat), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g458(.A(G50gat), .B1(new_n655_), .B2(new_n385_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n617_), .A2(new_n500_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT107), .Z(new_n662_));
  NAND2_X1  g461(.A1(new_n627_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n660_), .A2(new_n663_), .ZN(G1331gat));
  AOI21_X1  g463(.A(new_n455_), .B1(new_n597_), .B2(KEYINPUT110), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n493_), .A2(new_n532_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n404_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(new_n580_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT109), .Z(new_n669_));
  AOI211_X1 g468(.A(new_n665_), .B(new_n669_), .C1(KEYINPUT110), .C2(new_n455_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n667_), .A2(new_n594_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT108), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(G57gat), .B1(new_n673_), .B2(new_n597_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n670_), .A2(new_n674_), .ZN(G1332gat));
  INV_X1    g474(.A(KEYINPUT48), .ZN(new_n676_));
  INV_X1    g475(.A(new_n642_), .ZN(new_n677_));
  OAI21_X1  g476(.A(G64gat), .B1(new_n669_), .B2(new_n677_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n678_), .A2(KEYINPUT111), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n678_), .A2(KEYINPUT111), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n676_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n678_), .A2(KEYINPUT111), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n678_), .A2(KEYINPUT111), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(KEYINPUT48), .A3(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n673_), .A2(new_n456_), .A3(new_n642_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n681_), .A2(new_n684_), .A3(new_n685_), .ZN(G1333gat));
  OAI21_X1  g485(.A(G71gat), .B1(new_n669_), .B2(new_n612_), .ZN(new_n687_));
  XOR2_X1   g486(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(new_n689_));
  OR2_X1    g488(.A1(new_n612_), .A2(G71gat), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n689_), .B1(new_n672_), .B2(new_n690_), .ZN(G1334gat));
  OAI21_X1  g490(.A(G78gat), .B1(new_n669_), .B2(new_n618_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT50), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n618_), .A2(G78gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n693_), .B1(new_n672_), .B2(new_n694_), .ZN(G1335gat));
  AND2_X1   g494(.A1(new_n667_), .A2(new_n624_), .ZN(new_n696_));
  AOI21_X1  g495(.A(G85gat), .B1(new_n696_), .B2(new_n597_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n632_), .A2(KEYINPUT113), .A3(new_n579_), .A4(new_n666_), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n579_), .B(new_n666_), .C1(new_n634_), .C2(new_n635_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT113), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n698_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n597_), .A2(G85gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n697_), .B1(new_n703_), .B2(new_n704_), .ZN(G1336gat));
  AOI21_X1  g504(.A(G92gat), .B1(new_n696_), .B2(new_n606_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n703_), .A2(G92gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n707_), .B2(new_n642_), .ZN(G1337gat));
  OAI21_X1  g507(.A(G99gat), .B1(new_n702_), .B2(new_n612_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n612_), .B1(new_n436_), .B2(new_n439_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n696_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT51), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT51), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n709_), .A2(new_n714_), .A3(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1338gat));
  AND3_X1   g515(.A1(new_n696_), .A2(new_n407_), .A3(new_n401_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G106gat), .B1(new_n699_), .B2(new_n385_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT52), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT52), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n720_), .B(G106gat), .C1(new_n699_), .C2(new_n385_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n717_), .B1(new_n719_), .B2(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n722_), .B(new_n724_), .ZN(G1339gat));
  NAND2_X1  g524(.A1(new_n585_), .A2(new_n588_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT75), .ZN(new_n727_));
  INV_X1    g526(.A(new_n592_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n585_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n727_), .A2(new_n728_), .A3(new_n729_), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n730_), .A2(new_n623_), .A3(new_n533_), .A4(new_n493_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT54), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT58), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n483_), .A2(KEYINPUT115), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT55), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n472_), .A2(new_n480_), .A3(new_n482_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n736_), .A2(G230gat), .A3(G233gat), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT55), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n483_), .A2(KEYINPUT115), .A3(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n735_), .A2(new_n737_), .A3(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(new_n491_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT56), .ZN(new_n742_));
  AOI21_X1  g541(.A(KEYINPUT118), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT118), .ZN(new_n744_));
  AOI211_X1 g543(.A(new_n744_), .B(KEYINPUT56), .C1(new_n740_), .C2(new_n491_), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n740_), .A2(KEYINPUT56), .A3(new_n491_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n743_), .A2(new_n745_), .A3(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n519_), .A2(new_n495_), .A3(new_n522_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n512_), .B1(new_n516_), .B2(new_n511_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n528_), .B(new_n748_), .C1(new_n749_), .C2(new_n495_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n531_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT116), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n487_), .A2(new_n491_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n733_), .B1(new_n747_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n743_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n740_), .A2(KEYINPUT56), .A3(new_n491_), .ZN(new_n757_));
  AOI21_X1  g556(.A(KEYINPUT56), .B1(new_n740_), .B2(new_n491_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT118), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n756_), .A2(new_n757_), .A3(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n754_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(KEYINPUT58), .A3(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n593_), .A2(new_n755_), .A3(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n753_), .A2(new_n532_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n765_), .B1(new_n746_), .B2(new_n758_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n752_), .A2(new_n492_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n564_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT117), .ZN(new_n769_));
  OAI21_X1  g568(.A(KEYINPUT57), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n741_), .A2(new_n742_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n764_), .B1(new_n771_), .B2(new_n757_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n752_), .A2(new_n492_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n563_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT57), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(KEYINPUT117), .A3(new_n775_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n763_), .A2(KEYINPUT119), .A3(new_n770_), .A4(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n579_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n770_), .A2(new_n776_), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT119), .B1(new_n779_), .B2(new_n763_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n732_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n384_), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n782_), .A2(new_n249_), .A3(new_n606_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(G113gat), .B1(new_n785_), .B2(new_n532_), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n731_), .B(KEYINPUT54), .Z(new_n787_));
  AOI21_X1  g586(.A(new_n623_), .B1(new_n779_), .B2(new_n763_), .ZN(new_n788_));
  OR2_X1    g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT59), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n790_), .A3(new_n783_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n784_), .A2(KEYINPUT59), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n532_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n786_), .B1(new_n795_), .B2(G113gat), .ZN(G1340gat));
  NAND2_X1  g595(.A1(new_n791_), .A2(new_n792_), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT120), .B1(new_n797_), .B2(new_n493_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT120), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n791_), .A2(new_n792_), .A3(new_n799_), .A4(new_n494_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n798_), .A2(G120gat), .A3(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(G120gat), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n802_), .B1(new_n493_), .B2(KEYINPUT60), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n785_), .B(new_n803_), .C1(KEYINPUT60), .C2(new_n802_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n801_), .A2(new_n804_), .ZN(G1341gat));
  AOI21_X1  g604(.A(G127gat), .B1(new_n785_), .B2(new_n623_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT121), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n807_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n623_), .A2(G127gat), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(KEYINPUT122), .ZN(new_n811_));
  AOI22_X1  g610(.A1(new_n808_), .A2(new_n809_), .B1(new_n793_), .B2(new_n811_), .ZN(G1342gat));
  AND3_X1   g611(.A1(new_n793_), .A2(G134gat), .A3(new_n593_), .ZN(new_n813_));
  AOI21_X1  g612(.A(G134gat), .B1(new_n785_), .B2(new_n564_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n813_), .A2(new_n814_), .ZN(G1343gat));
  INV_X1    g614(.A(new_n781_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n816_), .A2(new_n249_), .A3(new_n642_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n386_), .ZN(new_n818_));
  OR3_X1    g617(.A1(new_n818_), .A2(G141gat), .A3(new_n533_), .ZN(new_n819_));
  OAI21_X1  g618(.A(G141gat), .B1(new_n818_), .B2(new_n533_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(G1344gat));
  OR3_X1    g620(.A1(new_n818_), .A2(G148gat), .A3(new_n493_), .ZN(new_n822_));
  OAI21_X1  g621(.A(G148gat), .B1(new_n818_), .B2(new_n493_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(G1345gat));
  XNOR2_X1  g623(.A(KEYINPUT61), .B(G155gat), .ZN(new_n825_));
  INV_X1    g624(.A(new_n818_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(new_n623_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n825_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n818_), .A2(new_n579_), .A3(new_n828_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n827_), .A2(new_n829_), .ZN(G1346gat));
  INV_X1    g629(.A(G162gat), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n818_), .A2(new_n831_), .A3(new_n730_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n826_), .A2(new_n564_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n832_), .B1(new_n831_), .B2(new_n833_), .ZN(G1347gat));
  AND2_X1   g633(.A1(new_n789_), .A2(new_n618_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n642_), .A2(new_n249_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n836_), .A2(new_n612_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n835_), .A2(new_n532_), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(G169gat), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT62), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n835_), .A2(new_n837_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n843_), .A2(new_n532_), .A3(new_n251_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n838_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n841_), .A2(new_n844_), .A3(new_n845_), .ZN(G1348gat));
  NOR3_X1   g645(.A1(new_n816_), .A2(new_n782_), .A3(new_n836_), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n847_), .A2(G176gat), .A3(new_n494_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n789_), .A2(new_n494_), .A3(new_n618_), .A4(new_n837_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n252_), .ZN(new_n850_));
  OR2_X1    g649(.A1(new_n850_), .A2(KEYINPUT123), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(KEYINPUT123), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n848_), .B1(new_n851_), .B2(new_n852_), .ZN(G1349gat));
  AOI21_X1  g652(.A(new_n259_), .B1(new_n847_), .B2(new_n623_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n623_), .A2(new_n301_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n843_), .B2(new_n855_), .ZN(G1350gat));
  OAI21_X1  g655(.A(G190gat), .B1(new_n842_), .B2(new_n730_), .ZN(new_n857_));
  OR2_X1    g656(.A1(new_n842_), .A2(new_n300_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n563_), .ZN(G1351gat));
  NAND2_X1  g658(.A1(new_n386_), .A2(new_n249_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(KEYINPUT124), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(new_n677_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n781_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT125), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n781_), .A2(KEYINPUT125), .A3(new_n862_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n532_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(KEYINPUT126), .B(G197gat), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n868_), .B(new_n869_), .ZN(G1352gat));
  NAND2_X1  g669(.A1(new_n867_), .A2(new_n494_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G204gat), .ZN(G1353gat));
  XNOR2_X1  g671(.A(KEYINPUT63), .B(G211gat), .ZN(new_n873_));
  AND3_X1   g672(.A1(new_n781_), .A2(KEYINPUT125), .A3(new_n862_), .ZN(new_n874_));
  AOI21_X1  g673(.A(KEYINPUT125), .B1(new_n781_), .B2(new_n862_), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n623_), .B(new_n873_), .C1(new_n874_), .C2(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n579_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n876_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(KEYINPUT127), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT127), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n876_), .B(new_n881_), .C1(new_n877_), .C2(new_n878_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(G1354gat));
  AOI21_X1  g682(.A(G218gat), .B1(new_n867_), .B2(new_n564_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n730_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(G218gat), .B2(new_n885_), .ZN(G1355gat));
endmodule


