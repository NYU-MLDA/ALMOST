//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 0 0 1 0 1 1 1 1 0 0 1 1 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n836_, new_n838_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n847_, new_n849_, new_n850_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT34), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(KEYINPUT35), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT6), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT65), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT65), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT6), .ZN(new_n208_));
  AND2_X1   g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  AND3_X1   g008(.A1(new_n206_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n209_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND4_X1  g011(.A1(KEYINPUT64), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT9), .ZN(new_n215_));
  INV_X1    g014(.A(G85gat), .ZN(new_n216_));
  INV_X1    g015(.A(G92gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n215_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  XOR2_X1   g017(.A(G85gat), .B(G92gat), .Z(new_n219_));
  OAI211_X1 g018(.A(new_n214_), .B(new_n218_), .C1(new_n219_), .C2(new_n215_), .ZN(new_n220_));
  XOR2_X1   g019(.A(KEYINPUT10), .B(G99gat), .Z(new_n221_));
  INV_X1    g020(.A(G106gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n212_), .A2(new_n213_), .A3(new_n220_), .A4(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G99gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT7), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n225_), .B(new_n222_), .C1(new_n226_), .C2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n225_), .A2(new_n222_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n226_), .A2(new_n227_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n229_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n228_), .B(new_n232_), .C1(new_n210_), .C2(new_n211_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT8), .ZN(new_n234_));
  AND3_X1   g033(.A1(new_n233_), .A2(new_n234_), .A3(new_n219_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n234_), .B1(new_n233_), .B2(new_n219_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n224_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(KEYINPUT69), .B(G29gat), .Z(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(G36gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT69), .B(G29gat), .ZN(new_n241_));
  INV_X1    g040(.A(G36gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(new_n243_), .ZN(new_n244_));
  XOR2_X1   g043(.A(G43gat), .B(G50gat), .Z(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n240_), .A2(new_n245_), .A3(new_n243_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n204_), .B1(new_n238_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT15), .ZN(new_n252_));
  INV_X1    g051(.A(new_n248_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n245_), .B1(new_n240_), .B2(new_n243_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n252_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n247_), .A2(KEYINPUT15), .A3(new_n248_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n203_), .A2(KEYINPUT35), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT68), .ZN(new_n259_));
  AOI22_X1  g058(.A1(new_n257_), .A2(new_n237_), .B1(KEYINPUT71), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT72), .ZN(new_n261_));
  OR2_X1    g060(.A1(new_n259_), .A2(KEYINPUT71), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n251_), .A2(new_n260_), .A3(new_n261_), .A4(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n257_), .A2(new_n237_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n259_), .A2(KEYINPUT71), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n204_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n262_), .B(new_n267_), .C1(new_n237_), .C2(new_n249_), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT72), .B1(new_n266_), .B2(new_n268_), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n263_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT36), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G190gat), .B(G218gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(G134gat), .ZN(new_n273_));
  INV_X1    g072(.A(G162gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n276_), .B1(new_n257_), .B2(new_n237_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n257_), .A2(new_n237_), .A3(new_n276_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(new_n251_), .A3(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(new_n259_), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n270_), .A2(new_n271_), .A3(new_n275_), .A4(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n275_), .A2(new_n271_), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n275_), .A2(new_n271_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n263_), .A2(new_n269_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n259_), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n257_), .A2(new_n237_), .A3(new_n276_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n287_), .A2(new_n277_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n286_), .B1(new_n288_), .B2(new_n251_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n283_), .B(new_n284_), .C1(new_n285_), .C2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n282_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G227gat), .A2(G233gat), .ZN(new_n293_));
  XOR2_X1   g092(.A(new_n293_), .B(KEYINPUT30), .Z(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G15gat), .B(G43gat), .ZN(new_n296_));
  XOR2_X1   g095(.A(G71gat), .B(G99gat), .Z(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT25), .B(G183gat), .ZN(new_n299_));
  INV_X1    g098(.A(G190gat), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n299_), .B1(KEYINPUT26), .B2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT77), .B(G190gat), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n301_), .B1(KEYINPUT26), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G183gat), .A2(G190gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT23), .ZN(new_n305_));
  INV_X1    g104(.A(G169gat), .ZN(new_n306_));
  INV_X1    g105(.A(G176gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n308_), .A2(KEYINPUT24), .A3(new_n309_), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n305_), .B(new_n310_), .C1(KEYINPUT24), .C2(new_n308_), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n303_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(G183gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n302_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(new_n305_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT22), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT78), .B1(new_n316_), .B2(G169gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT22), .B(G169gat), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n307_), .B(new_n317_), .C1(new_n318_), .C2(KEYINPUT78), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n315_), .A2(new_n309_), .A3(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n298_), .B1(new_n312_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n312_), .A2(new_n320_), .A3(new_n298_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n296_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n323_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n296_), .ZN(new_n326_));
  NOR3_X1   g125(.A1(new_n325_), .A2(new_n326_), .A3(new_n321_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n295_), .B1(new_n324_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT80), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n326_), .B1(new_n325_), .B2(new_n321_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n322_), .A2(new_n296_), .A3(new_n323_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n330_), .A2(new_n331_), .A3(new_n294_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n328_), .A2(new_n329_), .A3(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G127gat), .B(G134gat), .ZN(new_n334_));
  INV_X1    g133(.A(G113gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(G120gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n333_), .B(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G211gat), .B(G218gat), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n343_), .A2(KEYINPUT21), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n343_), .A2(KEYINPUT21), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G197gat), .B(G204gat), .ZN(new_n346_));
  OR3_X1    g145(.A1(new_n344_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n343_), .A2(new_n346_), .A3(KEYINPUT21), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(G155gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n274_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(G141gat), .A2(G148gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT3), .ZN(new_n353_));
  NAND3_X1  g152(.A1(KEYINPUT81), .A2(G141gat), .A3(G148gat), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT83), .ZN(new_n355_));
  AOI21_X1  g154(.A(KEYINPUT2), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(KEYINPUT2), .ZN(new_n357_));
  AOI22_X1  g156(.A1(new_n357_), .A2(KEYINPUT81), .B1(G141gat), .B2(G148gat), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n353_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT84), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n351_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  AOI22_X1  g161(.A1(new_n359_), .A2(new_n360_), .B1(G155gat), .B2(G162gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G155gat), .A2(G162gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT1), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT82), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n367_), .B(new_n351_), .C1(KEYINPUT1), .C2(new_n364_), .ZN(new_n368_));
  AOI21_X1  g167(.A(KEYINPUT81), .B1(G141gat), .B2(G148gat), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n369_), .A2(new_n352_), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n370_), .A2(new_n354_), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n362_), .A2(new_n363_), .B1(new_n368_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT29), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n349_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  AND2_X1   g173(.A1(KEYINPUT86), .A2(G228gat), .ZN(new_n375_));
  NOR2_X1   g174(.A1(KEYINPUT86), .A2(G228gat), .ZN(new_n376_));
  OAI21_X1  g175(.A(G233gat), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n377_), .B(KEYINPUT87), .Z(new_n378_));
  INV_X1    g177(.A(KEYINPUT88), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G78gat), .B(G106gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n374_), .B(new_n383_), .C1(new_n379_), .C2(new_n378_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n349_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n368_), .A2(new_n371_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n358_), .A2(new_n356_), .ZN(new_n387_));
  XOR2_X1   g186(.A(new_n352_), .B(KEYINPUT3), .Z(new_n388_));
  NOR2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n364_), .B1(new_n389_), .B2(KEYINPUT84), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n386_), .B1(new_n390_), .B2(new_n361_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n385_), .B1(new_n391_), .B2(KEYINPUT29), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n378_), .A2(new_n379_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n382_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n384_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n396_), .B1(new_n391_), .B2(KEYINPUT29), .ZN(new_n397_));
  INV_X1    g196(.A(new_n396_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n372_), .A2(new_n373_), .A3(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G22gat), .B(G50gat), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n397_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n400_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n395_), .B1(new_n403_), .B2(KEYINPUT89), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT89), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n405_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT90), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n397_), .A2(new_n399_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n400_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n397_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT90), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n412_), .A2(new_n405_), .A3(new_n413_), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n404_), .A2(new_n407_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n403_), .A2(KEYINPUT89), .ZN(new_n416_));
  INV_X1    g215(.A(new_n395_), .ZN(new_n417_));
  AOI22_X1  g216(.A1(new_n407_), .A2(new_n414_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n342_), .B1(new_n415_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n416_), .A2(new_n417_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n413_), .B1(new_n412_), .B2(new_n405_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n406_), .A2(KEYINPUT90), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n420_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n333_), .B(new_n340_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n404_), .A2(new_n407_), .A3(new_n414_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n419_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT92), .ZN(new_n428_));
  INV_X1    g227(.A(new_n338_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n391_), .A2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n428_), .B1(new_n430_), .B2(KEYINPUT4), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n372_), .A2(new_n338_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n432_), .A2(new_n430_), .A3(KEYINPUT4), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT4), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n391_), .A2(KEYINPUT92), .A3(new_n429_), .A4(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n431_), .A2(new_n433_), .A3(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G225gat), .A2(G233gat), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n391_), .B(new_n338_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n440_), .A2(new_n438_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n439_), .A2(new_n442_), .ZN(new_n443_));
  XOR2_X1   g242(.A(G1gat), .B(G29gat), .Z(new_n444_));
  XNOR2_X1  g243(.A(G57gat), .B(G85gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n447_));
  XOR2_X1   g246(.A(new_n446_), .B(new_n447_), .Z(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n443_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT95), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n441_), .B1(new_n438_), .B2(new_n436_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n448_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n450_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n452_), .A2(KEYINPUT95), .A3(new_n448_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(KEYINPUT96), .A3(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(new_n455_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT96), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT27), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n385_), .A2(new_n320_), .A3(new_n312_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT26), .B(G190gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n299_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n311_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT91), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n313_), .A2(new_n300_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n305_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n309_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n470_), .B1(new_n318_), .B2(new_n307_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n466_), .A2(new_n472_), .ZN(new_n473_));
  OAI211_X1 g272(.A(KEYINPUT20), .B(new_n461_), .C1(new_n473_), .C2(new_n385_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G226gat), .A2(G233gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT19), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT18), .B(G64gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(new_n217_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G8gat), .B(G36gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n473_), .A2(new_n385_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n476_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT20), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n312_), .A2(new_n320_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n484_), .B1(new_n485_), .B2(new_n349_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n482_), .A2(new_n483_), .A3(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n477_), .A2(new_n481_), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n481_), .B1(new_n477_), .B2(new_n487_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n460_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n472_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n492_), .A2(new_n385_), .A3(new_n465_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n483_), .B1(new_n486_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n474_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n494_), .B1(new_n495_), .B2(new_n483_), .ZN(new_n496_));
  OAI211_X1 g295(.A(KEYINPUT27), .B(new_n488_), .C1(new_n496_), .C2(new_n481_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n491_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n427_), .A2(new_n456_), .A3(new_n459_), .A4(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n481_), .A2(KEYINPUT32), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n496_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n477_), .A2(new_n501_), .A3(new_n487_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n454_), .A2(new_n455_), .A3(new_n502_), .A4(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n489_), .A2(new_n490_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT33), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n450_), .A2(new_n506_), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n436_), .A2(new_n438_), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n440_), .B(KEYINPUT94), .Z(new_n509_));
  OAI211_X1 g308(.A(new_n448_), .B(new_n508_), .C1(new_n509_), .C2(new_n437_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n443_), .A2(KEYINPUT33), .A3(new_n449_), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n505_), .A2(new_n507_), .A3(new_n510_), .A4(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n504_), .A2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n415_), .A2(new_n418_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n514_), .A2(new_n342_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n292_), .B1(new_n500_), .B2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G15gat), .B(G22gat), .ZN(new_n518_));
  INV_X1    g317(.A(G1gat), .ZN(new_n519_));
  INV_X1    g318(.A(G8gat), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT14), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n518_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G1gat), .B(G8gat), .ZN(new_n523_));
  XOR2_X1   g322(.A(new_n522_), .B(new_n523_), .Z(new_n524_));
  XNOR2_X1  g323(.A(G57gat), .B(G64gat), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n525_), .A2(KEYINPUT11), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(KEYINPUT11), .ZN(new_n527_));
  XOR2_X1   g326(.A(G71gat), .B(G78gat), .Z(new_n528_));
  NAND3_X1  g327(.A1(new_n526_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  OR2_X1    g328(.A1(new_n527_), .A2(new_n528_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n524_), .B(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G231gat), .A2(G233gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT17), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G127gat), .B(G155gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G183gat), .B(G211gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  OR3_X1    g340(.A1(new_n535_), .A2(new_n536_), .A3(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(KEYINPUT17), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n535_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n531_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n237_), .A2(new_n547_), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n224_), .B(new_n531_), .C1(new_n235_), .C2(new_n236_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n548_), .A2(KEYINPUT12), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT12), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n237_), .A2(new_n551_), .A3(new_n547_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G230gat), .A2(G233gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n548_), .A2(new_n549_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n554_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n555_), .A2(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(G120gat), .B(G148gat), .Z(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G176gat), .B(G204gat), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n562_), .B(new_n563_), .Z(new_n564_));
  XNOR2_X1  g363(.A(new_n559_), .B(new_n564_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n565_), .A2(KEYINPUT13), .ZN(new_n566_));
  INV_X1    g365(.A(new_n524_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n257_), .A2(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n567_), .A2(new_n249_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G229gat), .A2(G233gat), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n568_), .A2(new_n570_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n571_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n250_), .A2(new_n524_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n573_), .B1(new_n574_), .B2(new_n569_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G113gat), .B(G141gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(new_n306_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(G197gat), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n572_), .A2(new_n575_), .A3(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT74), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT75), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT75), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n579_), .A2(new_n580_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n572_), .A2(new_n575_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n586_), .A2(new_n578_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n585_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n585_), .A2(new_n588_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n565_), .A2(KEYINPUT13), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n566_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n517_), .A2(new_n546_), .A3(new_n595_), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n596_), .A2(KEYINPUT97), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(KEYINPUT97), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n459_), .A2(new_n456_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(G1gat), .B1(new_n599_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n500_), .A2(new_n516_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT37), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n291_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n282_), .A2(new_n290_), .A3(KEYINPUT37), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n607_), .A2(new_n545_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT13), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n565_), .B(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT76), .ZN(new_n612_));
  INV_X1    g411(.A(new_n591_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n612_), .B1(new_n613_), .B2(new_n589_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n590_), .A2(new_n591_), .A3(KEYINPUT76), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n611_), .A2(new_n616_), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n603_), .A2(new_n608_), .A3(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n618_), .A2(new_n519_), .A3(new_n600_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(KEYINPUT98), .A2(KEYINPUT38), .ZN(new_n620_));
  AND2_X1   g419(.A1(KEYINPUT98), .A2(KEYINPUT38), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n619_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n619_), .A2(new_n620_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n602_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT99), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(G1324gat));
  NAND4_X1  g425(.A1(new_n517_), .A2(new_n546_), .A3(new_n498_), .A4(new_n595_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  AOI211_X1 g428(.A(new_n292_), .B(new_n594_), .C1(new_n500_), .C2(new_n516_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n630_), .A2(KEYINPUT100), .A3(new_n546_), .A4(new_n498_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n629_), .A2(new_n631_), .A3(G8gat), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT39), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT39), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n629_), .A2(new_n631_), .A3(new_n634_), .A4(G8gat), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n618_), .A2(new_n520_), .A3(new_n498_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT101), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n636_), .A2(new_n640_), .A3(new_n637_), .ZN(new_n641_));
  AOI21_X1  g440(.A(KEYINPUT40), .B1(new_n639_), .B2(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n640_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n637_), .ZN(new_n644_));
  AOI211_X1 g443(.A(KEYINPUT101), .B(new_n644_), .C1(new_n633_), .C2(new_n635_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT40), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n643_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n642_), .A2(new_n647_), .ZN(G1325gat));
  OAI21_X1  g447(.A(G15gat), .B1(new_n599_), .B2(new_n424_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT41), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(G15gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n618_), .A2(new_n652_), .A3(new_n342_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(G1326gat));
  INV_X1    g453(.A(G22gat), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n618_), .A2(new_n655_), .A3(new_n514_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n514_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n657_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n658_));
  OR3_X1    g457(.A1(new_n658_), .A2(KEYINPUT102), .A3(new_n655_), .ZN(new_n659_));
  OAI21_X1  g458(.A(KEYINPUT102), .B1(new_n658_), .B2(new_n655_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n659_), .A2(KEYINPUT42), .A3(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT42), .B1(new_n659_), .B2(new_n660_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n656_), .B1(new_n661_), .B2(new_n662_), .ZN(G1327gat));
  NAND3_X1  g462(.A1(new_n610_), .A2(new_n545_), .A3(new_n592_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT103), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT43), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(new_n603_), .B2(new_n607_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n607_), .ZN(new_n668_));
  AOI211_X1 g467(.A(KEYINPUT43), .B(new_n668_), .C1(new_n500_), .C2(new_n516_), .ZN(new_n669_));
  OAI211_X1 g468(.A(new_n665_), .B(KEYINPUT104), .C1(new_n667_), .C2(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(KEYINPUT44), .B1(new_n670_), .B2(KEYINPUT105), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n672_), .B1(KEYINPUT105), .B2(KEYINPUT44), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n667_), .A2(new_n669_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n674_), .B2(new_n665_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n671_), .A2(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G29gat), .B1(new_n676_), .B2(new_n601_), .ZN(new_n677_));
  AOI211_X1 g476(.A(new_n291_), .B(new_n546_), .C1(new_n500_), .C2(new_n516_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(new_n617_), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n601_), .A2(G29gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n677_), .B1(new_n679_), .B2(new_n680_), .ZN(G1328gat));
  NAND3_X1  g480(.A1(new_n678_), .A2(new_n242_), .A3(new_n617_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n498_), .B(KEYINPUT106), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  OR3_X1    g484(.A1(new_n682_), .A2(new_n683_), .A3(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n683_), .B1(new_n682_), .B2(new_n685_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n498_), .B1(new_n671_), .B2(new_n675_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(G36gat), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT108), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT46), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n690_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n691_), .A2(new_n692_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n690_), .A2(new_n694_), .A3(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n693_), .A2(new_n696_), .ZN(G1329gat));
  OAI21_X1  g496(.A(G43gat), .B1(new_n676_), .B2(new_n424_), .ZN(new_n698_));
  OR3_X1    g497(.A1(new_n679_), .A2(G43gat), .A3(new_n424_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT47), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n698_), .A2(KEYINPUT47), .A3(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1330gat));
  OAI21_X1  g503(.A(G50gat), .B1(new_n676_), .B2(new_n657_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n657_), .A2(G50gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(new_n679_), .B2(new_n706_), .ZN(G1331gat));
  NAND2_X1  g506(.A1(new_n611_), .A2(new_n608_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT109), .Z(new_n709_));
  INV_X1    g508(.A(new_n592_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n709_), .A2(new_n710_), .A3(new_n603_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(G57gat), .B1(new_n712_), .B2(new_n600_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n545_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n517_), .A2(new_n611_), .A3(new_n714_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n715_), .A2(new_n600_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n713_), .B1(G57gat), .B2(new_n716_), .ZN(G1332gat));
  INV_X1    g516(.A(G64gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n715_), .B2(new_n684_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT48), .Z(new_n720_));
  NAND3_X1  g519(.A1(new_n712_), .A2(new_n718_), .A3(new_n684_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1333gat));
  INV_X1    g521(.A(G71gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n723_), .B1(new_n715_), .B2(new_n342_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT49), .Z(new_n725_));
  NAND3_X1  g524(.A1(new_n712_), .A2(new_n723_), .A3(new_n342_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1334gat));
  INV_X1    g526(.A(G78gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n715_), .B2(new_n514_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT50), .Z(new_n730_));
  NAND3_X1  g529(.A1(new_n712_), .A2(new_n728_), .A3(new_n514_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1335gat));
  NOR2_X1   g531(.A1(new_n610_), .A2(new_n592_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n674_), .A2(new_n545_), .A3(new_n733_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT110), .Z(new_n735_));
  OAI21_X1  g534(.A(G85gat), .B1(new_n735_), .B2(new_n601_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n678_), .A2(new_n733_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n738_), .A2(new_n216_), .A3(new_n600_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n736_), .A2(new_n739_), .ZN(G1336gat));
  OAI21_X1  g539(.A(G92gat), .B1(new_n735_), .B2(new_n685_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n738_), .A2(new_n217_), .A3(new_n498_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1337gat));
  OAI21_X1  g542(.A(G99gat), .B1(new_n734_), .B2(new_n424_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n738_), .A2(new_n221_), .A3(new_n342_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g546(.A1(new_n738_), .A2(new_n222_), .A3(new_n514_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G106gat), .B1(new_n734_), .B2(new_n657_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n749_), .A2(KEYINPUT52), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n751_), .B(G106gat), .C1(new_n734_), .C2(new_n657_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n748_), .B1(new_n750_), .B2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT53), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT53), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n756_), .B(new_n748_), .C1(new_n750_), .C2(new_n753_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1339gat));
  NAND3_X1  g557(.A1(new_n714_), .A2(new_n668_), .A3(new_n610_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT54), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n759_), .B(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT111), .ZN(new_n762_));
  INV_X1    g561(.A(new_n564_), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT55), .B1(new_n553_), .B2(new_n554_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n765_));
  AOI211_X1 g564(.A(new_n765_), .B(new_n557_), .C1(new_n550_), .C2(new_n552_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n553_), .A2(new_n554_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n763_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n762_), .B1(new_n770_), .B2(KEYINPUT56), .ZN(new_n771_));
  INV_X1    g570(.A(new_n764_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n553_), .A2(KEYINPUT55), .A3(new_n554_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n772_), .A2(new_n769_), .A3(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(KEYINPUT56), .A3(new_n564_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT56), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n764_), .A2(new_n766_), .A3(new_n768_), .ZN(new_n777_));
  OAI211_X1 g576(.A(KEYINPUT111), .B(new_n776_), .C1(new_n777_), .C2(new_n763_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n771_), .A2(new_n775_), .A3(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n559_), .A2(new_n763_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(new_n592_), .A3(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n568_), .A2(new_n570_), .A3(new_n573_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n578_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n571_), .B1(new_n574_), .B2(new_n569_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n782_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n579_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n579_), .A2(new_n785_), .A3(KEYINPUT112), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n565_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n781_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n291_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT57), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n793_), .A2(KEYINPUT57), .A3(new_n291_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n780_), .A2(new_n790_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n776_), .B1(new_n777_), .B2(new_n763_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(new_n775_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n607_), .B1(new_n800_), .B2(KEYINPUT58), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT113), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(KEYINPUT58), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT113), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n607_), .B(new_n804_), .C1(new_n800_), .C2(KEYINPUT58), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n802_), .A2(new_n803_), .A3(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n796_), .A2(new_n797_), .A3(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n761_), .B1(new_n807_), .B2(new_n545_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n600_), .A2(new_n499_), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n808_), .A2(new_n419_), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(G113gat), .B1(new_n810_), .B2(new_n592_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n812_), .A2(KEYINPUT59), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n807_), .A2(new_n545_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n761_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n419_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n809_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n813_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(KEYINPUT114), .B(KEYINPUT59), .ZN(new_n819_));
  NOR4_X1   g618(.A1(new_n808_), .A2(new_n419_), .A3(new_n809_), .A4(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(KEYINPUT115), .B1(new_n818_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n819_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n816_), .A2(new_n817_), .A3(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n823_), .B(new_n824_), .C1(new_n810_), .C2(new_n813_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n335_), .B1(new_n821_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n616_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n811_), .B1(new_n826_), .B2(new_n827_), .ZN(G1340gat));
  OAI21_X1  g627(.A(new_n337_), .B1(new_n610_), .B2(KEYINPUT60), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n810_), .B(new_n829_), .C1(KEYINPUT60), .C2(new_n337_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n818_), .A2(new_n820_), .A3(new_n610_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n831_), .B2(new_n337_), .ZN(G1341gat));
  AOI21_X1  g631(.A(G127gat), .B1(new_n810_), .B2(new_n546_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n821_), .A2(new_n825_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n546_), .A2(G127gat), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(KEYINPUT116), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n833_), .B1(new_n834_), .B2(new_n836_), .ZN(G1342gat));
  AOI21_X1  g636(.A(G134gat), .B1(new_n810_), .B2(new_n292_), .ZN(new_n838_));
  XOR2_X1   g637(.A(KEYINPUT117), .B(G134gat), .Z(new_n839_));
  NOR2_X1   g638(.A1(new_n668_), .A2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n838_), .B1(new_n834_), .B2(new_n840_), .ZN(G1343gat));
  NOR2_X1   g640(.A1(new_n808_), .A2(new_n426_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n842_), .A2(new_n600_), .A3(new_n685_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n843_), .A2(new_n710_), .ZN(new_n844_));
  XOR2_X1   g643(.A(KEYINPUT118), .B(G141gat), .Z(new_n845_));
  XNOR2_X1  g644(.A(new_n844_), .B(new_n845_), .ZN(G1344gat));
  NOR2_X1   g645(.A1(new_n843_), .A2(new_n610_), .ZN(new_n847_));
  XOR2_X1   g646(.A(new_n847_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g647(.A1(new_n843_), .A2(new_n545_), .ZN(new_n849_));
  XOR2_X1   g648(.A(KEYINPUT61), .B(G155gat), .Z(new_n850_));
  XNOR2_X1  g649(.A(new_n849_), .B(new_n850_), .ZN(G1346gat));
  NOR3_X1   g650(.A1(new_n843_), .A2(new_n274_), .A3(new_n668_), .ZN(new_n852_));
  OR2_X1    g651(.A1(new_n843_), .A2(new_n291_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n274_), .B2(new_n853_), .ZN(G1347gat));
  INV_X1    g653(.A(KEYINPUT62), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n601_), .A2(new_n684_), .ZN(new_n856_));
  NOR4_X1   g655(.A1(new_n808_), .A2(new_n710_), .A3(new_n419_), .A4(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n855_), .B1(new_n857_), .B2(new_n306_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n856_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n816_), .A2(new_n592_), .A3(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n860_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n857_), .A2(new_n318_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n858_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT119), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n858_), .A2(new_n861_), .A3(new_n865_), .A4(new_n862_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n866_), .ZN(G1348gat));
  NOR3_X1   g666(.A1(new_n808_), .A2(new_n419_), .A3(new_n856_), .ZN(new_n868_));
  AOI21_X1  g667(.A(G176gat), .B1(new_n868_), .B2(new_n611_), .ZN(new_n869_));
  OR2_X1    g668(.A1(new_n869_), .A2(KEYINPUT120), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(KEYINPUT120), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n868_), .A2(G176gat), .A3(new_n611_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n873_));
  OR2_X1    g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n872_), .A2(new_n873_), .ZN(new_n875_));
  AOI22_X1  g674(.A1(new_n870_), .A2(new_n871_), .B1(new_n874_), .B2(new_n875_), .ZN(G1349gat));
  NAND2_X1  g675(.A1(new_n868_), .A2(new_n546_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n877_), .A2(new_n878_), .A3(new_n299_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n313_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(KEYINPUT122), .ZN(new_n881_));
  OR2_X1    g680(.A1(new_n877_), .A2(new_n299_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n879_), .B1(new_n881_), .B2(new_n882_), .ZN(G1350gat));
  NAND3_X1  g682(.A1(new_n868_), .A2(new_n292_), .A3(new_n462_), .ZN(new_n884_));
  AOI21_X1  g683(.A(KEYINPUT57), .B1(new_n793_), .B2(new_n291_), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n802_), .A2(new_n803_), .A3(new_n805_), .ZN(new_n886_));
  AOI211_X1 g685(.A(new_n795_), .B(new_n292_), .C1(new_n781_), .C2(new_n792_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n885_), .A2(new_n886_), .A3(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n815_), .B1(new_n888_), .B2(new_n546_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n419_), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n889_), .A2(new_n607_), .A3(new_n890_), .A4(new_n859_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n891_), .A2(new_n892_), .A3(G190gat), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n892_), .B1(new_n891_), .B2(G190gat), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n884_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(KEYINPUT124), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT124), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n897_), .B(new_n884_), .C1(new_n893_), .C2(new_n894_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n896_), .A2(new_n898_), .ZN(G1351gat));
  NOR3_X1   g698(.A1(new_n808_), .A2(new_n426_), .A3(new_n856_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n592_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n611_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n903_), .A2(G204gat), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(KEYINPUT126), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT126), .ZN(new_n906_));
  NOR3_X1   g705(.A1(new_n903_), .A2(new_n906_), .A3(G204gat), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT125), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n908_), .B1(new_n903_), .B2(G204gat), .ZN(new_n909_));
  AND3_X1   g708(.A1(new_n903_), .A2(new_n908_), .A3(G204gat), .ZN(new_n910_));
  OAI22_X1  g709(.A1(new_n905_), .A2(new_n907_), .B1(new_n909_), .B2(new_n910_), .ZN(G1353gat));
  NAND2_X1  g710(.A1(new_n842_), .A2(new_n859_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n912_), .A2(new_n545_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n913_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n914_));
  XOR2_X1   g713(.A(KEYINPUT63), .B(G211gat), .Z(new_n915_));
  AOI21_X1  g714(.A(new_n914_), .B1(new_n913_), .B2(new_n915_), .ZN(G1354gat));
  XOR2_X1   g715(.A(KEYINPUT127), .B(G218gat), .Z(new_n917_));
  NOR3_X1   g716(.A1(new_n912_), .A2(new_n668_), .A3(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n900_), .A2(new_n292_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n918_), .B1(new_n919_), .B2(new_n917_), .ZN(G1355gat));
endmodule


