//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n591_, new_n592_, new_n593_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n600_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n788_, new_n789_,
    new_n790_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n809_, new_n810_, new_n811_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n838_, new_n839_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_;
  XOR2_X1   g000(.A(G85gat), .B(G92gat), .Z(new_n202_));
  NOR2_X1   g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT7), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n202_), .B1(new_n205_), .B2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT8), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT10), .B(G99gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT64), .ZN(new_n212_));
  INV_X1    g011(.A(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n208_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n202_), .A2(KEYINPUT9), .ZN(new_n216_));
  INV_X1    g015(.A(G85gat), .ZN(new_n217_));
  INV_X1    g016(.A(G92gat), .ZN(new_n218_));
  OR3_X1    g017(.A1(new_n217_), .A2(new_n218_), .A3(KEYINPUT9), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .A4(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n210_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G29gat), .B(G36gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G43gat), .B(G50gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n223_), .B(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT35), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G232gat), .A2(G233gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT34), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  AOI22_X1  g028(.A1(new_n222_), .A2(new_n225_), .B1(new_n226_), .B2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n210_), .B(KEYINPUT66), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(new_n220_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n225_), .B(KEYINPUT15), .ZN(new_n233_));
  AND3_X1   g032(.A1(new_n232_), .A2(KEYINPUT68), .A3(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT68), .B1(new_n232_), .B2(new_n233_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n230_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n229_), .A2(new_n226_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  OAI221_X1 g037(.A(new_n230_), .B1(new_n226_), .B2(new_n229_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(G190gat), .B(G218gat), .Z(new_n241_));
  XNOR2_X1  g040(.A(G134gat), .B(G162gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT36), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n240_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT70), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT37), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT71), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT36), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n243_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT69), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n238_), .A2(new_n239_), .A3(new_n251_), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n245_), .A2(new_n248_), .A3(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n248_), .B1(new_n245_), .B2(new_n252_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n247_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n245_), .A2(new_n252_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT71), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT37), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n258_), .B1(new_n245_), .B2(KEYINPUT70), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n245_), .A2(new_n248_), .A3(new_n252_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n257_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G57gat), .B(G64gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT11), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(KEYINPUT11), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT65), .B(G71gat), .ZN(new_n265_));
  INV_X1    g064(.A(G78gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  MUX2_X1   g066(.A(new_n263_), .B(new_n264_), .S(new_n267_), .Z(new_n268_));
  NAND3_X1  g067(.A1(new_n232_), .A2(KEYINPUT12), .A3(new_n268_), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n221_), .A2(new_n268_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT12), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n221_), .A2(new_n268_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G230gat), .A2(G233gat), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n269_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n270_), .A2(new_n272_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n276_), .A2(G230gat), .A3(G233gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G120gat), .B(G148gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT5), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G176gat), .B(G204gat), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n280_), .B(new_n281_), .Z(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT67), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n278_), .B(new_n283_), .Z(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT13), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT72), .B(G15gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(G22gat), .ZN(new_n287_));
  INV_X1    g086(.A(G1gat), .ZN(new_n288_));
  INV_X1    g087(.A(G8gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT14), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G1gat), .B(G8gat), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n292_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G231gat), .A2(G233gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n297_), .B(new_n268_), .Z(new_n298_));
  XOR2_X1   g097(.A(G127gat), .B(G155gat), .Z(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(G183gat), .B(G211gat), .Z(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT17), .B1(new_n298_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT74), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n303_), .B1(new_n298_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  OAI211_X1 g106(.A(KEYINPUT17), .B(new_n303_), .C1(new_n298_), .C2(new_n305_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n255_), .A2(new_n261_), .A3(new_n285_), .A4(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT75), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n295_), .B(new_n225_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT76), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G229gat), .A2(G233gat), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n295_), .A2(new_n233_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT77), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n293_), .A2(new_n294_), .A3(new_n225_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(new_n320_), .A3(new_n314_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G113gat), .B(G141gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT78), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G169gat), .B(G197gat), .ZN(new_n324_));
  XOR2_X1   g123(.A(new_n323_), .B(new_n324_), .Z(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n316_), .A2(new_n321_), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT79), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT79), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n316_), .A2(new_n329_), .A3(new_n321_), .A4(new_n326_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n316_), .A2(new_n321_), .ZN(new_n331_));
  AOI22_X1  g130(.A1(new_n328_), .A2(new_n330_), .B1(new_n331_), .B2(new_n325_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(G169gat), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT23), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(G183gat), .A3(G190gat), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT80), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(G183gat), .ZN(new_n340_));
  INV_X1    g139(.A(G190gat), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT23), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n336_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n339_), .B1(new_n343_), .B2(KEYINPUT80), .ZN(new_n344_));
  NOR2_X1   g143(.A1(G183gat), .A2(G190gat), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n334_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT25), .B(G183gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT26), .B(G190gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  OR2_X1    g148(.A1(G169gat), .A2(G176gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G169gat), .A2(G176gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(KEYINPUT24), .A3(new_n351_), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n350_), .A2(KEYINPUT24), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n349_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n343_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n346_), .A2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G71gat), .B(G99gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(G43gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n356_), .B(new_n358_), .ZN(new_n359_));
  XOR2_X1   g158(.A(KEYINPUT81), .B(KEYINPUT31), .Z(new_n360_));
  XOR2_X1   g159(.A(new_n359_), .B(new_n360_), .Z(new_n361_));
  XOR2_X1   g160(.A(G127gat), .B(G134gat), .Z(new_n362_));
  XOR2_X1   g161(.A(G113gat), .B(G120gat), .Z(new_n363_));
  XOR2_X1   g162(.A(new_n362_), .B(new_n363_), .Z(new_n364_));
  NAND2_X1  g163(.A1(G227gat), .A2(G233gat), .ZN(new_n365_));
  INV_X1    g164(.A(G15gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT30), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n364_), .B(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n361_), .B(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT82), .ZN(new_n371_));
  INV_X1    g170(.A(new_n364_), .ZN(new_n372_));
  XOR2_X1   g171(.A(G155gat), .B(G162gat), .Z(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT3), .ZN(new_n375_));
  INV_X1    g174(.A(G141gat), .ZN(new_n376_));
  INV_X1    g175(.A(G148gat), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G141gat), .A2(G148gat), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT83), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n379_), .B1(new_n380_), .B2(KEYINPUT2), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n380_), .A2(KEYINPUT2), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n374_), .B(new_n378_), .C1(new_n381_), .C2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT84), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n373_), .B1(new_n383_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT85), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT85), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n389_), .B(new_n373_), .C1(new_n383_), .C2(new_n386_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT1), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n373_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n376_), .A2(new_n377_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n393_), .A2(new_n379_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n392_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n388_), .A2(new_n390_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT94), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n372_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  AOI22_X1  g198(.A1(new_n387_), .A2(KEYINPUT85), .B1(new_n392_), .B2(new_n395_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n400_), .A2(KEYINPUT94), .A3(new_n390_), .A4(new_n364_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G225gat), .A2(G233gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n372_), .A2(KEYINPUT4), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n402_), .A2(KEYINPUT4), .B1(new_n397_), .B2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n405_), .B1(new_n407_), .B2(new_n404_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G1gat), .B(G29gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(G85gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT0), .B(G57gat), .ZN(new_n411_));
  XOR2_X1   g210(.A(new_n410_), .B(new_n411_), .Z(new_n412_));
  NAND2_X1  g211(.A1(new_n408_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n412_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n405_), .B(new_n414_), .C1(new_n407_), .C2(new_n404_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G8gat), .B(G36gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT18), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G64gat), .B(G92gat), .ZN(new_n419_));
  XOR2_X1   g218(.A(new_n418_), .B(new_n419_), .Z(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT32), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G226gat), .A2(G233gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT19), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT87), .ZN(new_n425_));
  INV_X1    g224(.A(G197gat), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n425_), .B1(new_n426_), .B2(G204gat), .ZN(new_n427_));
  INV_X1    g226(.A(G204gat), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n428_), .A2(KEYINPUT87), .A3(G197gat), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT21), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n426_), .A2(G204gat), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n427_), .A2(new_n429_), .A3(new_n430_), .A4(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n426_), .A2(G204gat), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n428_), .A2(G197gat), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT21), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(G218gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(G211gat), .ZN(new_n437_));
  INV_X1    g236(.A(G211gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(G218gat), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n437_), .A2(new_n439_), .A3(KEYINPUT88), .ZN(new_n440_));
  AOI21_X1  g239(.A(KEYINPUT88), .B1(new_n437_), .B2(new_n439_), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n432_), .B(new_n435_), .C1(new_n440_), .C2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT88), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n438_), .A2(G218gat), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n436_), .A2(G211gat), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n443_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n427_), .A2(new_n431_), .A3(new_n429_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n437_), .A2(new_n439_), .A3(KEYINPUT88), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n446_), .A2(new_n447_), .A3(KEYINPUT21), .A4(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT89), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n449_), .A2(new_n450_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n442_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT90), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n442_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n440_), .A2(new_n441_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n457_), .A2(KEYINPUT89), .A3(KEYINPUT21), .A4(new_n447_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n449_), .A2(new_n450_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n456_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT90), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n455_), .A2(new_n461_), .A3(new_n356_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT20), .ZN(new_n463_));
  INV_X1    g262(.A(new_n344_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n343_), .B1(G183gat), .B2(G190gat), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n464_), .A2(new_n354_), .B1(new_n334_), .B2(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n463_), .B1(new_n460_), .B2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n424_), .B1(new_n462_), .B2(new_n467_), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n468_), .A2(KEYINPUT97), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT20), .B1(new_n460_), .B2(new_n466_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  AOI211_X1 g270(.A(new_n454_), .B(new_n456_), .C1(new_n459_), .C2(new_n458_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n458_), .A2(new_n459_), .ZN(new_n473_));
  AOI21_X1  g272(.A(KEYINPUT90), .B1(new_n473_), .B2(new_n442_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  OAI211_X1 g274(.A(new_n424_), .B(new_n471_), .C1(new_n475_), .C2(new_n356_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n476_), .B1(new_n468_), .B2(KEYINPUT97), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n469_), .A2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n416_), .B1(new_n421_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT93), .ZN(new_n480_));
  INV_X1    g279(.A(new_n356_), .ZN(new_n481_));
  NOR3_X1   g280(.A1(new_n472_), .A2(new_n474_), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n467_), .A2(new_n424_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n480_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n356_), .B1(new_n455_), .B2(new_n461_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n423_), .B1(new_n485_), .B2(new_n470_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n462_), .A2(KEYINPUT93), .A3(new_n424_), .A4(new_n467_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n484_), .A2(new_n486_), .A3(new_n421_), .A4(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT96), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT33), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n413_), .A2(KEYINPUT95), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT95), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n408_), .B(new_n412_), .C1(new_n492_), .C2(KEYINPUT33), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n407_), .A2(new_n404_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n495_), .B(new_n414_), .C1(new_n404_), .C2(new_n403_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n484_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n420_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n484_), .A2(new_n486_), .A3(new_n420_), .A4(new_n487_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n496_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  OAI22_X1  g300(.A1(new_n479_), .A2(new_n489_), .B1(new_n494_), .B2(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(G22gat), .B(G50gat), .Z(new_n503_));
  INV_X1    g302(.A(KEYINPUT29), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n388_), .A2(new_n504_), .A3(new_n390_), .A4(new_n396_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT28), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT86), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT28), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n400_), .A2(new_n508_), .A3(new_n504_), .A4(new_n390_), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n506_), .A2(new_n507_), .A3(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n507_), .B1(new_n506_), .B2(new_n509_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n503_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n506_), .A2(new_n509_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT86), .ZN(new_n514_));
  INV_X1    g313(.A(new_n503_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n506_), .A2(new_n507_), .A3(new_n509_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n514_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  AND2_X1   g316(.A1(new_n512_), .A2(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n504_), .B1(new_n400_), .B2(new_n390_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G228gat), .A2(G233gat), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n475_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n397_), .A2(KEYINPUT29), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(new_n453_), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT91), .B1(new_n525_), .B2(new_n521_), .ZN(new_n526_));
  OAI211_X1 g325(.A(KEYINPUT91), .B(new_n521_), .C1(new_n519_), .C2(new_n460_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n523_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G78gat), .B(G106gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT92), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT91), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n460_), .B1(new_n397_), .B2(KEYINPUT29), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n534_), .B1(new_n535_), .B2(new_n520_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(new_n527_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n537_), .A2(new_n523_), .A3(new_n531_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n518_), .A2(new_n533_), .A3(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n512_), .A2(new_n517_), .ZN(new_n540_));
  AOI221_X4 g339(.A(new_n532_), .B1(new_n475_), .B2(new_n522_), .C1(new_n536_), .C2(new_n527_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n531_), .B1(new_n537_), .B2(new_n523_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n540_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n539_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n502_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT27), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n499_), .A2(new_n500_), .ZN(new_n548_));
  AND2_X1   g347(.A1(new_n500_), .A2(KEYINPUT27), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n498_), .B1(new_n469_), .B2(new_n477_), .ZN(new_n550_));
  AOI22_X1  g349(.A1(new_n547_), .A2(new_n548_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n416_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(new_n544_), .A3(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n371_), .B1(new_n546_), .B2(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n370_), .A2(new_n416_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n549_), .A2(new_n550_), .ZN(new_n556_));
  AOI21_X1  g355(.A(KEYINPUT27), .B1(new_n499_), .B2(new_n500_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT98), .ZN(new_n558_));
  NOR4_X1   g357(.A1(new_n556_), .A2(new_n544_), .A3(new_n557_), .A4(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(KEYINPUT98), .B1(new_n551_), .B2(new_n545_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n555_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT99), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n548_), .A2(new_n547_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n549_), .A2(new_n550_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n558_), .B1(new_n565_), .B2(new_n544_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n551_), .A2(new_n545_), .A3(KEYINPUT98), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT99), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(new_n569_), .A3(new_n555_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n554_), .B1(new_n562_), .B2(new_n570_), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n311_), .A2(new_n332_), .A3(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n572_), .A2(new_n288_), .A3(new_n416_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT38), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n332_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n285_), .A2(new_n576_), .A3(new_n309_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n577_), .A2(KEYINPUT100), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n577_), .A2(KEYINPUT100), .ZN(new_n579_));
  INV_X1    g378(.A(new_n256_), .ZN(new_n580_));
  NOR4_X1   g379(.A1(new_n578_), .A2(new_n579_), .A3(new_n571_), .A4(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n288_), .B1(new_n581_), .B2(new_n416_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n575_), .A2(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n583_), .B1(new_n574_), .B2(new_n573_), .ZN(G1324gat));
  AOI21_X1  g383(.A(new_n289_), .B1(new_n581_), .B2(new_n565_), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n585_), .B(KEYINPUT39), .Z(new_n586_));
  NAND3_X1  g385(.A1(new_n572_), .A2(new_n289_), .A3(new_n565_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT40), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(G1325gat));
  AOI21_X1  g389(.A(new_n366_), .B1(new_n581_), .B2(new_n371_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT41), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n572_), .A2(new_n366_), .A3(new_n371_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(G1326gat));
  INV_X1    g393(.A(G22gat), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n595_), .B1(new_n581_), .B2(new_n544_), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n596_), .B(KEYINPUT42), .Z(new_n597_));
  NAND3_X1  g396(.A1(new_n572_), .A2(new_n595_), .A3(new_n544_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT101), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(G1327gat));
  INV_X1    g400(.A(new_n285_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n309_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n580_), .A2(new_n603_), .ZN(new_n604_));
  NOR4_X1   g403(.A1(new_n571_), .A2(new_n332_), .A3(new_n602_), .A4(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(G29gat), .B1(new_n605_), .B2(new_n416_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n255_), .A2(new_n261_), .ZN(new_n607_));
  OAI21_X1  g406(.A(KEYINPUT43), .B1(new_n571_), .B2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n546_), .A2(new_n553_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n371_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n569_), .B1(new_n568_), .B2(new_n555_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n555_), .ZN(new_n613_));
  AOI211_X1 g412(.A(KEYINPUT99), .B(new_n613_), .C1(new_n566_), .C2(new_n567_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n611_), .B1(new_n612_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT43), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n255_), .A2(new_n261_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n615_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n608_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n285_), .A2(new_n576_), .A3(new_n603_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(KEYINPUT44), .B1(new_n619_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT44), .ZN(new_n623_));
  AOI211_X1 g422(.A(new_n623_), .B(new_n620_), .C1(new_n608_), .C2(new_n618_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n416_), .A2(G29gat), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n606_), .B1(new_n625_), .B2(new_n626_), .ZN(G1328gat));
  INV_X1    g426(.A(KEYINPUT103), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n571_), .A2(new_n607_), .A3(KEYINPUT43), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n616_), .B1(new_n615_), .B2(new_n617_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n621_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(new_n623_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n619_), .A2(KEYINPUT44), .A3(new_n621_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n632_), .A2(new_n565_), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT102), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n634_), .A2(new_n635_), .A3(G36gat), .ZN(new_n636_));
  INV_X1    g435(.A(G36gat), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n605_), .A2(new_n637_), .A3(new_n565_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT45), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n636_), .A2(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n635_), .B1(new_n634_), .B2(G36gat), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n628_), .B(KEYINPUT46), .C1(new_n640_), .C2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n622_), .A2(new_n624_), .A3(new_n551_), .ZN(new_n644_));
  OAI21_X1  g443(.A(KEYINPUT102), .B1(new_n644_), .B2(new_n637_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n645_), .A2(new_n636_), .A3(new_n639_), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT46), .B1(new_n646_), .B2(new_n628_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n643_), .A2(new_n647_), .ZN(G1329gat));
  AOI21_X1  g447(.A(G43gat), .B1(new_n605_), .B2(new_n371_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n370_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n650_), .A2(G43gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n649_), .B1(new_n625_), .B2(new_n651_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g452(.A(G50gat), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n605_), .A2(new_n654_), .A3(new_n544_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n625_), .A2(KEYINPUT104), .A3(new_n544_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(G50gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT104), .B1(new_n625_), .B2(new_n544_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n655_), .B1(new_n657_), .B2(new_n658_), .ZN(G1331gat));
  NAND3_X1  g458(.A1(new_n602_), .A2(new_n332_), .A3(new_n309_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n571_), .A2(new_n660_), .A3(new_n580_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n661_), .A2(G57gat), .A3(new_n416_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n662_), .A2(KEYINPUT105), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n571_), .A2(new_n576_), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n617_), .A2(new_n285_), .A3(new_n603_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(G57gat), .B1(new_n667_), .B2(new_n416_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n662_), .A2(KEYINPUT105), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n663_), .A2(new_n668_), .A3(new_n669_), .ZN(G1332gat));
  NAND2_X1  g469(.A1(new_n661_), .A2(new_n565_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(G64gat), .ZN(new_n672_));
  XNOR2_X1  g471(.A(KEYINPUT106), .B(KEYINPUT48), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n672_), .B(new_n673_), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n551_), .A2(G64gat), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n674_), .B1(new_n666_), .B2(new_n675_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT107), .Z(G1333gat));
  INV_X1    g476(.A(G71gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n678_), .B1(new_n661_), .B2(new_n371_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT49), .Z(new_n680_));
  NAND3_X1  g479(.A1(new_n667_), .A2(new_n678_), .A3(new_n371_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1334gat));
  NAND3_X1  g481(.A1(new_n667_), .A2(new_n266_), .A3(new_n544_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n661_), .A2(new_n544_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(G78gat), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT109), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT109), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n684_), .A2(new_n687_), .A3(G78gat), .ZN(new_n688_));
  XNOR2_X1  g487(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n686_), .A2(new_n688_), .A3(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n686_), .B2(new_n688_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n683_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT110), .ZN(G1335gat));
  NOR4_X1   g492(.A1(new_n571_), .A2(new_n576_), .A3(new_n285_), .A4(new_n604_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT111), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n695_), .A2(new_n217_), .A3(new_n416_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n602_), .A2(new_n332_), .A3(new_n603_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT112), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n619_), .A2(new_n698_), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n699_), .A2(KEYINPUT113), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(KEYINPUT113), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n552_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n696_), .B1(new_n702_), .B2(new_n217_), .ZN(G1336gat));
  NAND3_X1  g502(.A1(new_n695_), .A2(new_n218_), .A3(new_n565_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n551_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n704_), .B1(new_n705_), .B2(new_n218_), .ZN(G1337gat));
  NAND3_X1  g505(.A1(new_n695_), .A2(new_n650_), .A3(new_n212_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n610_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n708_));
  INV_X1    g507(.A(G99gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n707_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g510(.A1(new_n619_), .A2(new_n698_), .A3(new_n544_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT114), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(G106gat), .B1(new_n712_), .B2(KEYINPUT114), .ZN(new_n715_));
  OAI21_X1  g514(.A(KEYINPUT52), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n712_), .A2(KEYINPUT114), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT52), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n717_), .A2(new_n718_), .A3(G106gat), .A4(new_n713_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n545_), .A2(G106gat), .ZN(new_n720_));
  AOI22_X1  g519(.A1(new_n716_), .A2(new_n719_), .B1(new_n695_), .B2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n721_), .B(new_n723_), .ZN(G1339gat));
  OR3_X1    g523(.A1(new_n310_), .A2(KEYINPUT54), .A3(new_n576_), .ZN(new_n725_));
  OAI21_X1  g524(.A(KEYINPUT54), .B1(new_n310_), .B2(new_n576_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n282_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n274_), .B1(new_n269_), .B2(new_n273_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT55), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n275_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n269_), .A2(new_n273_), .A3(KEYINPUT55), .A4(new_n274_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT56), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n275_), .A2(new_n277_), .A3(new_n728_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n737_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n736_), .A2(new_n332_), .A3(new_n738_), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n319_), .A2(new_n320_), .A3(new_n315_), .ZN(new_n740_));
  AOI211_X1 g539(.A(new_n326_), .B(new_n740_), .C1(new_n313_), .C2(new_n314_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n742_), .A2(new_n284_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n256_), .B1(new_n739_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT57), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n736_), .A2(new_n738_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n747_), .A2(KEYINPUT58), .A3(new_n742_), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n733_), .A2(new_n734_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n749_), .A2(new_n742_), .A3(new_n735_), .A4(new_n737_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT58), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n617_), .A2(new_n748_), .A3(new_n752_), .ZN(new_n753_));
  OAI211_X1 g552(.A(KEYINPUT57), .B(new_n256_), .C1(new_n739_), .C2(new_n743_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n746_), .A2(new_n753_), .A3(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n603_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n727_), .A2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT59), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n568_), .A2(new_n416_), .A3(new_n650_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n757_), .A2(new_n758_), .A3(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT116), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n309_), .B1(new_n755_), .B2(new_n762_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n746_), .A2(new_n753_), .A3(KEYINPUT116), .A4(new_n754_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n759_), .B1(new_n765_), .B2(new_n727_), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n576_), .B(new_n761_), .C1(new_n766_), .C2(new_n758_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(G113gat), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT117), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n766_), .A2(new_n769_), .ZN(new_n770_));
  AOI22_X1  g569(.A1(new_n763_), .A2(new_n764_), .B1(new_n726_), .B2(new_n725_), .ZN(new_n771_));
  OAI21_X1  g570(.A(KEYINPUT117), .B1(new_n771_), .B2(new_n759_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n332_), .A2(G113gat), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n770_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n768_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT118), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n768_), .A2(KEYINPUT118), .A3(new_n774_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(G1340gat));
  AND2_X1   g578(.A1(new_n770_), .A2(new_n772_), .ZN(new_n780_));
  INV_X1    g579(.A(G120gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n781_), .B1(new_n285_), .B2(KEYINPUT60), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n780_), .B(new_n782_), .C1(KEYINPUT60), .C2(new_n781_), .ZN(new_n783_));
  OAI21_X1  g582(.A(KEYINPUT59), .B1(new_n771_), .B2(new_n759_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n761_), .ZN(new_n785_));
  OAI21_X1  g584(.A(G120gat), .B1(new_n785_), .B2(new_n285_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n783_), .A2(new_n786_), .ZN(G1341gat));
  INV_X1    g586(.A(G127gat), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n780_), .A2(new_n788_), .A3(new_n309_), .ZN(new_n789_));
  OAI21_X1  g588(.A(G127gat), .B1(new_n785_), .B2(new_n603_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(G1342gat));
  NAND2_X1  g590(.A1(new_n780_), .A2(new_n580_), .ZN(new_n792_));
  INV_X1    g591(.A(G134gat), .ZN(new_n793_));
  INV_X1    g592(.A(new_n785_), .ZN(new_n794_));
  XOR2_X1   g593(.A(KEYINPUT119), .B(G134gat), .Z(new_n795_));
  NAND2_X1  g594(.A1(new_n617_), .A2(new_n795_), .ZN(new_n796_));
  XOR2_X1   g595(.A(new_n796_), .B(KEYINPUT120), .Z(new_n797_));
  AOI22_X1  g596(.A1(new_n792_), .A2(new_n793_), .B1(new_n794_), .B2(new_n797_), .ZN(G1343gat));
  NAND3_X1  g597(.A1(new_n610_), .A2(new_n544_), .A3(new_n416_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n771_), .A2(new_n565_), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n576_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n602_), .ZN(new_n803_));
  XOR2_X1   g602(.A(KEYINPUT121), .B(G148gat), .Z(new_n804_));
  XNOR2_X1  g603(.A(new_n803_), .B(new_n804_), .ZN(G1345gat));
  NAND2_X1  g604(.A1(new_n800_), .A2(new_n309_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(KEYINPUT61), .B(G155gat), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n806_), .B(new_n807_), .ZN(G1346gat));
  AOI21_X1  g607(.A(G162gat), .B1(new_n800_), .B2(new_n580_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n617_), .A2(G162gat), .ZN(new_n810_));
  XOR2_X1   g609(.A(new_n810_), .B(KEYINPUT122), .Z(new_n811_));
  AOI21_X1  g610(.A(new_n809_), .B1(new_n800_), .B2(new_n811_), .ZN(G1347gat));
  AOI21_X1  g611(.A(new_n544_), .B1(new_n727_), .B2(new_n756_), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n610_), .A2(new_n416_), .A3(new_n551_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n576_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n817_));
  INV_X1    g616(.A(G169gat), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n818_), .B1(KEYINPUT123), .B2(KEYINPUT62), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n816_), .A2(new_n817_), .A3(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n817_), .B1(new_n816_), .B2(new_n819_), .ZN(new_n821_));
  XOR2_X1   g620(.A(KEYINPUT22), .B(G169gat), .Z(new_n822_));
  OAI22_X1  g621(.A1(new_n820_), .A2(new_n821_), .B1(new_n816_), .B2(new_n822_), .ZN(G1348gat));
  AOI21_X1  g622(.A(G176gat), .B1(new_n815_), .B2(new_n602_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n771_), .A2(new_n544_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n602_), .A2(G176gat), .A3(new_n814_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n824_), .B1(new_n825_), .B2(new_n827_), .ZN(G1349gat));
  INV_X1    g627(.A(new_n347_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n814_), .A2(new_n309_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n813_), .A2(new_n829_), .A3(new_n830_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n825_), .A2(new_n830_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(G183gat), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT124), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  OAI211_X1 g634(.A(KEYINPUT124), .B(new_n831_), .C1(new_n832_), .C2(G183gat), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(G1350gat));
  NAND3_X1  g636(.A1(new_n815_), .A2(new_n348_), .A3(new_n580_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n815_), .A2(new_n617_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n839_), .B2(new_n341_), .ZN(G1351gat));
  NAND2_X1  g639(.A1(new_n765_), .A2(new_n727_), .ZN(new_n841_));
  NOR4_X1   g640(.A1(new_n371_), .A2(new_n545_), .A3(new_n416_), .A4(new_n551_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT125), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n841_), .A2(KEYINPUT125), .A3(new_n842_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(KEYINPUT126), .B(G197gat), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n847_), .A2(new_n576_), .A3(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n848_), .B1(new_n847_), .B2(new_n576_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1352gat));
  AOI21_X1  g650(.A(new_n285_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(new_n428_), .ZN(G1353gat));
  XNOR2_X1  g652(.A(KEYINPUT63), .B(G211gat), .ZN(new_n854_));
  AOI211_X1 g653(.A(new_n603_), .B(new_n854_), .C1(new_n845_), .C2(new_n846_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n847_), .A2(new_n309_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n855_), .B1(new_n856_), .B2(new_n857_), .ZN(G1354gat));
  NAND2_X1  g657(.A1(new_n847_), .A2(new_n580_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(KEYINPUT127), .B(G218gat), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n607_), .A2(new_n860_), .ZN(new_n861_));
  AOI22_X1  g660(.A1(new_n859_), .A2(new_n860_), .B1(new_n847_), .B2(new_n861_), .ZN(G1355gat));
endmodule


