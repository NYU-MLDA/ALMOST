//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n615_, new_n616_, new_n617_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n877_, new_n879_, new_n880_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_;
  XOR2_X1   g000(.A(KEYINPUT81), .B(KEYINPUT28), .Z(new_n202_));
  INV_X1    g001(.A(KEYINPUT3), .ZN(new_n203_));
  INV_X1    g002(.A(G141gat), .ZN(new_n204_));
  INV_X1    g003(.A(G148gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT2), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n210_));
  AND3_X1   g009(.A1(new_n206_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT79), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G155gat), .ZN(new_n216_));
  INV_X1    g015(.A(G162gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n215_), .A2(new_n219_), .A3(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n204_), .A2(new_n205_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(new_n207_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n219_), .A2(KEYINPUT1), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT1), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n220_), .B1(new_n218_), .B2(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n224_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n222_), .A2(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT80), .B1(new_n230_), .B2(KEYINPUT29), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  NOR3_X1   g031(.A1(new_n230_), .A2(KEYINPUT80), .A3(KEYINPUT29), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n202_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n233_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n202_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(new_n231_), .A3(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n234_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G228gat), .A2(G233gat), .ZN(new_n239_));
  INV_X1    g038(.A(G78gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(G106gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n238_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n243_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n234_), .A2(new_n237_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G211gat), .B(G218gat), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT21), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT83), .ZN(new_n251_));
  INV_X1    g050(.A(G204gat), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n251_), .B1(new_n252_), .B2(G197gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(G197gat), .ZN(new_n254_));
  INV_X1    g053(.A(G197gat), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(KEYINPUT83), .A3(G204gat), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n253_), .A2(new_n254_), .A3(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n250_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n255_), .A2(G204gat), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n249_), .B1(new_n254_), .B2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT82), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n248_), .B1(new_n257_), .B2(KEYINPUT21), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n258_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n264_), .B1(KEYINPUT29), .B2(new_n230_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G22gat), .B(G50gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n247_), .A2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n244_), .A2(new_n267_), .A3(new_n246_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(G8gat), .B(G36gat), .Z(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT87), .B(KEYINPUT18), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G64gat), .B(G92gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT25), .B(G183gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT26), .B(G190gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(G169gat), .ZN(new_n281_));
  INV_X1    g080(.A(G176gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G169gat), .A2(G176gat), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n283_), .A2(KEYINPUT24), .A3(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n280_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT23), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n287_), .A2(G183gat), .A3(G190gat), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT78), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(G183gat), .ZN(new_n291_));
  INV_X1    g090(.A(G190gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT23), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(new_n289_), .A3(new_n288_), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n283_), .A2(KEYINPUT24), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n290_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT85), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT85), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n290_), .A2(new_n294_), .A3(new_n295_), .A4(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n286_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT86), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n293_), .A2(new_n288_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(G183gat), .A2(G190gat), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n301_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n293_), .A2(new_n288_), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n305_), .B(KEYINPUT86), .C1(G183gat), .C2(G190gat), .ZN(new_n306_));
  INV_X1    g105(.A(new_n284_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT22), .B(G169gat), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n307_), .B1(new_n308_), .B2(new_n282_), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n304_), .A2(new_n306_), .A3(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n263_), .B1(new_n300_), .B2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n295_), .A2(new_n305_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n312_), .B1(new_n286_), .B2(KEYINPUT77), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT77), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n280_), .A2(new_n314_), .A3(new_n285_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n290_), .A2(new_n294_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n309_), .B1(new_n317_), .B2(new_n303_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n311_), .B(KEYINPUT20), .C1(new_n263_), .C2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G226gat), .A2(G233gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n320_), .A2(new_n324_), .ZN(new_n325_));
  OR3_X1    g124(.A1(new_n300_), .A2(new_n263_), .A3(new_n310_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT20), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n327_), .B1(new_n319_), .B2(new_n263_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n323_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n277_), .B1(new_n325_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n320_), .A2(new_n324_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n277_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n326_), .A2(new_n328_), .A3(new_n323_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n331_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n330_), .A2(KEYINPUT27), .A3(new_n334_), .ZN(new_n335_));
  AND3_X1   g134(.A1(new_n326_), .A2(new_n328_), .A3(new_n323_), .ZN(new_n336_));
  OR2_X1    g135(.A1(new_n317_), .A2(new_n303_), .ZN(new_n337_));
  AOI22_X1  g136(.A1(new_n309_), .A2(new_n337_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n327_), .B1(new_n338_), .B2(new_n264_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n323_), .B1(new_n339_), .B2(new_n311_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n277_), .B1(new_n336_), .B2(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(KEYINPUT27), .B1(new_n341_), .B2(new_n334_), .ZN(new_n342_));
  NOR3_X1   g141(.A1(new_n335_), .A2(new_n342_), .A3(KEYINPUT91), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT91), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT27), .ZN(new_n345_));
  NOR3_X1   g144(.A1(new_n336_), .A2(new_n340_), .A3(new_n277_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n332_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n345_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n330_), .A2(KEYINPUT27), .A3(new_n334_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n344_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n272_), .B1(new_n343_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT92), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT91), .B1(new_n335_), .B2(new_n342_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n348_), .A2(new_n344_), .A3(new_n349_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT92), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n355_), .A2(new_n356_), .A3(new_n272_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n352_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G71gat), .B(G99gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(G43gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n319_), .B(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(G127gat), .B(G134gat), .Z(new_n362_));
  XOR2_X1   g161(.A(G113gat), .B(G120gat), .Z(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n361_), .B(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G227gat), .A2(G233gat), .ZN(new_n367_));
  INV_X1    g166(.A(G15gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT30), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT31), .ZN(new_n371_));
  XOR2_X1   g170(.A(new_n366_), .B(new_n371_), .Z(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G1gat), .B(G29gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(G85gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT0), .B(G57gat), .ZN(new_n376_));
  XOR2_X1   g175(.A(new_n375_), .B(new_n376_), .Z(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT4), .ZN(new_n379_));
  AOI211_X1 g178(.A(new_n218_), .B(new_n220_), .C1(new_n211_), .C2(new_n214_), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n365_), .B(KEYINPUT88), .C1(new_n380_), .C2(new_n228_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n222_), .A2(new_n229_), .A3(new_n364_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n379_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n364_), .B1(new_n222_), .B2(new_n229_), .ZN(new_n384_));
  AOI21_X1  g183(.A(KEYINPUT4), .B1(new_n384_), .B2(KEYINPUT88), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G225gat), .A2(G233gat), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n382_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n390_), .A2(new_n384_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n391_), .A2(new_n388_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n378_), .B1(new_n389_), .B2(new_n393_), .ZN(new_n394_));
  NOR3_X1   g193(.A1(new_n383_), .A2(new_n385_), .A3(new_n387_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n395_), .A2(new_n392_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n378_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n394_), .B1(new_n397_), .B2(KEYINPUT90), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT90), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n396_), .A2(new_n399_), .A3(new_n378_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n373_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n332_), .A2(KEYINPUT32), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n403_), .B1(new_n336_), .B2(new_n340_), .ZN(new_n404_));
  OR3_X1    g203(.A1(new_n325_), .A2(new_n329_), .A3(new_n403_), .ZN(new_n405_));
  AOI22_X1  g204(.A1(new_n398_), .A2(new_n400_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NOR3_X1   g205(.A1(new_n394_), .A2(KEYINPUT89), .A3(KEYINPUT33), .ZN(new_n407_));
  OAI211_X1 g206(.A(KEYINPUT33), .B(new_n377_), .C1(new_n395_), .C2(new_n392_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n377_), .B1(new_n391_), .B2(new_n388_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n409_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n408_), .A2(new_n341_), .A3(new_n334_), .A4(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT89), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n377_), .B1(new_n395_), .B2(new_n392_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT33), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n412_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NOR3_X1   g214(.A1(new_n407_), .A2(new_n411_), .A3(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n272_), .B1(new_n406_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n401_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n418_), .A2(new_n348_), .A3(new_n349_), .A4(new_n271_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n358_), .A2(new_n402_), .B1(new_n373_), .B2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G1gat), .B(G8gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT75), .ZN(new_n423_));
  INV_X1    g222(.A(G22gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n368_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G15gat), .A2(G22gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G1gat), .A2(G8gat), .ZN(new_n427_));
  AOI22_X1  g226(.A1(new_n425_), .A2(new_n426_), .B1(KEYINPUT14), .B2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n423_), .B(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G29gat), .B(G36gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT74), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G43gat), .B(G50gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n430_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n433_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n432_), .B(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n429_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n435_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G229gat), .A2(G233gat), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n434_), .A2(KEYINPUT15), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT15), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n437_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n443_), .A2(new_n445_), .A3(new_n430_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n446_), .A2(new_n438_), .A3(new_n440_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n442_), .A2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G113gat), .B(G141gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G169gat), .B(G197gat), .ZN(new_n450_));
  XOR2_X1   g249(.A(new_n449_), .B(new_n450_), .Z(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n448_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n442_), .A2(new_n447_), .A3(new_n451_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n421_), .A2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT10), .B(G99gat), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT65), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(new_n242_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G99gat), .A2(G106gat), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT6), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G85gat), .B(G92gat), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n466_), .B1(new_n467_), .B2(KEYINPUT9), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT66), .ZN(new_n469_));
  OR2_X1    g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n469_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n461_), .A2(new_n465_), .A3(new_n470_), .A4(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT8), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT69), .ZN(new_n474_));
  INV_X1    g273(.A(G99gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(new_n242_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n477_));
  OR2_X1    g276(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n476_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n480_), .B1(new_n475_), .B2(new_n242_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n474_), .B1(new_n479_), .B2(new_n481_), .ZN(new_n482_));
  AND2_X1   g281(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n475_), .B(new_n242_), .C1(new_n483_), .C2(new_n480_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n478_), .A2(new_n476_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n484_), .A2(KEYINPUT69), .A3(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n482_), .A2(new_n486_), .A3(new_n465_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G85gat), .B(G92gat), .Z(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT68), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT68), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n467_), .A2(new_n490_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n473_), .B1(new_n487_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n484_), .A2(new_n485_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n494_), .A2(new_n464_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n489_), .A2(new_n491_), .ZN(new_n496_));
  NOR3_X1   g295(.A1(new_n495_), .A2(new_n496_), .A3(KEYINPUT8), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n472_), .B1(new_n493_), .B2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(new_n443_), .A3(new_n445_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G232gat), .A2(G233gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  OAI221_X1 g302(.A(new_n499_), .B1(KEYINPUT35), .B2(new_n503_), .C1(new_n498_), .C2(new_n434_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(KEYINPUT35), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n504_), .A2(new_n506_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G190gat), .B(G218gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G134gat), .B(G162gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(new_n512_), .B(KEYINPUT36), .Z(new_n513_));
  NAND2_X1  g312(.A1(new_n509_), .A2(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n512_), .A2(KEYINPUT36), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n507_), .A2(new_n515_), .A3(new_n508_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT37), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT37), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n514_), .A2(new_n519_), .A3(new_n516_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  XOR2_X1   g320(.A(G127gat), .B(G155gat), .Z(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G183gat), .B(G211gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT17), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n526_), .A2(KEYINPUT17), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT11), .ZN(new_n529_));
  OR2_X1    g328(.A1(KEYINPUT70), .A2(G71gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(KEYINPUT70), .A2(G71gat), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n240_), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n240_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n529_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n534_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n536_), .A2(KEYINPUT11), .A3(new_n532_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G57gat), .B(G64gat), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n535_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n538_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n536_), .A2(KEYINPUT11), .A3(new_n532_), .A4(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G231gat), .A2(G233gat), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n542_), .A2(G231gat), .A3(G233gat), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n545_), .A2(new_n430_), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n430_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n527_), .B(new_n528_), .C1(new_n548_), .C2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n549_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n527_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(new_n547_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n550_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n521_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G230gat), .A2(G233gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT64), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n498_), .A2(new_n543_), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n472_), .B(new_n542_), .C1(new_n493_), .C2(new_n497_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n560_), .A2(KEYINPUT12), .A3(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(KEYINPUT12), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n492_), .B(new_n473_), .C1(new_n494_), .C2(new_n464_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n464_), .B1(new_n494_), .B2(new_n474_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n496_), .B1(new_n565_), .B2(new_n486_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n564_), .B1(new_n566_), .B2(new_n473_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n542_), .B1(new_n567_), .B2(new_n472_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n563_), .A2(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n559_), .B1(new_n562_), .B2(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n558_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G120gat), .B(G148gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT5), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G176gat), .B(G204gat), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n574_), .B(new_n575_), .Z(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n577_), .A2(KEYINPUT71), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT72), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n572_), .B(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT13), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n572_), .B(new_n579_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT13), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n556_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n457_), .A2(new_n587_), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n588_), .B(KEYINPUT93), .Z(new_n589_));
  INV_X1    g388(.A(G1gat), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n589_), .A2(new_n590_), .A3(new_n401_), .ZN(new_n591_));
  XOR2_X1   g390(.A(KEYINPUT94), .B(KEYINPUT38), .Z(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n586_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(new_n455_), .A3(new_n555_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT95), .ZN(new_n596_));
  INV_X1    g395(.A(new_n517_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n421_), .A2(new_n597_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n599_), .A2(new_n401_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n593_), .B1(new_n590_), .B2(new_n600_), .ZN(G1324gat));
  INV_X1    g400(.A(G8gat), .ZN(new_n602_));
  INV_X1    g401(.A(new_n355_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n602_), .B1(new_n599_), .B2(new_n603_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT39), .Z(new_n605_));
  NAND3_X1  g404(.A1(new_n589_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT40), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(G1325gat));
  AOI21_X1  g408(.A(new_n368_), .B1(new_n599_), .B2(new_n372_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT41), .ZN(new_n611_));
  INV_X1    g410(.A(new_n588_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n612_), .A2(new_n368_), .A3(new_n372_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(G1326gat));
  AOI21_X1  g413(.A(new_n424_), .B1(new_n599_), .B2(new_n271_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT42), .Z(new_n616_));
  NAND3_X1  g415(.A1(new_n612_), .A2(new_n424_), .A3(new_n271_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(G1327gat));
  NOR2_X1   g417(.A1(new_n517_), .A2(new_n555_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT97), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n620_), .A2(new_n586_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n457_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(G29gat), .B1(new_n623_), .B2(new_n401_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n586_), .A2(new_n456_), .A3(new_n555_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT43), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n356_), .B1(new_n355_), .B2(new_n272_), .ZN(new_n627_));
  AOI211_X1 g426(.A(KEYINPUT92), .B(new_n271_), .C1(new_n353_), .C2(new_n354_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n402_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n420_), .A2(new_n373_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n521_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n626_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  AOI211_X1 g432(.A(KEYINPUT43), .B(new_n521_), .C1(new_n629_), .C2(new_n630_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n625_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT96), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT44), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n625_), .ZN(new_n638_));
  OAI21_X1  g437(.A(KEYINPUT43), .B1(new_n421_), .B2(new_n521_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n631_), .A2(new_n626_), .A3(new_n632_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n638_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT96), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n637_), .A2(new_n642_), .ZN(new_n643_));
  OAI211_X1 g442(.A(KEYINPUT44), .B(new_n625_), .C1(new_n633_), .C2(new_n634_), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n644_), .A2(G29gat), .A3(new_n401_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n624_), .B1(new_n643_), .B2(new_n645_), .ZN(G1328gat));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n647_));
  XNOR2_X1  g446(.A(KEYINPUT99), .B(KEYINPUT45), .ZN(new_n648_));
  INV_X1    g447(.A(G36gat), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n603_), .A2(new_n649_), .ZN(new_n650_));
  OR3_X1    g449(.A1(new_n622_), .A2(new_n648_), .A3(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n648_), .B1(new_n622_), .B2(new_n650_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n355_), .B1(new_n641_), .B2(KEYINPUT44), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT44), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n655_), .B1(new_n641_), .B2(KEYINPUT96), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n635_), .A2(new_n636_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n654_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT98), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n649_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  OAI211_X1 g459(.A(KEYINPUT98), .B(new_n654_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n653_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  XOR2_X1   g461(.A(KEYINPUT100), .B(KEYINPUT46), .Z(new_n663_));
  OAI21_X1  g462(.A(new_n647_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n653_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n644_), .A2(new_n603_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(new_n637_), .B2(new_n642_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G36gat), .B1(new_n667_), .B2(KEYINPUT98), .ZN(new_n668_));
  INV_X1    g467(.A(new_n661_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n665_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n663_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n670_), .A2(KEYINPUT101), .A3(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n662_), .A2(KEYINPUT46), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n664_), .A2(new_n672_), .A3(new_n673_), .ZN(G1329gat));
  AOI21_X1  g473(.A(G43gat), .B1(new_n623_), .B2(new_n372_), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n644_), .A2(G43gat), .A3(new_n372_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n643_), .B2(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(KEYINPUT102), .B(KEYINPUT47), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n677_), .B(new_n678_), .ZN(G1330gat));
  OR3_X1    g478(.A1(new_n622_), .A2(G50gat), .A3(new_n272_), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n643_), .A2(new_n271_), .A3(new_n644_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G50gat), .B1(new_n681_), .B2(new_n682_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n680_), .B1(new_n684_), .B2(new_n685_), .ZN(G1331gat));
  NOR2_X1   g485(.A1(new_n556_), .A2(new_n594_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT104), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n688_), .A2(new_n421_), .A3(new_n455_), .ZN(new_n689_));
  INV_X1    g488(.A(G57gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n689_), .A2(new_n690_), .A3(new_n401_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n598_), .A2(new_n456_), .A3(new_n586_), .A4(new_n555_), .ZN(new_n692_));
  OAI21_X1  g491(.A(G57gat), .B1(new_n692_), .B2(new_n418_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1332gat));
  OAI21_X1  g493(.A(G64gat), .B1(new_n692_), .B2(new_n355_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT48), .ZN(new_n696_));
  INV_X1    g495(.A(G64gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n689_), .A2(new_n697_), .A3(new_n603_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(G1333gat));
  OAI21_X1  g498(.A(G71gat), .B1(new_n692_), .B2(new_n373_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT49), .ZN(new_n701_));
  INV_X1    g500(.A(G71gat), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n689_), .A2(new_n702_), .A3(new_n372_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT105), .Z(G1334gat));
  OAI21_X1  g504(.A(G78gat), .B1(new_n692_), .B2(new_n272_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT50), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n689_), .A2(new_n240_), .A3(new_n271_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1335gat));
  NOR2_X1   g508(.A1(new_n421_), .A2(new_n455_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n620_), .A2(new_n594_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(G85gat), .B1(new_n713_), .B2(new_n401_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n639_), .A2(new_n640_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n594_), .A2(new_n455_), .A3(new_n555_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n401_), .A2(G85gat), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT106), .Z(new_n720_));
  AOI21_X1  g519(.A(new_n714_), .B1(new_n718_), .B2(new_n720_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT107), .Z(G1336gat));
  OAI21_X1  g521(.A(G92gat), .B1(new_n717_), .B2(new_n355_), .ZN(new_n723_));
  OR2_X1    g522(.A1(new_n355_), .A2(G92gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n723_), .B1(new_n712_), .B2(new_n724_), .ZN(G1337gat));
  NAND2_X1  g524(.A1(new_n372_), .A2(new_n460_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT51), .ZN(new_n727_));
  OAI22_X1  g526(.A1(new_n712_), .A2(new_n726_), .B1(KEYINPUT108), .B2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n718_), .A2(new_n372_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(G99gat), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n727_), .A2(KEYINPUT108), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n730_), .B(new_n731_), .Z(G1338gat));
  XNOR2_X1  g531(.A(KEYINPUT109), .B(KEYINPUT53), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n718_), .A2(new_n271_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(G106gat), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT52), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n713_), .A2(new_n242_), .A3(new_n271_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n733_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n735_), .A2(KEYINPUT52), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT52), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n734_), .B2(G106gat), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n737_), .B(new_n733_), .C1(new_n739_), .C2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n738_), .A2(new_n743_), .ZN(G1339gat));
  INV_X1    g543(.A(KEYINPUT121), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n456_), .A2(new_n555_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT110), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n594_), .A2(new_n521_), .A3(new_n747_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n748_), .A2(KEYINPUT111), .A3(KEYINPUT54), .ZN(new_n749_));
  AOI21_X1  g548(.A(KEYINPUT111), .B1(new_n748_), .B2(KEYINPUT54), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n748_), .A2(KEYINPUT54), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n749_), .A2(new_n750_), .A3(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n439_), .A2(new_n440_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n446_), .A2(new_n438_), .A3(new_n441_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT115), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n753_), .A2(new_n754_), .A3(new_n755_), .A4(new_n452_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n753_), .A2(new_n754_), .A3(new_n452_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT115), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n581_), .A2(new_n454_), .A3(new_n756_), .A4(new_n758_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n570_), .A2(new_n571_), .A3(new_n576_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n456_), .A2(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n563_), .A2(new_n568_), .ZN(new_n762_));
  AOI211_X1 g561(.A(KEYINPUT12), .B(new_n542_), .C1(new_n567_), .C2(new_n472_), .ZN(new_n763_));
  OAI21_X1  g562(.A(KEYINPUT112), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n562_), .A2(new_n569_), .A3(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n764_), .A2(new_n559_), .A3(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n558_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n768_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n570_), .A2(new_n771_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n769_), .A2(new_n770_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n767_), .A2(new_n773_), .A3(new_n774_), .A4(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n576_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n778_), .A2(KEYINPUT56), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n761_), .B1(new_n777_), .B2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n779_), .B1(new_n776_), .B2(new_n576_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n759_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n783_), .A2(KEYINPUT57), .A3(new_n517_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT119), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n783_), .A2(KEYINPUT119), .A3(KEYINPUT57), .A4(new_n517_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n758_), .A2(new_n454_), .A3(new_n756_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n584_), .A2(new_n789_), .ZN(new_n790_));
  OR2_X1    g589(.A1(new_n456_), .A2(new_n760_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n775_), .B1(new_n570_), .B2(new_n771_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n768_), .A2(new_n772_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n577_), .B1(new_n794_), .B2(new_n767_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n791_), .B1(new_n795_), .B2(new_n779_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n782_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n790_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(KEYINPUT116), .B1(new_n798_), .B2(new_n597_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n783_), .A2(new_n801_), .A3(new_n517_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n799_), .A2(new_n800_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT56), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n776_), .A2(new_n804_), .A3(new_n576_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n789_), .A2(new_n760_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n804_), .B1(new_n776_), .B2(new_n576_), .ZN(new_n808_));
  OAI211_X1 g607(.A(KEYINPUT117), .B(KEYINPUT58), .C1(new_n807_), .C2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n777_), .A2(KEYINPUT56), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n811_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT58), .B1(new_n812_), .B2(KEYINPUT117), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n632_), .B1(new_n810_), .B2(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n788_), .A2(new_n803_), .A3(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n752_), .B1(new_n815_), .B2(new_n554_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n358_), .A2(new_n401_), .A3(new_n372_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n816_), .A2(KEYINPUT59), .A3(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(G113gat), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n456_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT118), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n814_), .A2(new_n822_), .ZN(new_n823_));
  OAI211_X1 g622(.A(KEYINPUT118), .B(new_n632_), .C1(new_n810_), .C2(new_n813_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n823_), .A2(new_n788_), .A3(new_n803_), .A4(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n752_), .B1(new_n825_), .B2(new_n554_), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT59), .B1(new_n826_), .B2(new_n817_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT120), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  OAI211_X1 g628(.A(KEYINPUT120), .B(KEYINPUT59), .C1(new_n826_), .C2(new_n817_), .ZN(new_n830_));
  AOI211_X1 g629(.A(new_n818_), .B(new_n821_), .C1(new_n829_), .C2(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n826_), .A2(new_n817_), .ZN(new_n832_));
  AOI21_X1  g631(.A(G113gat), .B1(new_n832_), .B2(new_n455_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n745_), .B1(new_n831_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n818_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n827_), .A2(new_n828_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n830_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n835_), .B(new_n820_), .C1(new_n836_), .C2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n833_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n838_), .A2(KEYINPUT121), .A3(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n834_), .A2(new_n840_), .ZN(G1340gat));
  INV_X1    g640(.A(KEYINPUT60), .ZN(new_n842_));
  AOI21_X1  g641(.A(G120gat), .B1(new_n586_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT122), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n843_), .A2(new_n844_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n846_), .B1(new_n842_), .B2(G120gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n832_), .A2(new_n845_), .A3(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n818_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n849_), .A2(new_n586_), .ZN(new_n850_));
  INV_X1    g649(.A(G120gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n848_), .B1(new_n850_), .B2(new_n851_), .ZN(G1341gat));
  AOI21_X1  g651(.A(G127gat), .B1(new_n832_), .B2(new_n555_), .ZN(new_n853_));
  XOR2_X1   g652(.A(KEYINPUT123), .B(G127gat), .Z(new_n854_));
  NAND2_X1  g653(.A1(new_n555_), .A2(new_n854_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(KEYINPUT124), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n853_), .B1(new_n849_), .B2(new_n856_), .ZN(G1342gat));
  INV_X1    g656(.A(G134gat), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n521_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  AOI211_X1 g659(.A(new_n818_), .B(new_n860_), .C1(new_n829_), .C2(new_n830_), .ZN(new_n861_));
  AOI21_X1  g660(.A(G134gat), .B1(new_n832_), .B2(new_n597_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT125), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n835_), .B(new_n859_), .C1(new_n836_), .C2(new_n837_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT125), .ZN(new_n865_));
  INV_X1    g664(.A(new_n862_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n864_), .A2(new_n865_), .A3(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n863_), .A2(new_n867_), .ZN(G1343gat));
  NOR2_X1   g667(.A1(new_n272_), .A2(new_n372_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n826_), .A2(new_n870_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n603_), .A2(new_n418_), .ZN(new_n872_));
  AND3_X1   g671(.A1(new_n871_), .A2(KEYINPUT126), .A3(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(KEYINPUT126), .B1(new_n871_), .B2(new_n872_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n455_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G141gat), .ZN(G1344gat));
  OAI21_X1  g675(.A(new_n586_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(G148gat), .ZN(G1345gat));
  OAI21_X1  g677(.A(new_n555_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(KEYINPUT61), .B(G155gat), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n879_), .B(new_n880_), .ZN(G1346gat));
  NOR2_X1   g680(.A1(new_n873_), .A2(new_n874_), .ZN(new_n882_));
  OAI21_X1  g681(.A(G162gat), .B1(new_n882_), .B2(new_n521_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n597_), .A2(new_n217_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n882_), .B2(new_n884_), .ZN(G1347gat));
  NOR2_X1   g684(.A1(new_n355_), .A2(new_n401_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n373_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n816_), .A2(new_n271_), .A3(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n281_), .B1(new_n890_), .B2(new_n455_), .ZN(new_n891_));
  OR2_X1    g690(.A1(new_n891_), .A2(KEYINPUT62), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n455_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n893_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n890_), .A2(new_n308_), .A3(new_n455_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n892_), .A2(new_n894_), .A3(new_n895_), .ZN(G1348gat));
  AOI21_X1  g695(.A(G176gat), .B1(new_n890_), .B2(new_n586_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n826_), .A2(new_n271_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n889_), .A2(new_n282_), .A3(new_n594_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n897_), .B1(new_n898_), .B2(new_n899_), .ZN(G1349gat));
  INV_X1    g699(.A(new_n890_), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n901_), .A2(new_n278_), .A3(new_n554_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n898_), .A2(new_n555_), .A3(new_n888_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n902_), .B1(new_n291_), .B2(new_n903_), .ZN(G1350gat));
  OAI21_X1  g703(.A(G190gat), .B1(new_n901_), .B2(new_n521_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n890_), .A2(new_n279_), .A3(new_n597_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1351gat));
  NOR3_X1   g706(.A1(new_n826_), .A2(new_n870_), .A3(new_n887_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(new_n455_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n586_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G204gat), .ZN(G1353gat));
  AND2_X1   g711(.A1(new_n908_), .A2(new_n555_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n914_));
  AND2_X1   g713(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n913_), .B1(new_n914_), .B2(new_n915_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n916_), .B1(new_n913_), .B2(new_n914_), .ZN(G1354gat));
  NAND2_X1  g716(.A1(new_n908_), .A2(new_n597_), .ZN(new_n918_));
  XOR2_X1   g717(.A(KEYINPUT127), .B(G218gat), .Z(new_n919_));
  NOR2_X1   g718(.A1(new_n521_), .A2(new_n919_), .ZN(new_n920_));
  AOI22_X1  g719(.A1(new_n918_), .A2(new_n919_), .B1(new_n908_), .B2(new_n920_), .ZN(G1355gat));
endmodule


