//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 0 1 1 1 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 0 1 0 1 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n757_, new_n758_,
    new_n759_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n914_, new_n915_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n922_, new_n923_, new_n924_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT94), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G197gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G204gat), .ZN(new_n206_));
  INV_X1    g005(.A(G204gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G197gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n209_), .A2(KEYINPUT21), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n204_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT92), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n206_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT91), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n208_), .A2(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n205_), .A2(KEYINPUT92), .A3(G204gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n207_), .A2(KEYINPUT91), .A3(G197gat), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n213_), .A2(new_n215_), .A3(new_n216_), .A4(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT21), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT93), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT93), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n218_), .A2(new_n221_), .A3(KEYINPUT21), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n211_), .A2(new_n220_), .A3(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n204_), .A2(KEYINPUT21), .A3(new_n209_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT95), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n223_), .A2(KEYINPUT95), .A3(new_n224_), .ZN(new_n228_));
  XOR2_X1   g027(.A(KEYINPUT25), .B(G183gat), .Z(new_n229_));
  XOR2_X1   g028(.A(KEYINPUT85), .B(KEYINPUT26), .Z(new_n230_));
  AOI21_X1  g029(.A(new_n229_), .B1(G190gat), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G190gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT26), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT84), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n231_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G169gat), .A2(G176gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT24), .ZN(new_n237_));
  NOR2_X1   g036(.A1(G169gat), .A2(G176gat), .ZN(new_n238_));
  MUX2_X1   g037(.A(new_n237_), .B(KEYINPUT24), .S(new_n238_), .Z(new_n239_));
  NAND2_X1  g038(.A1(G183gat), .A2(G190gat), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT23), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n235_), .A2(new_n239_), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(G176gat), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT86), .ZN(new_n246_));
  INV_X1    g045(.A(G169gat), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n246_), .B1(new_n247_), .B2(KEYINPUT22), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT22), .B(G169gat), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n245_), .B(new_n248_), .C1(new_n249_), .C2(new_n246_), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT87), .B1(new_n250_), .B2(new_n236_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(KEYINPUT87), .A3(new_n236_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(G183gat), .A2(G190gat), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n253_), .B1(new_n241_), .B2(new_n240_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n254_), .B1(new_n241_), .B2(new_n240_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n252_), .A2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n244_), .B1(new_n251_), .B2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n227_), .A2(new_n228_), .A3(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT26), .B(G190gat), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n260_), .A2(new_n229_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n261_), .A2(new_n242_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n236_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n263_), .B1(new_n249_), .B2(new_n245_), .ZN(new_n264_));
  AOI22_X1  g063(.A1(new_n262_), .A2(new_n239_), .B1(new_n255_), .B2(new_n264_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n223_), .A2(new_n265_), .A3(KEYINPUT97), .A4(new_n224_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G226gat), .A2(G233gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT19), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n266_), .A2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n223_), .A2(new_n224_), .A3(new_n265_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT97), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n258_), .A2(new_n270_), .A3(KEYINPUT20), .A4(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT98), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n273_), .A2(new_n269_), .A3(new_n266_), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n277_), .A2(KEYINPUT98), .A3(KEYINPUT20), .A4(new_n258_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n257_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n265_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n225_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT20), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n268_), .B1(new_n279_), .B2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n276_), .A2(new_n278_), .A3(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(G8gat), .B(G36gat), .Z(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G64gat), .B(G92gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n284_), .A2(new_n290_), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n276_), .A2(new_n278_), .A3(new_n283_), .A4(new_n289_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(KEYINPUT100), .A3(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT27), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT100), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n284_), .A2(new_n295_), .A3(new_n290_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n293_), .A2(new_n294_), .A3(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G127gat), .B(G134gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT88), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n298_), .A2(new_n299_), .ZN(new_n301_));
  XOR2_X1   g100(.A(G113gat), .B(G120gat), .Z(new_n302_));
  OR3_X1    g101(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n302_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306_));
  NOR2_X1   g105(.A1(G155gat), .A2(G162gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(G141gat), .A2(G148gat), .ZN(new_n309_));
  XOR2_X1   g108(.A(new_n309_), .B(KEYINPUT3), .Z(new_n310_));
  NAND2_X1  g109(.A1(G141gat), .A2(G148gat), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n311_), .B(KEYINPUT2), .Z(new_n312_));
  OAI211_X1 g111(.A(new_n306_), .B(new_n308_), .C1(new_n310_), .C2(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n307_), .B1(KEYINPUT1), .B2(new_n306_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n314_), .B1(KEYINPUT1), .B2(new_n306_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n309_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n315_), .A2(new_n316_), .A3(new_n311_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n313_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n305_), .A2(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT101), .B1(new_n319_), .B2(KEYINPUT4), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT101), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT4), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n305_), .A2(new_n318_), .A3(new_n321_), .A4(new_n322_), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n303_), .A2(new_n313_), .A3(new_n317_), .A4(new_n304_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n319_), .A2(new_n324_), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n320_), .B(new_n323_), .C1(new_n322_), .C2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G225gat), .A2(G233gat), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n325_), .A2(new_n327_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G1gat), .B(G29gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(G85gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT0), .B(G57gat), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n333_), .B(new_n334_), .Z(new_n335_));
  NAND2_X1  g134(.A1(new_n331_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n335_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n329_), .A2(new_n337_), .A3(new_n330_), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n258_), .A2(KEYINPUT20), .A3(new_n271_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(new_n268_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n257_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n228_), .ZN(new_n343_));
  AOI21_X1  g142(.A(KEYINPUT95), .B1(new_n223_), .B2(new_n224_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n342_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n345_), .A2(KEYINPUT20), .A3(new_n281_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n341_), .B1(new_n268_), .B2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n290_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n348_), .A2(KEYINPUT27), .A3(new_n292_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n297_), .A2(new_n339_), .A3(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n318_), .A2(KEYINPUT29), .ZN(new_n351_));
  XOR2_X1   g150(.A(G22gat), .B(G50gat), .Z(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NOR3_X1   g155(.A1(new_n318_), .A2(KEYINPUT29), .A3(new_n352_), .ZN(new_n357_));
  NOR3_X1   g156(.A1(new_n354_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT96), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n356_), .B1(new_n354_), .B2(new_n357_), .ZN(new_n361_));
  AND3_X1   g160(.A1(new_n359_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n360_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G228gat), .A2(G233gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n318_), .A2(KEYINPUT29), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n227_), .A2(new_n365_), .A3(new_n366_), .A4(new_n228_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n225_), .A2(new_n366_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n368_), .A2(G228gat), .A3(G233gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(G78gat), .ZN(new_n371_));
  INV_X1    g170(.A(G106gat), .ZN(new_n372_));
  INV_X1    g171(.A(G78gat), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n367_), .A2(new_n373_), .A3(new_n369_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n371_), .A2(new_n372_), .A3(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n372_), .B1(new_n371_), .B2(new_n374_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n364_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n377_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(new_n362_), .A3(new_n375_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n350_), .A2(new_n381_), .ZN(new_n382_));
  XOR2_X1   g181(.A(new_n305_), .B(KEYINPUT31), .Z(new_n383_));
  XNOR2_X1  g182(.A(G71gat), .B(G99gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(G43gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n257_), .B(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G227gat), .A2(G233gat), .ZN(new_n387_));
  INV_X1    g186(.A(G15gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT30), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n386_), .B(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT89), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n383_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n393_), .B1(new_n392_), .B2(new_n391_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n391_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n395_), .A2(KEYINPUT89), .A3(new_n383_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n337_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n319_), .A2(new_n328_), .A3(new_n324_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n337_), .B(new_n400_), .C1(new_n326_), .C2(new_n328_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n399_), .B1(KEYINPUT33), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT33), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT102), .B1(new_n336_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT102), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n399_), .A2(new_n405_), .A3(KEYINPUT33), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n402_), .B1(new_n404_), .B2(new_n406_), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n268_), .A2(new_n346_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n289_), .B1(new_n408_), .B2(new_n278_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n292_), .A2(KEYINPUT100), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n296_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n407_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n289_), .A2(KEYINPUT32), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  AOI22_X1  g214(.A1(new_n336_), .A2(new_n338_), .B1(new_n347_), .B2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n408_), .A2(new_n278_), .A3(new_n414_), .ZN(new_n417_));
  AOI22_X1  g216(.A1(new_n378_), .A2(new_n380_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n398_), .B1(new_n413_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n382_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT103), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n297_), .A2(new_n349_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n423_), .A2(new_n381_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n424_), .A2(new_n339_), .A3(new_n398_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n382_), .A2(new_n419_), .A3(KEYINPUT103), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n422_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G1gat), .B(G8gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G1gat), .A2(G8gat), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT78), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n429_), .A2(new_n430_), .A3(KEYINPUT14), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n388_), .A2(G22gat), .ZN(new_n432_));
  INV_X1    g231(.A(G22gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(G15gat), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n431_), .A2(new_n432_), .A3(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n430_), .B1(new_n429_), .B2(KEYINPUT14), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n428_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n428_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n436_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G15gat), .B(G22gat), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n438_), .A2(new_n439_), .A3(new_n431_), .A4(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n437_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G231gat), .A2(G233gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G71gat), .B(G78gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G57gat), .B(G64gat), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n445_), .B1(KEYINPUT11), .B2(new_n446_), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n446_), .A2(KEYINPUT11), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n446_), .A2(new_n445_), .A3(KEYINPUT11), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n444_), .B(new_n452_), .ZN(new_n453_));
  XOR2_X1   g252(.A(G127gat), .B(G155gat), .Z(new_n454_));
  XNOR2_X1  g253(.A(G183gat), .B(G211gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT17), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n453_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n453_), .A2(KEYINPUT17), .A3(new_n458_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT80), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n462_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n460_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  AND2_X1   g265(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n467_));
  NOR2_X1   g266(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n468_));
  OAI22_X1  g267(.A1(new_n467_), .A2(new_n468_), .B1(G99gat), .B2(G106gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G99gat), .A2(G106gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT6), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT6), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n472_), .A2(G99gat), .A3(G106gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(G99gat), .A2(G106gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n469_), .A2(new_n474_), .A3(new_n477_), .ZN(new_n478_));
  XOR2_X1   g277(.A(G85gat), .B(G92gat), .Z(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT8), .ZN(new_n481_));
  XOR2_X1   g280(.A(KEYINPUT10), .B(G99gat), .Z(new_n482_));
  XOR2_X1   g281(.A(KEYINPUT64), .B(G106gat), .Z(new_n483_));
  INV_X1    g282(.A(G85gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT65), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT65), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(G85gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(G92gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n489_), .A2(KEYINPUT9), .ZN(new_n490_));
  AOI22_X1  g289(.A1(new_n482_), .A2(new_n483_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n491_));
  AOI22_X1  g290(.A1(new_n479_), .A2(KEYINPUT9), .B1(new_n471_), .B2(new_n473_), .ZN(new_n492_));
  AOI22_X1  g291(.A1(new_n480_), .A2(new_n481_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT67), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT66), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT7), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n475_), .B1(new_n497_), .B2(new_n476_), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n475_), .A2(new_n476_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n494_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n469_), .A2(KEYINPUT67), .A3(new_n477_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(new_n501_), .A3(new_n474_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n479_), .A2(KEYINPUT8), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(G43gat), .B(G50gat), .Z(new_n506_));
  INV_X1    g305(.A(G36gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(G29gat), .ZN(new_n508_));
  INV_X1    g307(.A(G29gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(G36gat), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n508_), .A2(new_n510_), .A3(KEYINPUT71), .ZN(new_n511_));
  AOI21_X1  g310(.A(KEYINPUT71), .B1(new_n508_), .B2(new_n510_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n506_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT71), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n509_), .A2(G36gat), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n507_), .A2(G29gat), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n514_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n508_), .A2(new_n510_), .A3(KEYINPUT71), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G43gat), .B(G50gat), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n513_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n493_), .A2(new_n505_), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT72), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NOR3_X1   g323(.A1(new_n511_), .A2(new_n512_), .A3(new_n506_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n519_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT15), .ZN(new_n528_));
  AOI21_X1  g327(.A(KEYINPUT15), .B1(new_n513_), .B2(new_n520_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n480_), .A2(new_n481_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n491_), .A2(new_n492_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n474_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n469_), .A2(new_n477_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n534_), .B1(new_n535_), .B2(new_n494_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n503_), .B1(new_n536_), .B2(new_n501_), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n528_), .B(new_n530_), .C1(new_n533_), .C2(new_n537_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n493_), .A2(new_n505_), .A3(KEYINPUT72), .A4(new_n521_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G232gat), .A2(G233gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT34), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT35), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n524_), .A2(new_n538_), .A3(new_n539_), .A4(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n542_), .A2(new_n543_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT15), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n521_), .A2(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n549_), .A2(new_n529_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n493_), .A2(new_n505_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n550_), .A2(new_n551_), .B1(new_n543_), .B2(new_n542_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n546_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n552_), .A2(new_n553_), .A3(new_n539_), .A4(new_n524_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n547_), .A2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G190gat), .B(G218gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G134gat), .B(G162gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n558_), .B(KEYINPUT36), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT73), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n555_), .A2(KEYINPUT74), .A3(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n558_), .A2(KEYINPUT36), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n547_), .A2(new_n554_), .A3(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(KEYINPUT74), .B1(new_n555_), .B2(new_n560_), .ZN(new_n565_));
  OAI21_X1  g364(.A(KEYINPUT37), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT75), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  OAI211_X1 g367(.A(KEYINPUT75), .B(KEYINPUT37), .C1(new_n564_), .C2(new_n565_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT77), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT76), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n547_), .A2(new_n572_), .A3(new_n554_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(new_n560_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n572_), .B1(new_n547_), .B2(new_n554_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n571_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n555_), .A2(KEYINPUT76), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n577_), .A2(KEYINPUT77), .A3(new_n560_), .A4(new_n573_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n576_), .A2(new_n563_), .A3(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT37), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n466_), .B1(new_n570_), .B2(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(G120gat), .B(G148gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(G176gat), .B(G204gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(KEYINPUT69), .B(KEYINPUT5), .Z(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT70), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n551_), .A2(new_n452_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(KEYINPUT12), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT12), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n551_), .A2(new_n592_), .A3(new_n452_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT68), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n493_), .A2(new_n505_), .A3(new_n451_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G230gat), .A2(G233gat), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n595_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n596_), .A2(new_n595_), .A3(new_n597_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n594_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n590_), .A2(new_n596_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n597_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n589_), .B1(new_n601_), .B2(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n592_), .B1(new_n551_), .B2(new_n452_), .ZN(new_n606_));
  AOI211_X1 g405(.A(KEYINPUT12), .B(new_n451_), .C1(new_n493_), .C2(new_n505_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n600_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n604_), .B(new_n587_), .C1(new_n608_), .C2(new_n598_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n605_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT13), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(KEYINPUT13), .B1(new_n605_), .B2(new_n610_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT83), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n442_), .A2(new_n520_), .A3(new_n513_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n437_), .B(new_n441_), .C1(new_n525_), .C2(new_n526_), .ZN(new_n618_));
  AOI21_X1  g417(.A(KEYINPUT81), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n617_), .A2(new_n618_), .A3(KEYINPUT81), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n620_), .A2(G229gat), .A3(G233gat), .A4(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n550_), .A2(new_n442_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(G229gat), .A2(G233gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT82), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n623_), .A2(new_n618_), .A3(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G113gat), .B(G141gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G169gat), .B(G197gat), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n627_), .B(new_n628_), .Z(new_n629_));
  AND3_X1   g428(.A1(new_n622_), .A2(new_n626_), .A3(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n622_), .B2(new_n626_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n616_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n622_), .A2(new_n626_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n629_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n622_), .A2(new_n626_), .A3(new_n629_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n635_), .A2(KEYINPUT83), .A3(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n632_), .A2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n615_), .A2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n427_), .A2(new_n582_), .A3(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT104), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n339_), .A2(G1gat), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(KEYINPUT105), .B1(new_n641_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT104), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n640_), .B(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT105), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n646_), .A2(new_n647_), .A3(new_n642_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n644_), .A2(KEYINPUT38), .A3(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n426_), .A2(new_n425_), .ZN(new_n650_));
  AOI21_X1  g449(.A(KEYINPUT103), .B1(new_n382_), .B2(new_n419_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n652_), .A2(new_n579_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n639_), .B(KEYINPUT106), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n654_), .A2(new_n466_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G1gat), .B1(new_n656_), .B2(new_n339_), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT38), .B1(new_n644_), .B2(new_n648_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT107), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  AOI211_X1 g459(.A(KEYINPUT107), .B(KEYINPUT38), .C1(new_n644_), .C2(new_n648_), .ZN(new_n661_));
  OAI211_X1 g460(.A(new_n649_), .B(new_n657_), .C1(new_n660_), .C2(new_n661_), .ZN(G1324gat));
  INV_X1    g461(.A(new_n423_), .ZN(new_n663_));
  OR3_X1    g462(.A1(new_n641_), .A2(G8gat), .A3(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G8gat), .B1(new_n656_), .B2(new_n663_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n665_), .A2(KEYINPUT39), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT39), .ZN(new_n667_));
  OAI211_X1 g466(.A(new_n667_), .B(G8gat), .C1(new_n656_), .C2(new_n663_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n664_), .B1(new_n666_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT40), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n664_), .B(KEYINPUT40), .C1(new_n666_), .C2(new_n669_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1325gat));
  OAI21_X1  g473(.A(G15gat), .B1(new_n656_), .B2(new_n397_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT41), .Z(new_n676_));
  NAND3_X1  g475(.A1(new_n646_), .A2(new_n388_), .A3(new_n398_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(G1326gat));
  INV_X1    g477(.A(new_n381_), .ZN(new_n679_));
  OAI21_X1  g478(.A(G22gat), .B1(new_n656_), .B2(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT42), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n646_), .A2(new_n433_), .A3(new_n381_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1327gat));
  NOR2_X1   g482(.A1(new_n654_), .A2(new_n465_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n569_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n555_), .A2(new_n560_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT74), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(new_n563_), .A3(new_n561_), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT75), .B1(new_n690_), .B2(KEYINPUT37), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n576_), .A2(new_n563_), .A3(new_n578_), .ZN(new_n692_));
  OAI22_X1  g491(.A1(new_n686_), .A2(new_n691_), .B1(KEYINPUT37), .B2(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT43), .B1(new_n652_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n695_));
  AOI22_X1  g494(.A1(new_n568_), .A2(new_n569_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n695_), .B(new_n696_), .C1(new_n650_), .C2(new_n651_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n685_), .B1(new_n694_), .B2(new_n697_), .ZN(new_n698_));
  XOR2_X1   g497(.A(KEYINPUT108), .B(KEYINPUT44), .Z(new_n699_));
  OR2_X1    g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n339_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n697_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n695_), .B1(new_n427_), .B2(new_n696_), .ZN(new_n703_));
  OAI211_X1 g502(.A(KEYINPUT44), .B(new_n684_), .C1(new_n702_), .C2(new_n703_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n700_), .A2(G29gat), .A3(new_n701_), .A4(new_n704_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n692_), .A2(new_n465_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n427_), .A2(new_n639_), .A3(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n509_), .B1(new_n707_), .B2(new_n339_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n705_), .A2(new_n708_), .ZN(G1328gat));
  INV_X1    g508(.A(KEYINPUT110), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT46), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n704_), .B(new_n423_), .C1(new_n698_), .C2(new_n699_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(G36gat), .ZN(new_n715_));
  INV_X1    g514(.A(new_n639_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n650_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n717_), .B2(new_n422_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT109), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n663_), .A2(G36gat), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n718_), .A2(new_n719_), .A3(new_n706_), .A4(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n720_), .ZN(new_n722_));
  OAI21_X1  g521(.A(KEYINPUT109), .B1(new_n707_), .B2(new_n722_), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n721_), .A2(new_n723_), .A3(KEYINPUT45), .ZN(new_n724_));
  AOI21_X1  g523(.A(KEYINPUT45), .B1(new_n721_), .B2(new_n723_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  AOI211_X1 g525(.A(new_n712_), .B(new_n713_), .C1(new_n715_), .C2(new_n726_), .ZN(new_n727_));
  AND4_X1   g526(.A1(new_n710_), .A2(new_n715_), .A3(new_n711_), .A4(new_n726_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1329gat));
  INV_X1    g528(.A(G43gat), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n397_), .A2(new_n730_), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n704_), .B(new_n731_), .C1(new_n698_), .C2(new_n699_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n730_), .B1(new_n707_), .B2(new_n397_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g534(.A1(new_n700_), .A2(G50gat), .A3(new_n381_), .A4(new_n704_), .ZN(new_n736_));
  INV_X1    g535(.A(G50gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n737_), .B1(new_n707_), .B2(new_n679_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1331gat));
  INV_X1    g538(.A(new_n615_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n638_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n653_), .A2(new_n465_), .A3(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(G57gat), .B1(new_n743_), .B2(new_n339_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n427_), .A2(new_n742_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n582_), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n339_), .A2(G57gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n744_), .B1(new_n746_), .B2(new_n747_), .ZN(G1332gat));
  OAI21_X1  g547(.A(G64gat), .B1(new_n743_), .B2(new_n663_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT48), .ZN(new_n750_));
  OR2_X1    g549(.A1(new_n663_), .A2(G64gat), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n746_), .B2(new_n751_), .ZN(G1333gat));
  OAI21_X1  g551(.A(G71gat), .B1(new_n743_), .B2(new_n397_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT49), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n397_), .A2(G71gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n754_), .B1(new_n746_), .B2(new_n755_), .ZN(G1334gat));
  OAI21_X1  g555(.A(G78gat), .B1(new_n743_), .B2(new_n679_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT50), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n381_), .A2(new_n373_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n758_), .B1(new_n746_), .B2(new_n759_), .ZN(G1335gat));
  NAND2_X1  g559(.A1(new_n745_), .A2(new_n706_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(G85gat), .B1(new_n762_), .B2(new_n701_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n742_), .A2(new_n466_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT111), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n765_), .B1(new_n694_), .B2(new_n697_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n766_), .A2(KEYINPUT112), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(KEYINPUT112), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n339_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n763_), .B1(new_n769_), .B2(new_n770_), .ZN(G1336gat));
  NAND3_X1  g570(.A1(new_n762_), .A2(new_n489_), .A3(new_n423_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n767_), .A2(new_n768_), .A3(new_n663_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n772_), .B1(new_n773_), .B2(new_n489_), .ZN(G1337gat));
  NOR2_X1   g573(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n766_), .A2(new_n398_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(G99gat), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n762_), .A2(new_n482_), .A3(new_n398_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n775_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  AND2_X1   g578(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n779_), .B(new_n780_), .ZN(G1338gat));
  NAND3_X1  g580(.A1(new_n762_), .A2(new_n483_), .A3(new_n381_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n766_), .A2(new_n381_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n784_), .B2(G106gat), .ZN(new_n785_));
  AOI211_X1 g584(.A(KEYINPUT52), .B(new_n372_), .C1(new_n766_), .C2(new_n381_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n782_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT53), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT53), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n789_), .B(new_n782_), .C1(new_n785_), .C2(new_n786_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(G1339gat));
  INV_X1    g590(.A(KEYINPUT119), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n632_), .A2(new_n637_), .A3(new_n609_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n794_), .B1(new_n608_), .B2(new_n598_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n594_), .A2(new_n599_), .A3(KEYINPUT55), .A4(new_n600_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n596_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n603_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n795_), .A2(new_n796_), .A3(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n588_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT56), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n799_), .A2(KEYINPUT56), .A3(new_n588_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n793_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n617_), .A2(KEYINPUT81), .A3(new_n618_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n625_), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n805_), .A2(new_n619_), .A3(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT115), .B1(new_n807_), .B2(new_n629_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n620_), .A2(new_n621_), .A3(new_n625_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(new_n810_), .A3(new_n634_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n623_), .A2(new_n618_), .A3(new_n806_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n808_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT116), .B1(new_n813_), .B2(new_n636_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n813_), .A2(KEYINPUT116), .A3(new_n636_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n611_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n692_), .B1(new_n804_), .B2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT57), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT57), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n820_), .B(new_n692_), .C1(new_n804_), .C2(new_n817_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n802_), .A2(new_n803_), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n813_), .A2(KEYINPUT116), .A3(new_n636_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n609_), .B1(new_n824_), .B2(new_n814_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  OAI211_X1 g626(.A(KEYINPUT117), .B(new_n609_), .C1(new_n824_), .C2(new_n814_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n823_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n696_), .B1(new_n829_), .B2(KEYINPUT58), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT58), .ZN(new_n831_));
  AOI211_X1 g630(.A(new_n831_), .B(new_n823_), .C1(new_n827_), .C2(new_n828_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n822_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n465_), .B1(new_n833_), .B2(KEYINPUT118), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n822_), .B(new_n835_), .C1(new_n830_), .C2(new_n832_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n615_), .A2(new_n741_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n693_), .A2(new_n465_), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT54), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n582_), .A2(new_n840_), .A3(new_n841_), .A4(new_n837_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n839_), .A2(new_n842_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n693_), .A2(new_n841_), .A3(new_n465_), .A4(new_n837_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT114), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n834_), .A2(new_n836_), .B1(new_n843_), .B2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n424_), .A2(new_n701_), .A3(new_n398_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n792_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n833_), .A2(KEYINPUT118), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n849_), .A2(new_n466_), .A3(new_n836_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n845_), .A2(new_n839_), .A3(new_n842_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n847_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(KEYINPUT119), .A3(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n848_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(G113gat), .B1(new_n856_), .B2(new_n741_), .ZN(new_n857_));
  OAI21_X1  g656(.A(KEYINPUT59), .B1(new_n846_), .B2(new_n847_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n833_), .A2(new_n466_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n851_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n861_), .A3(new_n853_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n858_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n741_), .A2(G113gat), .ZN(new_n865_));
  XOR2_X1   g664(.A(new_n865_), .B(KEYINPUT120), .Z(new_n866_));
  AOI21_X1  g665(.A(new_n857_), .B1(new_n864_), .B2(new_n866_), .ZN(G1340gat));
  NAND3_X1  g666(.A1(new_n864_), .A2(KEYINPUT121), .A3(new_n615_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(new_n863_), .B2(new_n740_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n868_), .A2(G120gat), .A3(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(G120gat), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n872_), .B1(new_n740_), .B2(KEYINPUT60), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(KEYINPUT60), .B2(new_n872_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n871_), .B1(new_n855_), .B2(new_n874_), .ZN(G1341gat));
  NAND3_X1  g674(.A1(new_n864_), .A2(G127gat), .A3(new_n465_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n848_), .A2(new_n854_), .A3(new_n465_), .ZN(new_n877_));
  INV_X1    g676(.A(G127gat), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n877_), .A2(KEYINPUT122), .A3(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(KEYINPUT122), .B1(new_n877_), .B2(new_n878_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n876_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(KEYINPUT123), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT123), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n883_), .B(new_n876_), .C1(new_n879_), .C2(new_n880_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n882_), .A2(new_n884_), .ZN(G1342gat));
  OAI21_X1  g684(.A(G134gat), .B1(new_n863_), .B2(new_n693_), .ZN(new_n886_));
  OR2_X1    g685(.A1(new_n692_), .A2(G134gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n855_), .B2(new_n887_), .ZN(G1343gat));
  NOR3_X1   g687(.A1(new_n846_), .A2(new_n679_), .A3(new_n398_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n423_), .A2(new_n339_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n741_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g693(.A1(new_n891_), .A2(new_n740_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT124), .B(G148gat), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1345gat));
  NOR2_X1   g696(.A1(new_n891_), .A2(new_n466_), .ZN(new_n898_));
  XOR2_X1   g697(.A(KEYINPUT61), .B(G155gat), .Z(new_n899_));
  XNOR2_X1  g698(.A(new_n898_), .B(new_n899_), .ZN(G1346gat));
  OR3_X1    g699(.A1(new_n891_), .A2(G162gat), .A3(new_n692_), .ZN(new_n901_));
  OAI21_X1  g700(.A(G162gat), .B1(new_n891_), .B2(new_n693_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1347gat));
  NOR2_X1   g702(.A1(new_n663_), .A2(new_n701_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n398_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n905_), .A2(new_n381_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n860_), .A2(new_n906_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(new_n638_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n908_), .A2(new_n247_), .ZN(new_n909_));
  AOI22_X1  g708(.A1(new_n909_), .A2(KEYINPUT62), .B1(new_n249_), .B2(new_n908_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n910_), .B1(KEYINPUT62), .B2(new_n909_), .ZN(G1348gat));
  INV_X1    g710(.A(new_n907_), .ZN(new_n912_));
  AOI21_X1  g711(.A(G176gat), .B1(new_n912_), .B2(new_n615_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n846_), .A2(new_n381_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n905_), .A2(new_n245_), .A3(new_n740_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n913_), .B1(new_n914_), .B2(new_n915_), .ZN(G1349gat));
  NAND3_X1  g715(.A1(new_n912_), .A2(new_n465_), .A3(new_n229_), .ZN(new_n917_));
  XOR2_X1   g716(.A(new_n917_), .B(KEYINPUT125), .Z(new_n918_));
  NOR2_X1   g717(.A1(new_n905_), .A2(new_n466_), .ZN(new_n919_));
  AOI21_X1  g718(.A(G183gat), .B1(new_n914_), .B2(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n918_), .A2(new_n920_), .ZN(G1350gat));
  OAI21_X1  g720(.A(G190gat), .B1(new_n907_), .B2(new_n693_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n579_), .A2(new_n259_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(KEYINPUT126), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n922_), .B1(new_n907_), .B2(new_n924_), .ZN(G1351gat));
  NAND2_X1  g724(.A1(new_n889_), .A2(new_n904_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n926_), .A2(new_n638_), .ZN(new_n927_));
  OR2_X1    g726(.A1(new_n205_), .A2(KEYINPUT127), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n205_), .A2(KEYINPUT127), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n927_), .B1(new_n928_), .B2(new_n929_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n930_), .B1(new_n927_), .B2(new_n929_), .ZN(G1352gat));
  NOR2_X1   g730(.A1(new_n926_), .A2(new_n740_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(new_n207_), .ZN(G1353gat));
  INV_X1    g732(.A(new_n926_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(new_n465_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n936_));
  AND2_X1   g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  NOR3_X1   g736(.A1(new_n935_), .A2(new_n936_), .A3(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n938_), .B1(new_n935_), .B2(new_n936_), .ZN(G1354gat));
  OR3_X1    g738(.A1(new_n926_), .A2(G218gat), .A3(new_n692_), .ZN(new_n940_));
  OAI21_X1  g739(.A(G218gat), .B1(new_n926_), .B2(new_n693_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(G1355gat));
endmodule


