//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 0 0 0 1 0 0 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n909_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_, new_n939_;
  INV_X1    g000(.A(KEYINPUT67), .ZN(new_n202_));
  INV_X1    g001(.A(G85gat), .ZN(new_n203_));
  INV_X1    g002(.A(G92gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G85gat), .A2(G92gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NOR3_X1   g008(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT6), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  AOI211_X1 g015(.A(KEYINPUT8), .B(new_n207_), .C1(new_n211_), .C2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n214_), .B1(G99gat), .B2(G106gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n218_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n213_), .A2(new_n215_), .A3(KEYINPUT66), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(new_n222_), .A3(new_n211_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n207_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n217_), .B1(new_n225_), .B2(KEYINPUT8), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT9), .ZN(new_n227_));
  AND2_X1   g026(.A1(G85gat), .A2(G92gat), .ZN(new_n228_));
  OAI211_X1 g027(.A(new_n205_), .B(new_n227_), .C1(new_n228_), .C2(KEYINPUT64), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n205_), .A2(new_n230_), .A3(KEYINPUT9), .A4(new_n206_), .ZN(new_n231_));
  OR2_X1    g030(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n232_));
  INV_X1    g031(.A(G106gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n229_), .A2(new_n231_), .A3(new_n216_), .A4(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n202_), .B1(new_n226_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n236_), .A2(KEYINPUT65), .ZN(new_n240_));
  AND2_X1   g039(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n241_));
  NOR2_X1   g040(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  AOI22_X1  g042(.A1(new_n243_), .A2(new_n233_), .B1(new_n213_), .B2(new_n215_), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n244_), .A2(new_n237_), .A3(new_n229_), .A4(new_n231_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n240_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT8), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n247_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n246_), .B(KEYINPUT67), .C1(new_n248_), .C2(new_n217_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT12), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G57gat), .B(G64gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G71gat), .B(G78gat), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n251_), .A2(new_n252_), .A3(KEYINPUT11), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(KEYINPUT11), .ZN(new_n254_));
  INV_X1    g053(.A(new_n252_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n251_), .A2(KEYINPUT11), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n253_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT68), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  OAI211_X1 g059(.A(KEYINPUT68), .B(new_n253_), .C1(new_n256_), .C2(new_n257_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n250_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n239_), .A2(new_n249_), .A3(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT69), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n246_), .B1(new_n248_), .B2(new_n217_), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n256_), .A2(new_n257_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(new_n253_), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(new_n250_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n239_), .A2(new_n269_), .A3(new_n249_), .A4(new_n262_), .ZN(new_n270_));
  AND2_X1   g069(.A1(G230gat), .A2(G233gat), .ZN(new_n271_));
  INV_X1    g070(.A(new_n265_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n271_), .B1(new_n272_), .B2(new_n258_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n264_), .A2(new_n268_), .A3(new_n270_), .A4(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n258_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n267_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(new_n271_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n274_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G120gat), .B(G148gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT5), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G176gat), .B(G204gat), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n280_), .B(new_n281_), .Z(new_n282_));
  NAND2_X1  g081(.A1(new_n278_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n284_));
  INV_X1    g083(.A(new_n282_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n274_), .A2(new_n277_), .A3(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n283_), .A2(new_n284_), .A3(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n278_), .A2(KEYINPUT70), .A3(new_n282_), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT13), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(G183gat), .B(G211gat), .Z(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT79), .ZN(new_n293_));
  XOR2_X1   g092(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G127gat), .B(G155gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n297_), .A2(KEYINPUT17), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(KEYINPUT17), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G15gat), .B(G22gat), .ZN(new_n300_));
  INV_X1    g099(.A(G1gat), .ZN(new_n301_));
  INV_X1    g100(.A(G8gat), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT14), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n300_), .A2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G1gat), .B(G8gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G231gat), .A2(G233gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(new_n258_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n298_), .A2(new_n299_), .A3(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n310_), .B(KEYINPUT81), .Z(new_n311_));
  NAND2_X1  g110(.A1(new_n260_), .A2(new_n261_), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n308_), .B(new_n312_), .Z(new_n313_));
  AOI21_X1  g112(.A(new_n313_), .B1(KEYINPUT80), .B2(new_n299_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n314_), .B1(KEYINPUT80), .B2(new_n299_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n311_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G29gat), .B(G36gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G43gat), .B(G50gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT15), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n239_), .A2(new_n249_), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(KEYINPUT71), .B(KEYINPUT34), .Z(new_n323_));
  NAND2_X1  g122(.A1(G232gat), .A2(G233gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT35), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n326_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n319_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n328_), .B1(new_n265_), .B2(new_n329_), .ZN(new_n330_));
  NOR3_X1   g129(.A1(new_n322_), .A2(new_n327_), .A3(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  XOR2_X1   g131(.A(G190gat), .B(G218gat), .Z(new_n333_));
  XNOR2_X1  g132(.A(G134gat), .B(G162gat), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n334_), .ZN(new_n336_));
  AOI21_X1  g135(.A(KEYINPUT36), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n330_), .A2(KEYINPUT72), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT72), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n341_), .B(new_n328_), .C1(new_n265_), .C2(new_n329_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n340_), .A2(new_n321_), .A3(new_n342_), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n343_), .A2(KEYINPUT73), .A3(new_n327_), .ZN(new_n344_));
  AOI21_X1  g143(.A(KEYINPUT73), .B1(new_n343_), .B2(new_n327_), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n332_), .B(new_n339_), .C1(new_n344_), .C2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT37), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n343_), .A2(new_n327_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT73), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n343_), .A2(KEYINPUT73), .A3(new_n327_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n331_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n335_), .A2(new_n336_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT36), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n346_), .B(new_n347_), .C1(new_n352_), .C2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT77), .B1(new_n352_), .B2(new_n355_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n352_), .A2(new_n359_), .A3(new_n339_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n346_), .A2(KEYINPUT76), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n332_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT77), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(new_n363_), .A3(new_n354_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n358_), .A2(new_n360_), .A3(new_n361_), .A4(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n357_), .B1(new_n365_), .B2(KEYINPUT37), .ZN(new_n366_));
  NOR3_X1   g165(.A1(new_n291_), .A2(new_n316_), .A3(new_n366_), .ZN(new_n367_));
  OR2_X1    g166(.A1(new_n367_), .A2(KEYINPUT82), .ZN(new_n368_));
  NOR3_X1   g167(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G183gat), .A2(G190gat), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT23), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT84), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n374_), .B1(G169gat), .B2(G176gat), .ZN(new_n375_));
  AOI211_X1 g174(.A(new_n369_), .B(new_n372_), .C1(new_n373_), .C2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT25), .B(G183gat), .ZN(new_n377_));
  XOR2_X1   g176(.A(KEYINPUT83), .B(G190gat), .Z(new_n378_));
  INV_X1    g177(.A(KEYINPUT26), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n377_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n376_), .B(new_n382_), .C1(new_n373_), .C2(new_n375_), .ZN(new_n383_));
  INV_X1    g182(.A(G183gat), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n372_), .B1(new_n384_), .B2(new_n378_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n386_));
  INV_X1    g185(.A(G169gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n385_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n383_), .A2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G71gat), .B(G99gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(G43gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n390_), .B(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G227gat), .A2(G233gat), .ZN(new_n394_));
  INV_X1    g193(.A(G15gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT30), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT31), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n393_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT85), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G127gat), .B(G134gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G113gat), .B(G120gat), .ZN(new_n402_));
  XOR2_X1   g201(.A(new_n401_), .B(new_n402_), .Z(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n400_), .B(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT101), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G155gat), .A2(G162gat), .ZN(new_n407_));
  NOR2_X1   g206(.A1(G155gat), .A2(G162gat), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n410_));
  OR2_X1    g209(.A1(new_n410_), .A2(KEYINPUT86), .ZN(new_n411_));
  AND2_X1   g210(.A1(G141gat), .A2(G148gat), .ZN(new_n412_));
  NOR2_X1   g211(.A1(G141gat), .A2(G148gat), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT3), .ZN(new_n414_));
  AOI22_X1  g213(.A1(KEYINPUT2), .A2(new_n412_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n410_), .A2(KEYINPUT86), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n411_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT87), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n407_), .B(new_n409_), .C1(new_n417_), .C2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n408_), .B1(KEYINPUT1), .B2(new_n407_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n421_), .B1(KEYINPUT1), .B2(new_n407_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n412_), .A2(new_n413_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n420_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT88), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT88), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n425_), .A2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n427_), .A2(new_n429_), .A3(new_n403_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n426_), .A2(new_n404_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n430_), .A2(KEYINPUT4), .A3(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n430_), .A2(KEYINPUT4), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G225gat), .A2(G233gat), .ZN(new_n434_));
  XOR2_X1   g233(.A(new_n434_), .B(KEYINPUT94), .Z(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n433_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n430_), .A2(new_n431_), .A3(new_n434_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT96), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT96), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n430_), .A2(new_n440_), .A3(new_n431_), .A4(new_n434_), .ZN(new_n441_));
  AOI22_X1  g240(.A1(new_n432_), .A2(new_n437_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(G1gat), .B(G29gat), .Z(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT95), .B(G85gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT0), .B(G57gat), .ZN(new_n446_));
  XOR2_X1   g245(.A(new_n445_), .B(new_n446_), .Z(new_n447_));
  NOR2_X1   g246(.A1(new_n442_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n437_), .A2(new_n432_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n439_), .A2(new_n441_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(new_n450_), .A3(new_n447_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n406_), .B1(new_n448_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n449_), .A2(new_n450_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n447_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n456_), .A2(KEYINPUT101), .A3(new_n451_), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n453_), .A2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G211gat), .B(G218gat), .ZN(new_n459_));
  INV_X1    g258(.A(G204gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(G197gat), .ZN(new_n461_));
  INV_X1    g260(.A(G197gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(G204gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n461_), .A2(new_n463_), .A3(KEYINPUT90), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT21), .B1(new_n461_), .B2(KEYINPUT90), .ZN(new_n466_));
  OAI221_X1 g265(.A(new_n459_), .B1(KEYINPUT21), .B2(new_n464_), .C1(new_n465_), .C2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n464_), .A2(KEYINPUT21), .ZN(new_n468_));
  OR2_X1    g267(.A1(new_n468_), .A2(new_n459_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT29), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n470_), .B1(new_n426_), .B2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n472_), .A2(G228gat), .A3(G233gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n427_), .A2(new_n429_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n474_), .A2(new_n471_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G228gat), .A2(G233gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n470_), .A2(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n473_), .B1(new_n475_), .B2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G78gat), .B(G106gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n479_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n481_), .B(new_n473_), .C1(new_n475_), .C2(new_n477_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n474_), .A2(new_n471_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G22gat), .B(G50gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n484_), .B(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT91), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n490_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n483_), .B1(new_n489_), .B2(new_n491_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n480_), .A2(new_n488_), .A3(new_n490_), .A4(new_n482_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT20), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n370_), .B(KEYINPUT23), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n497_), .B1(G183gat), .B2(G190gat), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n388_), .B1(new_n498_), .B2(KEYINPUT92), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT92), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n497_), .B(new_n500_), .C1(G183gat), .C2(G190gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n375_), .A2(new_n369_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT26), .B(G190gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n377_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n503_), .A2(new_n497_), .A3(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n502_), .A2(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n496_), .B1(new_n507_), .B2(new_n470_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n470_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n383_), .A2(new_n509_), .A3(new_n389_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G226gat), .A2(G233gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT19), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G8gat), .B(G36gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT18), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G64gat), .B(G92gat), .ZN(new_n517_));
  XOR2_X1   g316(.A(new_n516_), .B(new_n517_), .Z(new_n518_));
  NAND2_X1  g317(.A1(new_n390_), .A2(new_n470_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n513_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n509_), .A2(new_n502_), .A3(new_n506_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n519_), .A2(KEYINPUT20), .A3(new_n520_), .A4(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n514_), .A2(new_n518_), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n518_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n520_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n521_), .A2(KEYINPUT20), .A3(new_n520_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n509_), .B1(new_n383_), .B2(new_n389_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n524_), .B1(new_n525_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n523_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT27), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n511_), .A2(new_n513_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT100), .B(KEYINPUT20), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n521_), .A2(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n520_), .B1(new_n535_), .B2(new_n519_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n533_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n518_), .B(KEYINPUT102), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  OAI211_X1 g338(.A(KEYINPUT27), .B(new_n523_), .C1(new_n537_), .C2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n532_), .A2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n495_), .A2(new_n541_), .ZN(new_n542_));
  AND3_X1   g341(.A1(new_n405_), .A2(new_n458_), .A3(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n494_), .A2(new_n541_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n458_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n518_), .A2(KEYINPUT32), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n514_), .A2(new_n522_), .A3(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n547_), .B1(new_n537_), .B2(new_n546_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n548_), .B1(new_n456_), .B2(new_n451_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n442_), .A2(KEYINPUT33), .A3(new_n447_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT93), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n523_), .A2(new_n529_), .A3(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n551_), .B1(new_n523_), .B2(new_n529_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n434_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n433_), .A2(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n447_), .B1(new_n556_), .B2(new_n432_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n430_), .A2(new_n431_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n436_), .B1(new_n558_), .B2(KEYINPUT98), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n559_), .B1(KEYINPUT98), .B2(new_n558_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT99), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n557_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n561_), .B1(new_n557_), .B2(new_n560_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n550_), .B(new_n554_), .C1(new_n562_), .C2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT97), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT33), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n451_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n566_), .B1(new_n451_), .B2(new_n567_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n549_), .B1(new_n565_), .B2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n545_), .B1(new_n571_), .B2(new_n495_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n405_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n543_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n320_), .A2(new_n306_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G229gat), .A2(G233gat), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n306_), .A2(new_n329_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n575_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n306_), .B(new_n329_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n579_), .A2(G229gat), .A3(G233gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G113gat), .B(G141gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G169gat), .B(G197gat), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n582_), .B(new_n583_), .Z(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n581_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n578_), .A2(new_n580_), .A3(new_n584_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n574_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n367_), .A2(KEYINPUT82), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n368_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n591_), .A2(KEYINPUT103), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(KEYINPUT103), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT38), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n453_), .A2(new_n457_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(new_n301_), .ZN(new_n597_));
  OR3_X1    g396(.A1(new_n594_), .A2(new_n595_), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n316_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n346_), .B1(new_n352_), .B2(new_n355_), .ZN(new_n600_));
  NOR3_X1   g399(.A1(new_n564_), .A2(new_n569_), .A3(new_n568_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n494_), .B1(new_n601_), .B2(new_n549_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n405_), .B1(new_n602_), .B2(new_n545_), .ZN(new_n603_));
  OAI211_X1 g402(.A(new_n599_), .B(new_n600_), .C1(new_n603_), .C2(new_n543_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n291_), .A2(new_n588_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(G1gat), .B1(new_n608_), .B2(new_n458_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n595_), .B1(new_n594_), .B2(new_n597_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n598_), .A2(new_n609_), .A3(new_n610_), .ZN(G1324gat));
  INV_X1    g410(.A(new_n600_), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n574_), .A2(new_n316_), .A3(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n613_), .A2(new_n541_), .A3(new_n605_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(G8gat), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT39), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT39), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n614_), .A2(new_n617_), .A3(G8gat), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n541_), .A2(new_n302_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n619_), .B1(new_n594_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT40), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n619_), .B(KEYINPUT40), .C1(new_n594_), .C2(new_n620_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1325gat));
  AOI21_X1  g424(.A(new_n395_), .B1(new_n607_), .B2(new_n405_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT41), .ZN(new_n627_));
  INV_X1    g426(.A(new_n591_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n628_), .A2(new_n395_), .A3(new_n405_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(G1326gat));
  INV_X1    g429(.A(KEYINPUT42), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n607_), .A2(new_n495_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n631_), .B1(new_n632_), .B2(G22gat), .ZN(new_n633_));
  INV_X1    g432(.A(G22gat), .ZN(new_n634_));
  AOI211_X1 g433(.A(KEYINPUT42), .B(new_n634_), .C1(new_n607_), .C2(new_n495_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n494_), .A2(G22gat), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT104), .Z(new_n637_));
  OAI22_X1  g436(.A1(new_n633_), .A2(new_n635_), .B1(new_n591_), .B2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT105), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(G1327gat));
  INV_X1    g439(.A(new_n366_), .ZN(new_n641_));
  OAI21_X1  g440(.A(KEYINPUT43), .B1(new_n574_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT43), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n643_), .B(new_n366_), .C1(new_n603_), .C2(new_n543_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n605_), .A2(new_n316_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT44), .B1(new_n645_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n649_));
  AOI211_X1 g448(.A(new_n649_), .B(new_n646_), .C1(new_n642_), .C2(new_n644_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n596_), .A2(G29gat), .ZN(new_n652_));
  INV_X1    g451(.A(G29gat), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n562_), .A2(new_n563_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n554_), .A2(new_n550_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n570_), .A2(new_n654_), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n549_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n495_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n596_), .A2(new_n494_), .A3(new_n541_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n573_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n543_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n316_), .A2(new_n612_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n663_), .A2(new_n605_), .A3(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT106), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n663_), .A2(KEYINPUT106), .A3(new_n605_), .A4(new_n665_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(new_n596_), .A3(new_n669_), .ZN(new_n670_));
  AOI22_X1  g469(.A1(new_n651_), .A2(new_n652_), .B1(new_n653_), .B2(new_n670_), .ZN(G1328gat));
  INV_X1    g470(.A(KEYINPUT46), .ZN(new_n672_));
  INV_X1    g471(.A(G36gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n673_), .B1(new_n651_), .B2(new_n541_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n541_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n675_), .A2(G36gat), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n668_), .A2(new_n669_), .A3(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n678_), .B(KEYINPUT108), .Z(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n677_), .B(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n672_), .B1(new_n674_), .B2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n677_), .B(new_n679_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n648_), .A2(new_n650_), .A3(new_n675_), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n683_), .B(KEYINPUT46), .C1(new_n673_), .C2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n682_), .A2(new_n685_), .ZN(G1329gat));
  INV_X1    g485(.A(G43gat), .ZN(new_n687_));
  NOR4_X1   g486(.A1(new_n648_), .A2(new_n650_), .A3(new_n687_), .A4(new_n573_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n668_), .A2(new_n405_), .A3(new_n669_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(new_n687_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(KEYINPUT47), .B1(new_n688_), .B2(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n651_), .A2(G43gat), .A3(new_n405_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT47), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(new_n694_), .A3(new_n690_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n692_), .A2(new_n695_), .ZN(G1330gat));
  INV_X1    g495(.A(KEYINPUT109), .ZN(new_n697_));
  INV_X1    g496(.A(G50gat), .ZN(new_n698_));
  NOR4_X1   g497(.A1(new_n648_), .A2(new_n650_), .A3(new_n698_), .A4(new_n494_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n668_), .A2(new_n495_), .A3(new_n669_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n698_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n697_), .B1(new_n699_), .B2(new_n702_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n651_), .A2(G50gat), .A3(new_n495_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n704_), .A2(KEYINPUT109), .A3(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(G1331gat));
  NAND2_X1  g505(.A1(new_n291_), .A2(new_n588_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n604_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G57gat), .B1(new_n709_), .B2(new_n458_), .ZN(new_n710_));
  NOR4_X1   g509(.A1(new_n574_), .A2(new_n316_), .A3(new_n707_), .A4(new_n366_), .ZN(new_n711_));
  INV_X1    g510(.A(G57gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n711_), .A2(new_n712_), .A3(new_n596_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n710_), .A2(new_n713_), .ZN(G1332gat));
  INV_X1    g513(.A(G64gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n708_), .B2(new_n541_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT48), .Z(new_n717_));
  NAND3_X1  g516(.A1(new_n711_), .A2(new_n715_), .A3(new_n541_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1333gat));
  INV_X1    g518(.A(G71gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n720_), .B1(new_n708_), .B2(new_n405_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT49), .Z(new_n722_));
  NAND3_X1  g521(.A1(new_n711_), .A2(new_n720_), .A3(new_n405_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1334gat));
  NOR2_X1   g523(.A1(new_n494_), .A2(G78gat), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT110), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n711_), .A2(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(G78gat), .B1(new_n709_), .B2(new_n494_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n728_), .A2(KEYINPUT50), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n728_), .A2(KEYINPUT50), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n727_), .B1(new_n729_), .B2(new_n730_), .ZN(G1335gat));
  NOR3_X1   g530(.A1(new_n574_), .A2(new_n664_), .A3(new_n707_), .ZN(new_n732_));
  AOI21_X1  g531(.A(G85gat), .B1(new_n732_), .B2(new_n596_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n645_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n707_), .A2(new_n599_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n734_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n596_), .A2(G85gat), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT111), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n733_), .B1(new_n737_), .B2(new_n739_), .ZN(G1336gat));
  NAND3_X1  g539(.A1(new_n732_), .A2(new_n204_), .A3(new_n541_), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n734_), .A2(new_n675_), .A3(new_n736_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n741_), .B1(new_n742_), .B2(new_n204_), .ZN(G1337gat));
  NAND3_X1  g542(.A1(new_n732_), .A2(new_n243_), .A3(new_n405_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n734_), .A2(new_n573_), .A3(new_n736_), .ZN(new_n745_));
  INV_X1    g544(.A(G99gat), .ZN(new_n746_));
  OAI211_X1 g545(.A(KEYINPUT112), .B(new_n744_), .C1(new_n745_), .C2(new_n746_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g547(.A1(new_n732_), .A2(new_n233_), .A3(new_n495_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n645_), .A2(new_n495_), .A3(new_n735_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n750_), .A2(new_n751_), .A3(G106gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n750_), .B2(G106gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n749_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(KEYINPUT53), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT53), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n756_), .B(new_n749_), .C1(new_n752_), .C2(new_n753_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1339gat));
  INV_X1    g557(.A(KEYINPUT118), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n366_), .A2(new_n316_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n760_), .A2(new_n290_), .A3(new_n588_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n760_), .A2(new_n290_), .A3(new_n588_), .A4(new_n762_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT116), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT115), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n575_), .A2(new_n577_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT114), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n576_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n575_), .A2(KEYINPUT114), .A3(new_n577_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n579_), .A2(new_n576_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n585_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n768_), .B(new_n587_), .C1(new_n773_), .C2(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n587_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT115), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n776_), .A2(new_n779_), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n287_), .A2(new_n288_), .A3(new_n780_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n264_), .A2(new_n275_), .A3(new_n268_), .A4(new_n270_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n271_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n274_), .A2(new_n784_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n270_), .A2(new_n268_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n786_), .A2(KEYINPUT55), .A3(new_n264_), .A4(new_n273_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n783_), .A2(new_n785_), .A3(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n282_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT56), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n788_), .A2(KEYINPUT56), .A3(new_n282_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n588_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n794_), .A2(new_n286_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n781_), .B1(new_n793_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n600_), .A2(KEYINPUT57), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n767_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n788_), .A2(KEYINPUT56), .A3(new_n282_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT56), .B1(new_n788_), .B2(new_n282_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n795_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n287_), .A2(new_n288_), .A3(new_n780_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n797_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n803_), .A2(KEYINPUT116), .A3(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n798_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n807_), .B1(new_n796_), .B2(new_n612_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n780_), .A2(new_n286_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n793_), .A2(KEYINPUT58), .A3(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT58), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n366_), .A2(new_n810_), .A3(new_n813_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n806_), .A2(KEYINPUT117), .A3(new_n808_), .A4(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT116), .B1(new_n803_), .B2(new_n804_), .ZN(new_n816_));
  AOI211_X1 g615(.A(new_n767_), .B(new_n797_), .C1(new_n801_), .C2(new_n802_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n808_), .B(new_n814_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT117), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n599_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n766_), .B1(new_n815_), .B2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n405_), .A2(new_n542_), .A3(new_n596_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n759_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n818_), .A2(new_n819_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n824_), .A2(new_n815_), .A3(new_n316_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n764_), .A2(new_n765_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n822_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n827_), .A2(KEYINPUT118), .A3(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(G113gat), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n823_), .A2(new_n829_), .A3(new_n830_), .A4(new_n794_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n822_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n818_), .A2(new_n316_), .ZN(new_n834_));
  OR2_X1    g633(.A1(new_n834_), .A2(new_n766_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n822_), .A2(KEYINPUT59), .ZN(new_n836_));
  AOI22_X1  g635(.A1(new_n833_), .A2(KEYINPUT59), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n794_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n831_), .B1(new_n839_), .B2(new_n830_), .ZN(G1340gat));
  OAI21_X1  g639(.A(new_n836_), .B1(new_n834_), .B2(new_n766_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT59), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n291_), .B(new_n841_), .C1(new_n832_), .C2(new_n842_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(KEYINPUT119), .B(G120gat), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(new_n846_));
  OR2_X1    g645(.A1(new_n844_), .A2(KEYINPUT60), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n844_), .B1(new_n290_), .B2(KEYINPUT60), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n823_), .A2(new_n829_), .A3(new_n847_), .A4(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n846_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(KEYINPUT120), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n846_), .A2(new_n852_), .A3(new_n849_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(G1341gat));
  NAND2_X1  g653(.A1(new_n599_), .A2(G127gat), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(KEYINPUT121), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n823_), .A2(new_n599_), .A3(new_n829_), .ZN(new_n857_));
  INV_X1    g656(.A(G127gat), .ZN(new_n858_));
  AOI22_X1  g657(.A1(new_n837_), .A2(new_n856_), .B1(new_n857_), .B2(new_n858_), .ZN(G1342gat));
  OAI211_X1 g658(.A(new_n366_), .B(new_n841_), .C1(new_n832_), .C2(new_n842_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(G134gat), .ZN(new_n861_));
  INV_X1    g660(.A(G134gat), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n823_), .A2(new_n829_), .A3(new_n862_), .A4(new_n612_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n861_), .A2(KEYINPUT122), .A3(new_n863_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(G1343gat));
  NAND2_X1  g667(.A1(new_n596_), .A2(new_n544_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n821_), .A2(new_n405_), .A3(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n794_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n291_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g673(.A(new_n869_), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n827_), .A2(new_n599_), .A3(new_n573_), .A4(new_n875_), .ZN(new_n876_));
  OR2_X1    g675(.A1(new_n876_), .A2(KEYINPUT123), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(KEYINPUT123), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(KEYINPUT61), .B(G155gat), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n877_), .A2(new_n878_), .A3(new_n880_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1346gat));
  INV_X1    g683(.A(G162gat), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n870_), .A2(new_n885_), .A3(new_n612_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n870_), .A2(new_n366_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(new_n885_), .ZN(G1347gat));
  NOR2_X1   g687(.A1(new_n573_), .A2(new_n596_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n541_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n494_), .B(new_n891_), .C1(new_n834_), .C2(new_n766_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(new_n794_), .ZN(new_n894_));
  OAI21_X1  g693(.A(KEYINPUT62), .B1(new_n894_), .B2(KEYINPUT22), .ZN(new_n895_));
  OAI21_X1  g694(.A(G169gat), .B1(new_n894_), .B2(KEYINPUT62), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n897_), .B1(new_n387_), .B2(new_n895_), .ZN(G1348gat));
  AOI21_X1  g697(.A(G176gat), .B1(new_n893_), .B2(new_n291_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n821_), .A2(new_n495_), .ZN(new_n900_));
  AND3_X1   g699(.A1(new_n891_), .A2(G176gat), .A3(new_n291_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n899_), .B1(new_n900_), .B2(new_n901_), .ZN(G1349gat));
  NAND2_X1  g701(.A1(new_n835_), .A2(new_n494_), .ZN(new_n903_));
  NOR4_X1   g702(.A1(new_n903_), .A2(new_n316_), .A3(new_n377_), .A4(new_n890_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n890_), .A2(new_n316_), .ZN(new_n905_));
  AOI21_X1  g704(.A(G183gat), .B1(new_n900_), .B2(new_n905_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n904_), .A2(new_n906_), .ZN(G1350gat));
  OAI21_X1  g706(.A(G190gat), .B1(new_n892_), .B2(new_n641_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n612_), .A2(new_n504_), .ZN(new_n909_));
  XOR2_X1   g708(.A(new_n909_), .B(KEYINPUT124), .Z(new_n910_));
  OAI21_X1  g709(.A(new_n908_), .B1(new_n892_), .B2(new_n910_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(KEYINPUT125), .ZN(G1351gat));
  NOR3_X1   g711(.A1(new_n596_), .A2(new_n494_), .A3(new_n675_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n827_), .A2(new_n573_), .A3(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT126), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  NAND4_X1  g715(.A1(new_n827_), .A2(KEYINPUT126), .A3(new_n573_), .A4(new_n913_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  AOI21_X1  g717(.A(G197gat), .B1(new_n918_), .B2(new_n794_), .ZN(new_n919_));
  AOI211_X1 g718(.A(new_n462_), .B(new_n588_), .C1(new_n916_), .C2(new_n917_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n919_), .A2(new_n920_), .ZN(G1352gat));
  NOR2_X1   g720(.A1(new_n821_), .A2(new_n405_), .ZN(new_n922_));
  AOI21_X1  g721(.A(KEYINPUT126), .B1(new_n922_), .B2(new_n913_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n917_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n291_), .B1(new_n923_), .B2(new_n924_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(G204gat), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n918_), .A2(new_n460_), .A3(new_n291_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(G1353gat));
  AOI21_X1  g727(.A(new_n316_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n929_), .B1(new_n923_), .B2(new_n924_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(KEYINPUT127), .ZN(new_n932_));
  INV_X1    g731(.A(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n930_), .A2(new_n933_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n918_), .A2(new_n929_), .A3(new_n932_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(G1354gat));
  INV_X1    g735(.A(G218gat), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n918_), .A2(new_n937_), .A3(new_n612_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n641_), .B1(new_n916_), .B2(new_n917_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n938_), .B1(new_n937_), .B2(new_n939_), .ZN(G1355gat));
endmodule


