//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 1 1 1 1 0 0 0 1 0 0 0 0 0 1 1 0 0 1 0 0 1 1 0 0 0 1 1 1 1 1 0 1 0 0 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n632_, new_n633_, new_n634_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n799_, new_n800_, new_n801_,
    new_n803_, new_n804_, new_n805_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n821_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n860_, new_n861_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_;
  XOR2_X1   g000(.A(G127gat), .B(G155gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT16), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G183gat), .B(G211gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT17), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT75), .B(G15gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(G22gat), .ZN(new_n209_));
  INV_X1    g008(.A(G1gat), .ZN(new_n210_));
  INV_X1    g009(.A(G8gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT14), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  XOR2_X1   g012(.A(G1gat), .B(G8gat), .Z(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n209_), .A2(new_n214_), .A3(new_n212_), .ZN(new_n217_));
  AND2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G231gat), .A2(G233gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n218_), .B(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G57gat), .B(G64gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT67), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n221_), .A2(new_n222_), .A3(KEYINPUT11), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n222_), .B1(new_n221_), .B2(KEYINPUT11), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n221_), .A2(KEYINPUT11), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G71gat), .B(G78gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n225_), .A2(new_n228_), .ZN(new_n229_));
  OAI22_X1  g028(.A1(new_n223_), .A2(new_n224_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n220_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n220_), .A2(new_n232_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n207_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n220_), .A2(new_n232_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n205_), .B(new_n206_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(new_n238_), .A3(new_n233_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT76), .ZN(new_n240_));
  AND3_X1   g039(.A1(new_n236_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n240_), .B1(new_n236_), .B2(new_n239_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(G233gat), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT90), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n245_), .A2(G228gat), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(G228gat), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n244_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT87), .B(KEYINPUT88), .ZN(new_n251_));
  OR2_X1    g050(.A1(G155gat), .A2(G162gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G155gat), .A2(G162gat), .ZN(new_n254_));
  XOR2_X1   g053(.A(new_n254_), .B(KEYINPUT1), .Z(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  OR2_X1    g055(.A1(G141gat), .A2(G148gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G141gat), .A2(G148gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n257_), .A2(KEYINPUT3), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT2), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n257_), .A2(KEYINPUT3), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n260_), .A2(new_n262_), .A3(new_n263_), .A4(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n253_), .A2(new_n254_), .A3(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n259_), .A2(new_n266_), .ZN(new_n267_));
  XOR2_X1   g066(.A(KEYINPUT92), .B(KEYINPUT29), .Z(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT91), .ZN(new_n270_));
  INV_X1    g069(.A(G211gat), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n270_), .B1(new_n271_), .B2(G218gat), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n272_), .B1(new_n271_), .B2(G218gat), .ZN(new_n273_));
  XOR2_X1   g072(.A(G197gat), .B(G204gat), .Z(new_n274_));
  OAI21_X1  g073(.A(new_n273_), .B1(new_n274_), .B2(KEYINPUT21), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(KEYINPUT21), .ZN(new_n276_));
  XOR2_X1   g075(.A(new_n275_), .B(new_n276_), .Z(new_n277_));
  AOI21_X1  g076(.A(new_n250_), .B1(new_n269_), .B2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n267_), .A2(KEYINPUT29), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT89), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n277_), .A2(new_n250_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n278_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(G78gat), .B(G106gat), .Z(new_n283_));
  OR2_X1    g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n283_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT94), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT93), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n285_), .A2(new_n288_), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n267_), .A2(KEYINPUT29), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G22gat), .B(G50gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT28), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n290_), .B(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n287_), .B1(new_n289_), .B2(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT93), .B1(new_n282_), .B2(new_n283_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n293_), .ZN(new_n296_));
  NOR3_X1   g095(.A1(new_n295_), .A2(KEYINPUT94), .A3(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n286_), .B1(new_n294_), .B2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n289_), .A2(new_n287_), .A3(new_n293_), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT94), .B1(new_n295_), .B2(new_n296_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n299_), .A2(new_n300_), .A3(new_n285_), .A4(new_n284_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT85), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G183gat), .A2(G190gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT23), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n306_), .B1(G183gat), .B2(G190gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT22), .B(G169gat), .ZN(new_n310_));
  INV_X1    g109(.A(G176gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT81), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n309_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT26), .B(G190gat), .ZN(new_n315_));
  INV_X1    g114(.A(G183gat), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT25), .B1(new_n316_), .B2(KEYINPUT79), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT25), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(G183gat), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n315_), .B(new_n317_), .C1(KEYINPUT79), .C2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT80), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(G169gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n311_), .ZN(new_n324_));
  OR2_X1    g123(.A1(new_n324_), .A2(KEYINPUT24), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n324_), .A2(KEYINPUT24), .A3(new_n308_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n306_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n320_), .A2(new_n321_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n322_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n314_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT30), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT83), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G71gat), .B(G99gat), .ZN(new_n335_));
  INV_X1    g134(.A(G43gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  AND2_X1   g136(.A1(G227gat), .A2(G233gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n334_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT82), .B(G15gat), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n332_), .A2(new_n333_), .A3(new_n339_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  OR2_X1    g143(.A1(new_n332_), .A2(new_n333_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n342_), .B1(new_n341_), .B2(new_n343_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n304_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT86), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT86), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n304_), .B(new_n350_), .C1(new_n346_), .C2(new_n347_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G127gat), .B(G134gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT84), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G113gat), .B(G120gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  XOR2_X1   g154(.A(new_n355_), .B(KEYINPUT31), .Z(new_n356_));
  NAND3_X1  g155(.A1(new_n349_), .A2(new_n351_), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n349_), .A2(new_n351_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n356_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n303_), .A2(new_n357_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n357_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n356_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n302_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n361_), .A2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G1gat), .B(G29gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(G85gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT0), .B(G57gat), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n367_), .B(new_n368_), .Z(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT4), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n267_), .A2(new_n371_), .A3(new_n355_), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n372_), .B(KEYINPUT99), .Z(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G225gat), .A2(G233gat), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n267_), .A2(new_n355_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT98), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  OR2_X1    g178(.A1(new_n267_), .A2(new_n355_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n374_), .B(new_n376_), .C1(new_n371_), .C2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n381_), .A2(new_n376_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n370_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n384_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n382_), .A2(new_n386_), .A3(new_n369_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n331_), .A2(new_n277_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n309_), .A2(new_n312_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n316_), .A2(KEYINPUT25), .ZN(new_n392_));
  AND3_X1   g191(.A1(new_n315_), .A2(new_n319_), .A3(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n391_), .B1(new_n327_), .B2(new_n393_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n390_), .B(KEYINPUT20), .C1(new_n277_), .C2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G226gat), .A2(G233gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT19), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n394_), .A2(new_n277_), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n399_), .B(KEYINPUT20), .C1(new_n277_), .C2(new_n331_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n398_), .B1(new_n397_), .B2(new_n400_), .ZN(new_n401_));
  XOR2_X1   g200(.A(G8gat), .B(G36gat), .Z(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT96), .ZN(new_n403_));
  XOR2_X1   g202(.A(G64gat), .B(G92gat), .Z(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n401_), .A2(new_n407_), .ZN(new_n408_));
  XOR2_X1   g207(.A(new_n408_), .B(KEYINPUT102), .Z(new_n409_));
  AND2_X1   g208(.A1(new_n400_), .A2(new_n397_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n395_), .A2(new_n397_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n407_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n409_), .A2(KEYINPUT27), .A3(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n412_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT97), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(new_n417_), .A3(new_n407_), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT97), .B1(new_n412_), .B2(new_n413_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n414_), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT27), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n389_), .A2(new_n415_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n365_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n381_), .ZN(new_n426_));
  AOI211_X1 g225(.A(new_n376_), .B(new_n373_), .C1(new_n426_), .C2(KEYINPUT4), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT100), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n369_), .B1(new_n426_), .B2(new_n376_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n427_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  OR2_X1    g229(.A1(new_n429_), .A2(new_n428_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n420_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n387_), .B(KEYINPUT33), .ZN(new_n433_));
  AND2_X1   g232(.A1(new_n413_), .A2(KEYINPUT32), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n401_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT101), .ZN(new_n436_));
  OAI22_X1  g235(.A1(new_n435_), .A2(new_n436_), .B1(new_n416_), .B2(new_n434_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n437_), .B1(new_n436_), .B2(new_n435_), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n432_), .A2(new_n433_), .B1(new_n388_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n360_), .A2(new_n357_), .ZN(new_n440_));
  OR3_X1    g239(.A1(new_n439_), .A2(new_n440_), .A3(new_n303_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n243_), .B1(new_n425_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT13), .ZN(new_n443_));
  INV_X1    g242(.A(G230gat), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n444_), .A2(new_n244_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G99gat), .A2(G106gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(KEYINPUT6), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT6), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n448_), .A2(G99gat), .A3(G106gat), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT7), .ZN(new_n451_));
  INV_X1    g250(.A(G99gat), .ZN(new_n452_));
  INV_X1    g251(.A(G106gat), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n451_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n450_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT65), .ZN(new_n458_));
  AND2_X1   g257(.A1(G85gat), .A2(G92gat), .ZN(new_n459_));
  NOR2_X1   g258(.A1(G85gat), .A2(G92gat), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n458_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(G85gat), .ZN(new_n462_));
  INV_X1    g261(.A(G92gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G85gat), .A2(G92gat), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(KEYINPUT65), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n461_), .A2(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT8), .B1(new_n457_), .B2(new_n467_), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n461_), .A2(new_n466_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT8), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n448_), .B1(G99gat), .B2(G106gat), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n446_), .A2(KEYINPUT6), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n455_), .B(new_n454_), .C1(new_n471_), .C2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n469_), .A2(new_n470_), .A3(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n468_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT66), .ZN(new_n476_));
  OR2_X1    g275(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(new_n453_), .A3(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n464_), .A2(KEYINPUT9), .A3(new_n465_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT9), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n459_), .A2(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n483_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT64), .B1(new_n481_), .B2(new_n484_), .ZN(new_n485_));
  AOI22_X1  g284(.A1(new_n447_), .A2(new_n449_), .B1(new_n459_), .B2(new_n482_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT64), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n486_), .A2(new_n487_), .A3(new_n479_), .A4(new_n480_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n485_), .A2(new_n488_), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n475_), .A2(new_n476_), .A3(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n476_), .B1(new_n475_), .B2(new_n489_), .ZN(new_n491_));
  NOR3_X1   g290(.A1(new_n490_), .A2(new_n491_), .A3(new_n231_), .ZN(new_n492_));
  NOR3_X1   g291(.A1(new_n457_), .A2(KEYINPUT8), .A3(new_n467_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n470_), .B1(new_n469_), .B2(new_n473_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n489_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT66), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n475_), .A2(new_n476_), .A3(new_n489_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n232_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n445_), .B1(new_n492_), .B2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G120gat), .B(G148gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT5), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G176gat), .B(G204gat), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n501_), .B(new_n502_), .Z(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT12), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n232_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(new_n495_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n507_), .B1(new_n498_), .B2(KEYINPUT12), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n496_), .A2(new_n497_), .A3(new_n232_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n509_), .B1(new_n444_), .B2(new_n244_), .ZN(new_n510_));
  OAI211_X1 g309(.A(new_n499_), .B(new_n504_), .C1(new_n508_), .C2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT69), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n231_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n514_));
  AOI22_X1  g313(.A1(new_n514_), .A2(new_n505_), .B1(new_n495_), .B2(new_n506_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n492_), .A2(new_n445_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n509_), .ZN(new_n517_));
  AOI22_X1  g316(.A1(new_n515_), .A2(new_n516_), .B1(new_n445_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT68), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n503_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n499_), .B(new_n519_), .C1(new_n508_), .C2(new_n510_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n513_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT70), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n499_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n504_), .B1(new_n525_), .B2(KEYINPUT68), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n526_), .A2(new_n512_), .A3(new_n521_), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n523_), .A2(new_n524_), .A3(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n524_), .B1(new_n523_), .B2(new_n527_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n443_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n526_), .A2(new_n512_), .A3(new_n521_), .ZN(new_n531_));
  AOI22_X1  g330(.A1(new_n526_), .A2(new_n521_), .B1(new_n512_), .B2(new_n511_), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT70), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n523_), .A2(new_n524_), .A3(new_n527_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(KEYINPUT13), .A3(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n530_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n216_), .A2(new_n217_), .ZN(new_n537_));
  XOR2_X1   g336(.A(G29gat), .B(G36gat), .Z(new_n538_));
  XOR2_X1   g337(.A(G43gat), .B(G50gat), .Z(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n537_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT77), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n216_), .A2(new_n217_), .A3(new_n540_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n537_), .A2(KEYINPUT77), .A3(new_n541_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n545_), .A2(G229gat), .A3(G233gat), .A4(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n540_), .B(KEYINPUT15), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(new_n537_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G229gat), .A2(G233gat), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(new_n550_), .A3(new_n544_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n547_), .A2(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(G113gat), .B(G141gat), .Z(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT78), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G169gat), .B(G197gat), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n554_), .B(new_n555_), .Z(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n552_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n547_), .A2(new_n551_), .A3(new_n556_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n536_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n548_), .A2(new_n495_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n563_), .A2(KEYINPUT72), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n496_), .A2(new_n540_), .A3(new_n497_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(KEYINPUT72), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n564_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G232gat), .A2(G233gat), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n568_), .B(KEYINPUT34), .Z(new_n569_));
  XOR2_X1   g368(.A(KEYINPUT71), .B(KEYINPUT35), .Z(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n569_), .B(new_n570_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n565_), .A2(new_n563_), .A3(new_n573_), .ZN(new_n574_));
  AOI22_X1  g373(.A1(new_n567_), .A2(new_n571_), .B1(new_n574_), .B2(KEYINPUT74), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n574_), .A2(KEYINPUT74), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G190gat), .B(G218gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT73), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G134gat), .B(G162gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT36), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n581_), .A2(new_n582_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n577_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n575_), .A2(new_n582_), .A3(new_n581_), .A4(new_n576_), .ZN(new_n586_));
  AND3_X1   g385(.A1(new_n585_), .A2(KEYINPUT37), .A3(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(KEYINPUT37), .B1(new_n585_), .B2(new_n586_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n442_), .A2(new_n562_), .A3(new_n589_), .ZN(new_n590_));
  NOR3_X1   g389(.A1(new_n590_), .A2(G1gat), .A3(new_n389_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(KEYINPUT38), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n585_), .A2(new_n586_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n442_), .A2(new_n562_), .A3(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(G1gat), .B1(new_n594_), .B2(new_n389_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n591_), .A2(KEYINPUT38), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT103), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n591_), .A2(KEYINPUT103), .A3(KEYINPUT38), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n592_), .B(new_n595_), .C1(new_n598_), .C2(new_n599_), .ZN(G1324gat));
  INV_X1    g399(.A(new_n243_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n423_), .B1(new_n361_), .B2(new_n364_), .ZN(new_n602_));
  NOR3_X1   g401(.A1(new_n439_), .A2(new_n440_), .A3(new_n303_), .ZN(new_n603_));
  OAI211_X1 g402(.A(new_n593_), .B(new_n601_), .C1(new_n602_), .C2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n562_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n415_), .A2(new_n422_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n604_), .A2(new_n605_), .A3(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(KEYINPUT39), .B1(new_n608_), .B2(new_n211_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(KEYINPUT104), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n442_), .A2(new_n562_), .A3(new_n593_), .A4(new_n606_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT39), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(new_n612_), .A3(G8gat), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(KEYINPUT105), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT104), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n615_), .B(KEYINPUT39), .C1(new_n608_), .C2(new_n211_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT105), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n611_), .A2(new_n617_), .A3(new_n612_), .A4(G8gat), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n610_), .A2(new_n614_), .A3(new_n616_), .A4(new_n618_), .ZN(new_n619_));
  OR3_X1    g418(.A1(new_n590_), .A2(G8gat), .A3(new_n607_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n619_), .A2(new_n620_), .A3(new_n622_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(G1325gat));
  INV_X1    g425(.A(new_n440_), .ZN(new_n627_));
  OAI21_X1  g426(.A(G15gat), .B1(new_n594_), .B2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT41), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n590_), .A2(G15gat), .A3(new_n627_), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n629_), .A2(new_n630_), .ZN(G1326gat));
  OAI21_X1  g430(.A(G22gat), .B1(new_n594_), .B2(new_n302_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT42), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n302_), .A2(G22gat), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n633_), .B1(new_n590_), .B2(new_n634_), .ZN(G1327gat));
  NOR2_X1   g434(.A1(new_n601_), .A2(new_n593_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n637_), .B1(new_n425_), .B2(new_n441_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(new_n562_), .ZN(new_n639_));
  OR3_X1    g438(.A1(new_n639_), .A2(G29gat), .A3(new_n389_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n589_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n641_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT43), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n601_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  OAI211_X1 g443(.A(KEYINPUT43), .B(new_n641_), .C1(new_n602_), .C2(new_n603_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n644_), .A2(new_n562_), .A3(new_n645_), .ZN(new_n646_));
  XOR2_X1   g445(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n644_), .A2(KEYINPUT44), .A3(new_n645_), .A4(new_n562_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n648_), .A2(new_n388_), .A3(new_n649_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n650_), .A2(KEYINPUT108), .ZN(new_n651_));
  OAI21_X1  g450(.A(G29gat), .B1(new_n650_), .B2(KEYINPUT108), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n640_), .B1(new_n651_), .B2(new_n652_), .ZN(G1328gat));
  NOR2_X1   g452(.A1(new_n607_), .A2(G36gat), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n638_), .A2(new_n562_), .A3(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n655_), .B(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n648_), .A2(new_n606_), .A3(new_n649_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n658_), .B2(G36gat), .ZN(new_n659_));
  XNOR2_X1  g458(.A(KEYINPUT110), .B(KEYINPUT46), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n660_), .ZN(new_n662_));
  AOI211_X1 g461(.A(new_n662_), .B(new_n657_), .C1(new_n658_), .C2(G36gat), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n661_), .A2(new_n663_), .ZN(G1329gat));
  NAND4_X1  g463(.A1(new_n648_), .A2(G43gat), .A3(new_n440_), .A4(new_n649_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n336_), .B1(new_n639_), .B2(new_n627_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g467(.A(new_n639_), .ZN(new_n669_));
  AOI21_X1  g468(.A(G50gat), .B1(new_n669_), .B2(new_n303_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n648_), .A2(new_n649_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n303_), .A2(G50gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n670_), .B1(new_n671_), .B2(new_n672_), .ZN(G1331gat));
  NAND2_X1  g472(.A1(new_n536_), .A2(new_n561_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n604_), .A2(new_n389_), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(G57gat), .ZN(new_n676_));
  INV_X1    g475(.A(new_n674_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n442_), .A2(new_n589_), .A3(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n388_), .A2(new_n676_), .ZN(new_n679_));
  OAI22_X1  g478(.A1(new_n675_), .A2(new_n676_), .B1(new_n678_), .B2(new_n679_), .ZN(G1332gat));
  NAND4_X1  g479(.A1(new_n442_), .A2(new_n593_), .A3(new_n606_), .A4(new_n677_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT48), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n681_), .A2(new_n682_), .A3(G64gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n682_), .B1(new_n681_), .B2(G64gat), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n607_), .A2(G64gat), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n685_), .B(KEYINPUT111), .Z(new_n686_));
  OAI22_X1  g485(.A1(new_n683_), .A2(new_n684_), .B1(new_n678_), .B2(new_n686_), .ZN(G1333gat));
  OR3_X1    g486(.A1(new_n678_), .A2(G71gat), .A3(new_n627_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n442_), .A2(new_n593_), .A3(new_n440_), .A4(new_n677_), .ZN(new_n689_));
  XOR2_X1   g488(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n690_));
  AND3_X1   g489(.A1(new_n689_), .A2(G71gat), .A3(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n689_), .B2(G71gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n688_), .B1(new_n691_), .B2(new_n692_), .ZN(G1334gat));
  OR3_X1    g492(.A1(new_n678_), .A2(G78gat), .A3(new_n302_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n442_), .A2(new_n593_), .A3(new_n303_), .A4(new_n677_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT50), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n695_), .A2(new_n696_), .A3(G78gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n695_), .B2(G78gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n694_), .B1(new_n697_), .B2(new_n698_), .ZN(G1335gat));
  NAND3_X1  g498(.A1(new_n644_), .A2(new_n645_), .A3(new_n677_), .ZN(new_n700_));
  OAI21_X1  g499(.A(G85gat), .B1(new_n700_), .B2(new_n389_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n638_), .A2(new_n677_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n702_), .A2(new_n462_), .A3(new_n388_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(G1336gat));
  INV_X1    g503(.A(KEYINPUT113), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n702_), .A2(new_n606_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n706_), .B2(new_n463_), .ZN(new_n707_));
  AOI211_X1 g506(.A(KEYINPUT113), .B(G92gat), .C1(new_n702_), .C2(new_n606_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n606_), .A2(G92gat), .ZN(new_n709_));
  OAI22_X1  g508(.A1(new_n707_), .A2(new_n708_), .B1(new_n700_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT114), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n710_), .B(new_n711_), .ZN(G1337gat));
  OAI21_X1  g511(.A(G99gat), .B1(new_n700_), .B2(new_n627_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n702_), .A2(new_n477_), .A3(new_n478_), .A4(new_n440_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g515(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT52), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n644_), .A2(new_n303_), .A3(new_n645_), .A4(new_n677_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n719_), .B2(G106gat), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n719_), .A2(new_n718_), .A3(G106gat), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n702_), .A2(new_n453_), .A3(new_n303_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n717_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n722_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n724_), .B(new_n717_), .C1(new_n726_), .C2(new_n720_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n725_), .A2(new_n728_), .ZN(G1339gat));
  NOR2_X1   g528(.A1(new_n243_), .A2(new_n560_), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n530_), .A2(new_n535_), .A3(new_n589_), .A4(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT54), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n731_), .B(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n550_), .B1(new_n218_), .B2(new_n540_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n556_), .B1(new_n735_), .B2(new_n549_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n545_), .A2(new_n546_), .A3(new_n550_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n559_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n560_), .A2(new_n511_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT116), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n560_), .A2(KEYINPUT116), .A3(new_n511_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n515_), .A2(KEYINPUT117), .A3(new_n509_), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n507_), .B(new_n509_), .C1(new_n498_), .C2(KEYINPUT12), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT117), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n747_), .A2(new_n750_), .A3(new_n445_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT55), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n752_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n515_), .A2(new_n516_), .A3(KEYINPUT55), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n751_), .A2(new_n753_), .A3(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT56), .B1(new_n755_), .B2(new_n503_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n755_), .A2(KEYINPUT56), .A3(new_n503_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n746_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  OAI211_X1 g558(.A(KEYINPUT57), .B(new_n593_), .C1(new_n741_), .C2(new_n759_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n739_), .A2(new_n511_), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n755_), .A2(KEYINPUT56), .A3(new_n503_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n761_), .B1(new_n762_), .B2(new_n756_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT58), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  OAI211_X1 g564(.A(KEYINPUT58), .B(new_n761_), .C1(new_n762_), .C2(new_n756_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n765_), .A2(new_n641_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n760_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT57), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n593_), .B1(new_n741_), .B2(new_n759_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n768_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n734_), .B1(new_n771_), .B2(new_n601_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n606_), .A2(new_n389_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n774_), .A2(KEYINPUT59), .A3(new_n364_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n772_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n593_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n739_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n744_), .B(new_n745_), .C1(new_n762_), .C2(new_n756_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n777_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT118), .B1(new_n780_), .B2(KEYINPUT57), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT118), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n770_), .A2(new_n782_), .A3(new_n769_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n781_), .A2(new_n783_), .A3(new_n760_), .A4(new_n767_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n733_), .B1(new_n784_), .B2(new_n243_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n785_), .A2(new_n364_), .A3(new_n774_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT59), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n776_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(G113gat), .B1(new_n788_), .B2(new_n561_), .ZN(new_n789_));
  INV_X1    g588(.A(G113gat), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n786_), .A2(new_n790_), .A3(new_n560_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(G1340gat));
  INV_X1    g591(.A(new_n536_), .ZN(new_n793_));
  OAI21_X1  g592(.A(G120gat), .B1(new_n788_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(G120gat), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n795_), .B1(new_n793_), .B2(KEYINPUT60), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n786_), .B(new_n796_), .C1(KEYINPUT60), .C2(new_n795_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n794_), .A2(new_n797_), .ZN(G1341gat));
  OAI21_X1  g597(.A(G127gat), .B1(new_n788_), .B2(new_n243_), .ZN(new_n799_));
  INV_X1    g598(.A(G127gat), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n786_), .A2(new_n800_), .A3(new_n601_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(G1342gat));
  XNOR2_X1  g601(.A(KEYINPUT119), .B(G134gat), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n788_), .A2(new_n589_), .A3(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(G134gat), .B1(new_n786_), .B2(new_n777_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n804_), .A2(new_n805_), .ZN(G1343gat));
  INV_X1    g605(.A(new_n361_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n782_), .B1(new_n770_), .B2(new_n769_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n808_), .A2(new_n768_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n601_), .B1(new_n809_), .B2(new_n783_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n807_), .B(new_n773_), .C1(new_n810_), .C2(new_n733_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT120), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n784_), .A2(new_n243_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n734_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n815_), .A2(KEYINPUT120), .A3(new_n807_), .A4(new_n773_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n813_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n560_), .ZN(new_n818_));
  XOR2_X1   g617(.A(KEYINPUT121), .B(G141gat), .Z(new_n819_));
  XNOR2_X1  g618(.A(new_n818_), .B(new_n819_), .ZN(G1344gat));
  NAND2_X1  g619(.A1(new_n817_), .A2(new_n536_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g621(.A(KEYINPUT61), .B(G155gat), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT122), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n825_), .B1(new_n817_), .B2(new_n601_), .ZN(new_n826_));
  AOI211_X1 g625(.A(KEYINPUT122), .B(new_n243_), .C1(new_n813_), .C2(new_n816_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n824_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n361_), .B1(new_n814_), .B2(new_n734_), .ZN(new_n829_));
  AOI21_X1  g628(.A(KEYINPUT120), .B1(new_n829_), .B2(new_n773_), .ZN(new_n830_));
  NOR4_X1   g629(.A1(new_n785_), .A2(new_n812_), .A3(new_n361_), .A4(new_n774_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n601_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT122), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n817_), .A2(new_n825_), .A3(new_n601_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(new_n834_), .A3(new_n823_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n828_), .A2(new_n835_), .ZN(G1346gat));
  INV_X1    g635(.A(new_n817_), .ZN(new_n837_));
  OR3_X1    g636(.A1(new_n837_), .A2(G162gat), .A3(new_n593_), .ZN(new_n838_));
  OAI21_X1  g637(.A(G162gat), .B1(new_n837_), .B2(new_n589_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(G1347gat));
  NOR3_X1   g639(.A1(new_n627_), .A2(new_n388_), .A3(new_n607_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(KEYINPUT123), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n842_), .A2(new_n302_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n843_), .A2(new_n772_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n323_), .B1(new_n844_), .B2(new_n560_), .ZN(new_n845_));
  OR2_X1    g644(.A1(new_n845_), .A2(KEYINPUT62), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n844_), .A2(new_n560_), .A3(new_n310_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(KEYINPUT62), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n846_), .A2(new_n847_), .A3(new_n848_), .ZN(G1348gat));
  AOI21_X1  g648(.A(G176gat), .B1(new_n844_), .B2(new_n536_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n815_), .A2(KEYINPUT124), .A3(new_n302_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT124), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n852_), .B1(new_n785_), .B2(new_n303_), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n851_), .A2(new_n842_), .A3(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n793_), .A2(new_n311_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n850_), .B1(new_n854_), .B2(new_n855_), .ZN(G1349gat));
  AOI21_X1  g655(.A(G183gat), .B1(new_n854_), .B2(new_n601_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n243_), .B1(new_n319_), .B2(new_n392_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n857_), .B1(new_n844_), .B2(new_n858_), .ZN(G1350gat));
  INV_X1    g658(.A(new_n844_), .ZN(new_n860_));
  OAI21_X1  g659(.A(G190gat), .B1(new_n860_), .B2(new_n589_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n844_), .A2(new_n777_), .A3(new_n315_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1351gat));
  NOR2_X1   g662(.A1(new_n607_), .A2(new_n388_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n829_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT125), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT125), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n829_), .A2(new_n867_), .A3(new_n864_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n868_), .ZN(new_n869_));
  AND3_X1   g668(.A1(new_n869_), .A2(G197gat), .A3(new_n560_), .ZN(new_n870_));
  AOI21_X1  g669(.A(G197gat), .B1(new_n869_), .B2(new_n560_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1352gat));
  INV_X1    g671(.A(KEYINPUT126), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n793_), .B1(new_n873_), .B2(G204gat), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n875_), .B1(new_n866_), .B2(new_n868_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n873_), .A2(G204gat), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n876_), .B(new_n877_), .ZN(G1353gat));
  AOI21_X1  g677(.A(new_n243_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n880_), .B1(new_n866_), .B2(new_n868_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n881_), .B(new_n882_), .ZN(G1354gat));
  AOI21_X1  g682(.A(G218gat), .B1(new_n869_), .B2(new_n777_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n641_), .A2(G218gat), .ZN(new_n885_));
  XOR2_X1   g684(.A(new_n885_), .B(KEYINPUT127), .Z(new_n886_));
  AOI21_X1  g685(.A(new_n884_), .B1(new_n869_), .B2(new_n886_), .ZN(G1355gat));
endmodule


