//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 1 0 0 0 0 1 1 0 1 0 0 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n821_, new_n822_, new_n823_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n830_, new_n831_, new_n833_, new_n834_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n861_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT18), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G64gat), .B(G92gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  XNOR2_X1  g005(.A(G211gat), .B(G218gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT92), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n208_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G197gat), .B(G204gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT21), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT93), .ZN(new_n214_));
  AND3_X1   g013(.A1(new_n211_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT21), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n212_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n209_), .A2(new_n210_), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(new_n214_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n211_), .A2(new_n213_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n216_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(KEYINPUT23), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n225_), .B1(G183gat), .B2(G190gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227_));
  INV_X1    g026(.A(G176gat), .ZN(new_n228_));
  INV_X1    g027(.A(G169gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT83), .B1(new_n229_), .B2(KEYINPUT22), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT22), .B(G169gat), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n228_), .B(new_n230_), .C1(new_n231_), .C2(KEYINPUT83), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n226_), .A2(new_n227_), .A3(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT26), .B(G190gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT82), .ZN(new_n235_));
  INV_X1    g034(.A(G183gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT25), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT25), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(G183gat), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n234_), .B(new_n237_), .C1(new_n235_), .C2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n229_), .A2(new_n228_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n241_), .A2(KEYINPUT24), .A3(new_n227_), .ZN(new_n242_));
  OR2_X1    g041(.A1(new_n241_), .A2(KEYINPUT24), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n240_), .A2(new_n225_), .A3(new_n242_), .A4(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n233_), .A2(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT20), .B1(new_n223_), .B2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n231_), .A2(new_n228_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n226_), .A2(new_n227_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT98), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT97), .ZN(new_n250_));
  XOR2_X1   g049(.A(KEYINPUT26), .B(G190gat), .Z(new_n251_));
  INV_X1    g050(.A(KEYINPUT95), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n236_), .A2(KEYINPUT25), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n238_), .A2(G183gat), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n252_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n236_), .A2(KEYINPUT25), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n239_), .A2(new_n256_), .A3(KEYINPUT95), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n251_), .B1(new_n255_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n241_), .A2(new_n227_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT96), .B(KEYINPUT24), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n250_), .B1(new_n258_), .B2(new_n261_), .ZN(new_n262_));
  AND3_X1   g061(.A1(new_n239_), .A2(new_n256_), .A3(KEYINPUT95), .ZN(new_n263_));
  AOI21_X1  g062(.A(KEYINPUT95), .B1(new_n239_), .B2(new_n256_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n234_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n261_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(new_n266_), .A3(KEYINPUT97), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n262_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n260_), .A2(new_n229_), .A3(new_n228_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(new_n225_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n249_), .B1(new_n268_), .B2(new_n271_), .ZN(new_n272_));
  AOI211_X1 g071(.A(KEYINPUT98), .B(new_n270_), .C1(new_n262_), .C2(new_n267_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n248_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n246_), .B1(new_n274_), .B2(new_n223_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G226gat), .A2(G233gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT19), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT99), .B1(new_n275_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT99), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n219_), .A2(new_n214_), .B1(new_n211_), .B2(new_n213_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n281_), .A2(new_n215_), .ZN(new_n282_));
  NOR3_X1   g081(.A1(new_n258_), .A2(new_n250_), .A3(new_n261_), .ZN(new_n283_));
  AOI21_X1  g082(.A(KEYINPUT97), .B1(new_n265_), .B2(new_n266_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n271_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT98), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n268_), .A2(new_n249_), .A3(new_n271_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n282_), .B1(new_n288_), .B2(new_n248_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n280_), .B(new_n277_), .C1(new_n289_), .C2(new_n246_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n279_), .A2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n288_), .A2(new_n248_), .A3(new_n282_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n278_), .A2(KEYINPUT20), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n245_), .B1(new_n281_), .B2(new_n215_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT100), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  OAI211_X1 g095(.A(KEYINPUT100), .B(new_n245_), .C1(new_n281_), .C2(new_n215_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n293_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n292_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n206_), .B1(new_n291_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n206_), .ZN(new_n302_));
  AOI211_X1 g101(.A(new_n302_), .B(new_n299_), .C1(new_n279_), .C2(new_n290_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n202_), .B1(new_n301_), .B2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n291_), .A2(new_n206_), .A3(new_n300_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT20), .ZN(new_n306_));
  INV_X1    g105(.A(new_n245_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n306_), .B1(new_n282_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n248_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n309_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n308_), .B1(new_n310_), .B2(new_n282_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n278_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n296_), .A2(new_n297_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n282_), .A2(new_n285_), .A3(new_n248_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n313_), .A2(KEYINPUT20), .A3(new_n277_), .A4(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n312_), .A2(new_n302_), .A3(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n305_), .A2(KEYINPUT27), .A3(new_n316_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n304_), .A2(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(G15gat), .B(G43gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT85), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n245_), .B(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G227gat), .A2(G233gat), .ZN(new_n322_));
  INV_X1    g121(.A(G71gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(G99gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT84), .B(KEYINPUT30), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n321_), .B(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT87), .ZN(new_n329_));
  XOR2_X1   g128(.A(G127gat), .B(G134gat), .Z(new_n330_));
  XOR2_X1   g129(.A(G113gat), .B(G120gat), .Z(new_n331_));
  XOR2_X1   g130(.A(new_n330_), .B(new_n331_), .Z(new_n332_));
  XOR2_X1   g131(.A(new_n332_), .B(KEYINPUT86), .Z(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT31), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n329_), .A2(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n328_), .A2(KEYINPUT87), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n329_), .A2(new_n334_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n335_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(G141gat), .ZN(new_n339_));
  INV_X1    g138(.A(G148gat), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(G141gat), .A2(G148gat), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT88), .ZN(new_n345_));
  INV_X1    g144(.A(G155gat), .ZN(new_n346_));
  INV_X1    g145(.A(G162gat), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n345_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT88), .B1(G155gat), .B2(G162gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G155gat), .A2(G162gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT89), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT89), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n353_), .A2(G155gat), .A3(G162gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n350_), .B1(KEYINPUT1), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT1), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n352_), .A2(new_n354_), .A3(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n344_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT2), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n360_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT3), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n342_), .A2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n361_), .A2(new_n363_), .A3(new_n364_), .A4(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n350_), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n366_), .A2(new_n367_), .A3(new_n355_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n359_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT29), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  OAI211_X1 g170(.A(G228gat), .B(G233gat), .C1(new_n371_), .C2(new_n282_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G228gat), .A2(G233gat), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT90), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n374_), .B1(new_n359_), .B2(new_n368_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n355_), .A2(KEYINPUT1), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n376_), .A2(new_n367_), .A3(new_n358_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(new_n343_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n366_), .A2(new_n367_), .A3(new_n355_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n378_), .A2(KEYINPUT90), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n375_), .A2(new_n380_), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n223_), .B(new_n373_), .C1(new_n381_), .C2(new_n370_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G78gat), .B(G106gat), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n372_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n383_), .B1(new_n372_), .B2(new_n382_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  XOR2_X1   g185(.A(G22gat), .B(G50gat), .Z(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n390_), .B1(new_n381_), .B2(new_n370_), .ZN(new_n391_));
  AOI211_X1 g190(.A(KEYINPUT29), .B(new_n389_), .C1(new_n375_), .C2(new_n380_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n388_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n359_), .A2(new_n374_), .A3(new_n368_), .ZN(new_n394_));
  AOI21_X1  g193(.A(KEYINPUT90), .B1(new_n378_), .B2(new_n379_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n370_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n389_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n381_), .A2(new_n370_), .A3(new_n390_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n397_), .A2(new_n387_), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT94), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n393_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n400_), .B1(new_n393_), .B2(new_n399_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n386_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n393_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n404_), .B1(new_n385_), .B2(new_n384_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT4), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n375_), .A2(new_n407_), .A3(new_n380_), .A4(new_n332_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G225gat), .A2(G233gat), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n375_), .A2(new_n332_), .A3(new_n380_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n332_), .ZN(new_n413_));
  AOI21_X1  g212(.A(KEYINPUT101), .B1(new_n369_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n375_), .A2(KEYINPUT101), .A3(new_n380_), .A4(new_n332_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n411_), .B1(new_n417_), .B2(KEYINPUT4), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  XOR2_X1   g218(.A(G1gat), .B(G29gat), .Z(new_n420_));
  XNOR2_X1  g219(.A(G57gat), .B(G85gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT102), .B(KEYINPUT0), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n417_), .A2(new_n409_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n419_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n426_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n424_), .B1(new_n428_), .B2(new_n418_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n338_), .A2(new_n406_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n318_), .A2(new_n431_), .ZN(new_n432_));
  XOR2_X1   g231(.A(new_n432_), .B(KEYINPUT107), .Z(new_n433_));
  INV_X1    g232(.A(KEYINPUT105), .ZN(new_n434_));
  NOR3_X1   g233(.A1(new_n275_), .A2(KEYINPUT99), .A3(new_n278_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n280_), .B1(new_n311_), .B2(new_n277_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n300_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(new_n302_), .ZN(new_n438_));
  AOI21_X1  g237(.A(KEYINPUT27), .B1(new_n438_), .B2(new_n305_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n427_), .A2(new_n429_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n316_), .A2(KEYINPUT27), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n440_), .B(new_n406_), .C1(new_n303_), .C2(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n434_), .B1(new_n439_), .B2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n430_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n304_), .A2(KEYINPUT105), .A3(new_n317_), .A4(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n426_), .A2(new_n425_), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT33), .B1(new_n446_), .B2(new_n418_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT33), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n419_), .A2(new_n448_), .A3(new_n425_), .A4(new_n426_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n417_), .A2(new_n410_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n424_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT103), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n417_), .A2(KEYINPUT4), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n408_), .A2(new_n409_), .ZN(new_n454_));
  AOI22_X1  g253(.A1(new_n451_), .A2(new_n452_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n450_), .A2(KEYINPUT103), .A3(new_n424_), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n447_), .A2(new_n449_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n457_), .A2(new_n305_), .A3(new_n438_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n206_), .A2(KEYINPUT32), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n312_), .A2(new_n315_), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n460_), .A2(new_n461_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n291_), .A2(new_n300_), .A3(new_n459_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n406_), .B1(new_n458_), .B2(new_n464_), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n443_), .B(new_n445_), .C1(new_n465_), .C2(KEYINPUT104), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n301_), .A2(new_n303_), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n467_), .A2(new_n457_), .B1(new_n463_), .B2(new_n462_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT104), .ZN(new_n469_));
  NOR3_X1   g268(.A1(new_n468_), .A2(new_n469_), .A3(new_n406_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n338_), .B1(new_n466_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT106), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  OAI211_X1 g272(.A(KEYINPUT106), .B(new_n338_), .C1(new_n466_), .C2(new_n470_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n433_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G85gat), .B(G92gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT69), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G99gat), .A2(G106gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT6), .ZN(new_n479_));
  OR3_X1    g278(.A1(KEYINPUT67), .A2(G99gat), .A3(G106gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(KEYINPUT7), .ZN(new_n481_));
  OR4_X1    g280(.A1(KEYINPUT67), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n479_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n477_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT68), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT70), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT8), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT10), .B(G99gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT66), .ZN(new_n490_));
  INV_X1    g289(.A(G106gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT9), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n476_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(G85gat), .A3(G92gat), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n492_), .A2(new_n479_), .A3(new_n494_), .A4(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n484_), .A2(KEYINPUT70), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT8), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n488_), .B(new_n496_), .C1(new_n486_), .C2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G57gat), .B(G64gat), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n500_), .A2(KEYINPUT11), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(KEYINPUT11), .ZN(new_n502_));
  XOR2_X1   g301(.A(G71gat), .B(G78gat), .Z(new_n503_));
  NAND3_X1  g302(.A1(new_n501_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n502_), .A2(new_n503_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n499_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT71), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n509_), .A2(KEYINPUT12), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G230gat), .A2(G233gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n499_), .A2(new_n507_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n514_), .B1(new_n509_), .B2(KEYINPUT12), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n510_), .A2(new_n513_), .A3(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n513_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n508_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n517_), .B1(new_n518_), .B2(new_n514_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n516_), .A2(new_n519_), .ZN(new_n520_));
  XOR2_X1   g319(.A(G120gat), .B(G148gat), .Z(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G176gat), .B(G204gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n525_), .B(KEYINPUT73), .Z(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n520_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT74), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n516_), .A2(new_n519_), .A3(new_n525_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n529_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n534_), .A2(KEYINPUT13), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(KEYINPUT13), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G1gat), .B(G8gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT80), .ZN(new_n540_));
  OR2_X1    g339(.A1(G15gat), .A2(G22gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G15gat), .A2(G22gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G1gat), .A2(G8gat), .ZN(new_n543_));
  AOI22_X1  g342(.A1(new_n541_), .A2(new_n542_), .B1(KEYINPUT14), .B2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n540_), .B(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G29gat), .B(G36gat), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(G43gat), .B(G50gat), .Z(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n545_), .B(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n551_), .A2(G229gat), .A3(G233gat), .ZN(new_n552_));
  XOR2_X1   g351(.A(KEYINPUT75), .B(KEYINPUT15), .Z(new_n553_));
  XNOR2_X1  g352(.A(new_n549_), .B(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(new_n545_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G229gat), .A2(G233gat), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n555_), .B(new_n556_), .C1(new_n545_), .C2(new_n550_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n552_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G113gat), .B(G141gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G169gat), .B(G197gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n559_), .B(new_n560_), .Z(new_n561_));
  XNOR2_X1  g360(.A(new_n558_), .B(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT81), .Z(new_n563_));
  NOR3_X1   g362(.A1(new_n475_), .A2(new_n538_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT37), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n499_), .A2(new_n550_), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n566_), .B(KEYINPUT76), .Z(new_n567_));
  INV_X1    g366(.A(KEYINPUT35), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G232gat), .A2(G233gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT34), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  AOI22_X1  g370(.A1(new_n499_), .A2(new_n554_), .B1(new_n568_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n567_), .A2(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n571_), .A2(new_n568_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n567_), .B(new_n572_), .C1(new_n568_), .C2(new_n571_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(G190gat), .B(G218gat), .Z(new_n578_));
  XNOR2_X1  g377(.A(G134gat), .B(G162gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT36), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT79), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n577_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT78), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n565_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n580_), .A2(new_n581_), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n587_), .B(KEYINPUT77), .Z(new_n588_));
  NAND3_X1  g387(.A1(new_n575_), .A2(new_n576_), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n584_), .A2(new_n589_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n586_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n586_), .A2(new_n590_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G231gat), .A2(G233gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n506_), .B(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(new_n545_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT17), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G127gat), .B(G155gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT16), .ZN(new_n600_));
  XOR2_X1   g399(.A(G183gat), .B(G211gat), .Z(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  NOR3_X1   g401(.A1(new_n597_), .A2(new_n598_), .A3(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(KEYINPUT17), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n603_), .B1(new_n597_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n594_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n564_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT108), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n564_), .A2(KEYINPUT108), .A3(new_n607_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n440_), .A2(G1gat), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n612_), .A2(KEYINPUT38), .A3(new_n613_), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n614_), .A2(KEYINPUT109), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(KEYINPUT109), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n612_), .A2(new_n613_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n590_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n475_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n562_), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n538_), .A2(new_n606_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(G1gat), .B1(new_n622_), .B2(new_n440_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n623_), .A2(KEYINPUT38), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n615_), .B(new_n616_), .C1(new_n617_), .C2(new_n624_), .ZN(G1324gat));
  INV_X1    g424(.A(G8gat), .ZN(new_n626_));
  INV_X1    g425(.A(new_n318_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n612_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n619_), .A2(new_n621_), .A3(new_n627_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(G8gat), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT110), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT110), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n629_), .A2(new_n633_), .A3(G8gat), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n631_), .A2(new_n632_), .A3(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n632_), .B1(new_n631_), .B2(new_n634_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n628_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT40), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n628_), .B(KEYINPUT40), .C1(new_n635_), .C2(new_n636_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1325gat));
  OAI21_X1  g440(.A(G15gat), .B1(new_n622_), .B2(new_n338_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT41), .Z(new_n643_));
  INV_X1    g442(.A(new_n612_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n338_), .A2(G15gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n643_), .B1(new_n644_), .B2(new_n645_), .ZN(G1326gat));
  INV_X1    g445(.A(new_n406_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G22gat), .B1(new_n622_), .B2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT42), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n647_), .A2(G22gat), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n649_), .B1(new_n644_), .B2(new_n650_), .ZN(G1327gat));
  NOR2_X1   g450(.A1(new_n590_), .A2(new_n605_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n564_), .A2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(G29gat), .B1(new_n653_), .B2(new_n430_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n538_), .A2(new_n605_), .A3(new_n620_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n475_), .A2(KEYINPUT43), .A3(new_n593_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT43), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n432_), .B(KEYINPUT107), .ZN(new_n658_));
  INV_X1    g457(.A(new_n474_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n469_), .B1(new_n468_), .B2(new_n406_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n458_), .A2(new_n464_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n661_), .A2(KEYINPUT104), .A3(new_n647_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n660_), .A2(new_n662_), .A3(new_n443_), .A4(new_n445_), .ZN(new_n663_));
  AOI21_X1  g462(.A(KEYINPUT106), .B1(new_n663_), .B2(new_n338_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n658_), .B1(new_n659_), .B2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n657_), .B1(new_n665_), .B2(new_n594_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n655_), .B1(new_n656_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(KEYINPUT43), .B1(new_n475_), .B2(new_n593_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n665_), .A2(new_n657_), .A3(new_n594_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n672_), .A2(KEYINPUT44), .A3(new_n655_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n669_), .A2(new_n673_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n430_), .A2(G29gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n654_), .B1(new_n674_), .B2(new_n675_), .ZN(G1328gat));
  INV_X1    g475(.A(KEYINPUT46), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n669_), .A2(new_n627_), .A3(new_n673_), .ZN(new_n678_));
  INV_X1    g477(.A(G36gat), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n318_), .B(KEYINPUT111), .Z(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n653_), .A2(new_n679_), .A3(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT45), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n683_), .B(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n677_), .B1(new_n680_), .B2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n683_), .B(KEYINPUT45), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n687_), .B(KEYINPUT46), .C1(new_n679_), .C2(new_n678_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(G1329gat));
  INV_X1    g488(.A(new_n338_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(G43gat), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n669_), .A2(new_n673_), .A3(KEYINPUT112), .A4(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n669_), .A2(new_n673_), .A3(new_n692_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT112), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(G43gat), .B1(new_n653_), .B2(new_n690_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n699_));
  AND4_X1   g498(.A1(new_n693_), .A2(new_n696_), .A3(new_n698_), .A4(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n697_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n699_), .B1(new_n701_), .B2(new_n693_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n700_), .A2(new_n702_), .ZN(G1330gat));
  INV_X1    g502(.A(G50gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n653_), .A2(new_n704_), .A3(new_n406_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n669_), .A2(new_n406_), .A3(new_n673_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT114), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n706_), .A2(new_n707_), .A3(G50gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n706_), .B2(G50gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n705_), .B1(new_n708_), .B2(new_n709_), .ZN(G1331gat));
  NOR3_X1   g509(.A1(new_n475_), .A2(new_n537_), .A3(new_n562_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n607_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT115), .Z(new_n713_));
  AOI21_X1  g512(.A(G57gat), .B1(new_n713_), .B2(new_n430_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n563_), .A2(new_n605_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n537_), .A2(new_n715_), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n619_), .A2(G57gat), .A3(new_n430_), .A4(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT116), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n714_), .A2(new_n718_), .ZN(G1332gat));
  INV_X1    g518(.A(G64gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n713_), .A2(new_n720_), .A3(new_n682_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n619_), .A2(new_n716_), .ZN(new_n722_));
  OAI21_X1  g521(.A(G64gat), .B1(new_n722_), .B2(new_n681_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT48), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n721_), .A2(new_n724_), .ZN(G1333gat));
  NAND3_X1  g524(.A1(new_n713_), .A2(new_n323_), .A3(new_n690_), .ZN(new_n726_));
  OAI21_X1  g525(.A(G71gat), .B1(new_n722_), .B2(new_n338_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT49), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1334gat));
  INV_X1    g528(.A(G78gat), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n713_), .A2(new_n730_), .A3(new_n406_), .ZN(new_n731_));
  OAI21_X1  g530(.A(G78gat), .B1(new_n722_), .B2(new_n647_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT50), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1335gat));
  NOR2_X1   g533(.A1(new_n562_), .A2(new_n605_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n538_), .A2(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n736_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(G85gat), .B1(new_n738_), .B2(new_n440_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n711_), .A2(new_n652_), .ZN(new_n740_));
  INV_X1    g539(.A(G85gat), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n740_), .A2(new_n741_), .A3(new_n430_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(new_n742_), .ZN(G1336gat));
  OAI21_X1  g542(.A(G92gat), .B1(new_n738_), .B2(new_n681_), .ZN(new_n744_));
  INV_X1    g543(.A(G92gat), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n740_), .A2(new_n745_), .A3(new_n627_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(G1337gat));
  NAND3_X1  g546(.A1(new_n740_), .A2(new_n490_), .A3(new_n690_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n738_), .A2(new_n338_), .ZN(new_n749_));
  INV_X1    g548(.A(G99gat), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n748_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g551(.A1(new_n740_), .A2(new_n491_), .A3(new_n406_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n737_), .A2(new_n406_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n755_), .B2(G106gat), .ZN(new_n756_));
  AOI211_X1 g555(.A(KEYINPUT52), .B(new_n491_), .C1(new_n737_), .C2(new_n406_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n753_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT53), .ZN(G1339gat));
  XNOR2_X1  g558(.A(new_n715_), .B(KEYINPUT117), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n760_), .B1(new_n592_), .B2(new_n591_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT54), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n761_), .A2(new_n762_), .A3(new_n537_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n761_), .B2(new_n537_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n516_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n516_), .A2(new_n766_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n510_), .A2(new_n515_), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n767_), .B(new_n768_), .C1(new_n513_), .C2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n527_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT56), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n771_), .A2(new_n772_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n558_), .A2(new_n561_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n545_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n556_), .B1(new_n778_), .B2(new_n549_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n561_), .B1(new_n779_), .B2(new_n555_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n551_), .A2(new_n556_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n777_), .B1(KEYINPUT119), .B2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(KEYINPUT119), .B2(new_n782_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n530_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n776_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT58), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n776_), .A2(KEYINPUT58), .A3(new_n786_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n594_), .A3(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n530_), .A2(new_n562_), .ZN(new_n793_));
  XOR2_X1   g592(.A(new_n793_), .B(KEYINPUT118), .Z(new_n794_));
  AOI21_X1  g593(.A(new_n794_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n534_), .A2(new_n784_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n792_), .B1(new_n797_), .B2(new_n618_), .ZN(new_n798_));
  OAI211_X1 g597(.A(KEYINPUT57), .B(new_n590_), .C1(new_n795_), .C2(new_n796_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n791_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n765_), .B1(new_n800_), .B2(new_n606_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n318_), .A2(new_n690_), .A3(new_n430_), .A4(new_n647_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(G113gat), .B1(new_n803_), .B2(new_n562_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(KEYINPUT59), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT59), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n806_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n807_), .ZN(new_n808_));
  XOR2_X1   g607(.A(KEYINPUT120), .B(G113gat), .Z(new_n809_));
  NOR2_X1   g608(.A1(new_n563_), .A2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n804_), .B1(new_n808_), .B2(new_n810_), .ZN(G1340gat));
  INV_X1    g610(.A(G120gat), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n812_), .B1(new_n537_), .B2(KEYINPUT60), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n803_), .B(new_n813_), .C1(KEYINPUT60), .C2(new_n812_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n537_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n814_), .B1(new_n815_), .B2(new_n812_), .ZN(G1341gat));
  INV_X1    g615(.A(G127gat), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n803_), .A2(new_n817_), .A3(new_n605_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n606_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n818_), .B1(new_n819_), .B2(new_n817_), .ZN(G1342gat));
  INV_X1    g619(.A(G134gat), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n803_), .A2(new_n821_), .A3(new_n618_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n593_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n823_), .B2(new_n821_), .ZN(G1343gat));
  NOR4_X1   g623(.A1(new_n682_), .A2(new_n690_), .A3(new_n440_), .A4(new_n647_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n801_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n562_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n538_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(KEYINPUT121), .B(G148gat), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n830_), .B(new_n831_), .ZN(G1345gat));
  NAND2_X1  g631(.A1(new_n827_), .A2(new_n605_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(KEYINPUT61), .B(G155gat), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n833_), .B(new_n834_), .ZN(G1346gat));
  INV_X1    g634(.A(new_n801_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n836_), .A2(new_n347_), .A3(new_n618_), .A4(new_n825_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n801_), .A2(new_n593_), .A3(new_n826_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(new_n347_), .B2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT122), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT122), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n837_), .B(new_n841_), .C1(new_n347_), .C2(new_n838_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(G1347gat));
  NOR2_X1   g642(.A1(new_n801_), .A2(new_n681_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n431_), .ZN(new_n845_));
  OAI211_X1 g644(.A(KEYINPUT62), .B(G169gat), .C1(new_n845_), .C2(new_n620_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT62), .ZN(new_n847_));
  INV_X1    g646(.A(new_n431_), .ZN(new_n848_));
  NOR4_X1   g647(.A1(new_n801_), .A2(new_n848_), .A3(new_n620_), .A4(new_n681_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n847_), .B1(new_n849_), .B2(new_n229_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n231_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n846_), .A2(new_n850_), .A3(new_n851_), .ZN(G1348gat));
  NAND3_X1  g651(.A1(new_n844_), .A2(new_n431_), .A3(new_n538_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(G176gat), .ZN(G1349gat));
  NAND4_X1  g653(.A1(new_n765_), .A2(new_n605_), .A3(new_n431_), .A4(new_n682_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(G183gat), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n263_), .A2(new_n264_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(new_n855_), .ZN(new_n858_));
  XOR2_X1   g657(.A(new_n858_), .B(KEYINPUT123), .Z(G1350gat));
  OAI21_X1  g658(.A(G190gat), .B1(new_n845_), .B2(new_n593_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n618_), .A2(new_n234_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n845_), .B2(new_n861_), .ZN(G1351gat));
  NAND2_X1  g661(.A1(new_n444_), .A2(new_n338_), .ZN(new_n863_));
  XOR2_X1   g662(.A(new_n863_), .B(KEYINPUT124), .Z(new_n864_));
  NAND3_X1  g663(.A1(new_n844_), .A2(new_n562_), .A3(new_n864_), .ZN(new_n865_));
  XOR2_X1   g664(.A(KEYINPUT125), .B(G197gat), .Z(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1352gat));
  NAND3_X1  g666(.A1(new_n844_), .A2(new_n538_), .A3(new_n864_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT126), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(G204gat), .ZN(new_n870_));
  XOR2_X1   g669(.A(new_n868_), .B(new_n870_), .Z(G1353gat));
  NAND3_X1  g670(.A1(new_n844_), .A2(new_n605_), .A3(new_n864_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT63), .B(G211gat), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n872_), .B2(new_n875_), .ZN(G1354gat));
  NOR2_X1   g675(.A1(new_n590_), .A2(G218gat), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n836_), .A2(new_n682_), .A3(new_n864_), .A4(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n864_), .ZN(new_n879_));
  NOR4_X1   g678(.A1(new_n801_), .A2(new_n593_), .A3(new_n681_), .A4(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(G218gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n878_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT127), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n878_), .B(KEYINPUT127), .C1(new_n880_), .C2(new_n881_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1355gat));
endmodule


