//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 1 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n623_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n866_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  INV_X1    g001(.A(G197gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(G204gat), .ZN(new_n204_));
  INV_X1    g003(.A(G204gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n205_), .A2(G197gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT21), .B1(new_n204_), .B2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT87), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n206_), .B1(new_n209_), .B2(new_n204_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n210_), .B1(new_n209_), .B2(new_n204_), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n207_), .B(new_n208_), .C1(new_n211_), .C2(KEYINPUT21), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT21), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT88), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n213_), .B1(new_n208_), .B2(new_n214_), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n211_), .B(new_n215_), .C1(new_n214_), .C2(new_n208_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n212_), .A2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT26), .B(G190gat), .ZN(new_n218_));
  INV_X1    g017(.A(G183gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT79), .B1(new_n219_), .B2(KEYINPUT25), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT25), .B(G183gat), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n218_), .B(new_n220_), .C1(new_n221_), .C2(KEYINPUT79), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(KEYINPUT80), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT23), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(KEYINPUT81), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n225_), .B1(new_n226_), .B2(KEYINPUT23), .ZN(new_n227_));
  NOR2_X1   g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT24), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT24), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n230_), .B1(new_n232_), .B2(new_n228_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n227_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n223_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT22), .B(G169gat), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n231_), .B1(new_n239_), .B2(G176gat), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n226_), .A2(KEYINPUT23), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n224_), .A2(KEYINPUT23), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT82), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(G183gat), .A2(G190gat), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n240_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n217_), .B1(new_n237_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n217_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n227_), .A2(new_n246_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n238_), .B(KEYINPUT92), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n250_), .B(new_n231_), .C1(G176gat), .C2(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n233_), .B1(new_n221_), .B2(new_n218_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n244_), .A2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n249_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n248_), .A2(KEYINPUT20), .A3(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G226gat), .A2(G233gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT19), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(KEYINPUT91), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n241_), .A2(new_n243_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n261_), .A2(new_n245_), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n249_), .B(new_n236_), .C1(new_n262_), .C2(new_n240_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n254_), .A2(new_n252_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(new_n217_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n263_), .A2(KEYINPUT20), .A3(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n259_), .B1(new_n260_), .B2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G8gat), .B(G36gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT18), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G64gat), .B(G92gat), .ZN(new_n270_));
  XOR2_X1   g069(.A(new_n269_), .B(new_n270_), .Z(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n267_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT97), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n266_), .A2(new_n260_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n258_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n248_), .A2(KEYINPUT20), .A3(new_n276_), .A4(new_n255_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(new_n271_), .A3(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n273_), .A2(new_n274_), .A3(new_n278_), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n278_), .A2(new_n274_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n202_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT93), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n278_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n278_), .A2(new_n282_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n275_), .A2(new_n277_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(new_n272_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n283_), .A2(new_n284_), .A3(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n281_), .B1(new_n202_), .B2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G127gat), .B(G134gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G113gat), .B(G120gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT84), .ZN(new_n292_));
  AND2_X1   g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293_));
  NOR2_X1   g092(.A1(G155gat), .A2(G162gat), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(G141gat), .A2(G148gat), .ZN(new_n296_));
  XOR2_X1   g095(.A(new_n296_), .B(KEYINPUT3), .Z(new_n297_));
  NAND2_X1  g096(.A1(G141gat), .A2(G148gat), .ZN(new_n298_));
  XOR2_X1   g097(.A(new_n298_), .B(KEYINPUT2), .Z(new_n299_));
  OAI21_X1  g098(.A(new_n295_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT1), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n294_), .B1(new_n293_), .B2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n302_), .B1(new_n301_), .B2(new_n293_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n296_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n303_), .A2(new_n298_), .A3(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n300_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(KEYINPUT94), .B(KEYINPUT4), .Z(new_n308_));
  OR3_X1    g107(.A1(new_n292_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n291_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n310_), .B1(new_n292_), .B2(new_n307_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT4), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n309_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G225gat), .A2(G233gat), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n311_), .A2(new_n314_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G1gat), .B(G29gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(G85gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT0), .B(G57gat), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n320_), .B(new_n321_), .Z(new_n322_));
  NAND2_X1  g121(.A1(new_n318_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n322_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n316_), .A2(new_n324_), .A3(new_n317_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(KEYINPUT89), .B(KEYINPUT29), .Z(new_n327_));
  OAI21_X1  g126(.A(new_n217_), .B1(new_n307_), .B2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n328_), .A2(G228gat), .A3(G233gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G228gat), .A2(G233gat), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT29), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n217_), .B(new_n330_), .C1(new_n307_), .C2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n329_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G78gat), .B(G106gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n334_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n329_), .A2(new_n336_), .A3(new_n332_), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n335_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(G50gat), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n307_), .A2(KEYINPUT28), .A3(new_n331_), .ZN(new_n340_));
  INV_X1    g139(.A(G22gat), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT28), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n342_), .B1(new_n306_), .B2(KEYINPUT29), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n340_), .A2(new_n341_), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n341_), .B1(new_n340_), .B2(new_n343_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n339_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT90), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n337_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n346_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n350_), .A2(G50gat), .A3(new_n344_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n338_), .A2(new_n347_), .A3(new_n349_), .A4(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n349_), .A2(new_n347_), .A3(new_n351_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n335_), .A2(new_n337_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n352_), .A2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G71gat), .B(G99gat), .ZN(new_n357_));
  INV_X1    g156(.A(G43gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT30), .ZN(new_n360_));
  XOR2_X1   g159(.A(KEYINPUT83), .B(G15gat), .Z(new_n361_));
  NAND2_X1  g160(.A1(G227gat), .A2(G233gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n360_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n360_), .A2(new_n363_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n237_), .A2(new_n247_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n364_), .B(new_n365_), .C1(new_n237_), .C2(new_n247_), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n292_), .B(KEYINPUT31), .Z(new_n370_));
  NAND4_X1  g169(.A1(new_n368_), .A2(KEYINPUT85), .A3(new_n369_), .A4(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n368_), .A2(new_n369_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n292_), .B(KEYINPUT31), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT85), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n371_), .B1(new_n373_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n356_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(KEYINPUT86), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT86), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n371_), .B(new_n381_), .C1(new_n373_), .C2(new_n376_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n380_), .A2(new_n382_), .A3(new_n352_), .A4(new_n355_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n326_), .B1(new_n379_), .B2(new_n383_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n271_), .A2(KEYINPUT32), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n267_), .A2(new_n385_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n326_), .B(new_n386_), .C1(new_n285_), .C2(new_n385_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT33), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n323_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n318_), .A2(KEYINPUT33), .A3(new_n322_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT96), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n324_), .B1(new_n311_), .B2(new_n314_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT95), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n309_), .B(new_n314_), .C1(new_n311_), .C2(new_n312_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT95), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n396_), .B(new_n324_), .C1(new_n311_), .C2(new_n314_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n391_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  AND4_X1   g197(.A1(new_n391_), .A2(new_n393_), .A3(new_n397_), .A4(new_n394_), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n389_), .B(new_n390_), .C1(new_n398_), .C2(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n387_), .B1(new_n400_), .B2(new_n287_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n356_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n380_), .A2(new_n382_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  AOI22_X1  g203(.A1(new_n288_), .A2(new_n384_), .B1(new_n401_), .B2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G113gat), .B(G141gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G169gat), .B(G197gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  XOR2_X1   g209(.A(new_n410_), .B(KEYINPUT78), .Z(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G43gat), .B(G50gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(G36gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(G29gat), .ZN(new_n416_));
  INV_X1    g215(.A(G29gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(G36gat), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n416_), .A2(new_n418_), .A3(KEYINPUT67), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT67), .B1(new_n416_), .B2(new_n418_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n414_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT67), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n417_), .A2(G36gat), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n415_), .A2(G29gat), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n422_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n416_), .A2(new_n418_), .A3(KEYINPUT67), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n426_), .A3(new_n413_), .ZN(new_n427_));
  AOI21_X1  g226(.A(KEYINPUT15), .B1(new_n421_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G15gat), .B(G22gat), .ZN(new_n430_));
  INV_X1    g229(.A(G1gat), .ZN(new_n431_));
  INV_X1    g230(.A(G8gat), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT14), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n430_), .A2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G1gat), .B(G8gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n421_), .A2(new_n427_), .A3(KEYINPUT15), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n429_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G229gat), .A2(G233gat), .ZN(new_n439_));
  XOR2_X1   g238(.A(new_n434_), .B(new_n435_), .Z(new_n440_));
  NAND2_X1  g239(.A1(new_n421_), .A2(new_n427_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n438_), .A2(new_n439_), .A3(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n436_), .A2(new_n427_), .A3(new_n421_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n439_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n443_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT77), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n412_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n411_), .A2(KEYINPUT77), .A3(new_n448_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n405_), .A2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G57gat), .B(G64gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G71gat), .B(G78gat), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n454_), .A2(new_n455_), .A3(KEYINPUT11), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(KEYINPUT11), .ZN(new_n457_));
  INV_X1    g256(.A(new_n455_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n454_), .A2(KEYINPUT11), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n456_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G231gat), .A2(G233gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT72), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(new_n436_), .ZN(new_n465_));
  XOR2_X1   g264(.A(G127gat), .B(G155gat), .Z(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G183gat), .B(G211gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(new_n470_), .B(KEYINPUT17), .Z(new_n471_));
  NAND2_X1  g270(.A1(new_n465_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT74), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n465_), .A2(KEYINPUT74), .A3(new_n471_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n470_), .A2(KEYINPUT17), .ZN(new_n476_));
  OR2_X1    g275(.A1(new_n465_), .A2(new_n476_), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n474_), .A2(new_n475_), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  OR2_X1    g282(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n484_));
  INV_X1    g283(.A(G106gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n484_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(G85gat), .ZN(new_n488_));
  INV_X1    g287(.A(G92gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(G85gat), .A2(G92gat), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(KEYINPUT9), .A3(new_n491_), .ZN(new_n492_));
  OR2_X1    g291(.A1(new_n491_), .A2(KEYINPUT9), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n483_), .A2(new_n487_), .A3(new_n492_), .A4(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT7), .ZN(new_n495_));
  INV_X1    g294(.A(G99gat), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n495_), .A2(new_n496_), .A3(new_n485_), .A4(KEYINPUT65), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT65), .ZN(new_n498_));
  OAI22_X1  g297(.A1(new_n498_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G99gat), .A2(G106gat), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT6), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n497_), .A2(new_n499_), .A3(new_n502_), .A4(new_n480_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT8), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n490_), .A2(new_n491_), .ZN(new_n505_));
  AND3_X1   g304(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n504_), .B1(new_n503_), .B2(new_n505_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n494_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT66), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  OAI211_X1 g309(.A(KEYINPUT66), .B(new_n494_), .C1(new_n506_), .C2(new_n507_), .ZN(new_n511_));
  OAI211_X1 g310(.A(KEYINPUT12), .B(new_n456_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n510_), .A2(new_n511_), .A3(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G230gat), .A2(G233gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT64), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n461_), .B(new_n494_), .C1(new_n507_), .C2(new_n506_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT12), .ZN(new_n519_));
  INV_X1    g318(.A(new_n494_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n503_), .A2(new_n505_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT8), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n520_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n519_), .B1(new_n524_), .B2(new_n461_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n514_), .A2(new_n517_), .A3(new_n518_), .A4(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n524_), .A2(new_n461_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n518_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n516_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G120gat), .B(G148gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT5), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G176gat), .B(G204gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n526_), .A2(new_n529_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n533_), .B1(new_n526_), .B2(new_n529_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n537_), .A2(KEYINPUT13), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(KEYINPUT13), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n421_), .A2(KEYINPUT15), .A3(new_n427_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n542_), .A2(new_n428_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n510_), .A2(new_n543_), .A3(new_n511_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G232gat), .A2(G233gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT34), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n546_), .A2(KEYINPUT35), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n547_), .B1(new_n524_), .B2(new_n441_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n544_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n546_), .A2(KEYINPUT35), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n550_), .A2(KEYINPUT68), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n550_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT68), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n549_), .A2(new_n552_), .A3(new_n556_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n544_), .A2(new_n554_), .A3(new_n553_), .A4(new_n548_), .ZN(new_n558_));
  XOR2_X1   g357(.A(G190gat), .B(G218gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT69), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G134gat), .B(G162gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT36), .Z(new_n563_));
  AND3_X1   g362(.A1(new_n557_), .A2(new_n558_), .A3(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n562_), .A2(KEYINPUT36), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n566_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT37), .B1(new_n564_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT70), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT37), .ZN(new_n571_));
  AOI211_X1 g370(.A(new_n551_), .B(new_n555_), .C1(new_n544_), .C2(new_n548_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n558_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n565_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n557_), .A2(new_n563_), .A3(new_n558_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n571_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT70), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT71), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n557_), .A2(new_n563_), .A3(KEYINPUT71), .A4(new_n558_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n567_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  AOI22_X1  g380(.A1(new_n570_), .A2(new_n577_), .B1(new_n571_), .B2(new_n581_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n479_), .A2(new_n541_), .A3(new_n582_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n453_), .A2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n326_), .B(KEYINPUT98), .ZN(new_n585_));
  AND3_X1   g384(.A1(new_n584_), .A2(new_n431_), .A3(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n586_), .A2(KEYINPUT38), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT100), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT99), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n589_), .B1(new_n541_), .B2(new_n452_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n452_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n540_), .A2(KEYINPUT99), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  NOR4_X1   g392(.A1(new_n405_), .A2(new_n593_), .A3(new_n581_), .A4(new_n479_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n431_), .B1(new_n594_), .B2(new_n326_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n595_), .B1(new_n586_), .B2(KEYINPUT38), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n588_), .A2(new_n596_), .ZN(G1324gat));
  INV_X1    g396(.A(new_n281_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n287_), .A2(new_n202_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n584_), .A2(new_n432_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT39), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n594_), .A2(new_n600_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n602_), .B1(new_n603_), .B2(G8gat), .ZN(new_n604_));
  AOI211_X1 g403(.A(KEYINPUT39), .B(new_n432_), .C1(new_n594_), .C2(new_n600_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n601_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n606_), .B(KEYINPUT40), .Z(G1325gat));
  NAND2_X1  g406(.A1(new_n594_), .A2(new_n403_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(G15gat), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(KEYINPUT101), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT101), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n608_), .A2(new_n611_), .A3(G15gat), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n610_), .A2(KEYINPUT41), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(G15gat), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n584_), .A2(new_n614_), .A3(new_n403_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(KEYINPUT41), .B1(new_n610_), .B2(new_n612_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n616_), .A2(new_n617_), .ZN(G1326gat));
  AOI21_X1  g417(.A(new_n341_), .B1(new_n594_), .B2(new_n402_), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n619_), .B(KEYINPUT42), .Z(new_n620_));
  NAND2_X1  g419(.A1(new_n402_), .A2(new_n341_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT102), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n584_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n620_), .A2(new_n623_), .ZN(G1327gat));
  NAND2_X1  g423(.A1(new_n479_), .A2(new_n581_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n625_), .A2(new_n541_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n453_), .A2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n627_), .A2(new_n417_), .A3(new_n326_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n585_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n590_), .A2(new_n479_), .A3(new_n592_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT43), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n631_), .B1(new_n582_), .B2(KEYINPUT103), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n581_), .A2(new_n571_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n568_), .A2(new_n569_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n576_), .A2(KEYINPUT70), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n633_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n632_), .B1(new_n405_), .B2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n379_), .A2(new_n383_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n326_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n638_), .A2(new_n598_), .A3(new_n599_), .A4(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n401_), .A2(new_n404_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n632_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n642_), .A2(new_n582_), .A3(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n630_), .B1(new_n637_), .B2(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n629_), .B1(new_n645_), .B2(KEYINPUT44), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n637_), .A2(new_n644_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n630_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n650_));
  AOI21_X1  g449(.A(KEYINPUT104), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT104), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n645_), .A2(new_n652_), .A3(KEYINPUT44), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n646_), .B1(new_n651_), .B2(new_n653_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n654_), .A2(KEYINPUT105), .A3(G29gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT105), .B1(new_n654_), .B2(G29gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n628_), .B1(new_n655_), .B2(new_n656_), .ZN(G1328gat));
  OR2_X1    g456(.A1(new_n600_), .A2(KEYINPUT106), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n600_), .A2(KEYINPUT106), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  AND4_X1   g459(.A1(new_n415_), .A2(new_n660_), .A3(new_n453_), .A4(new_n626_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT45), .Z(new_n662_));
  AOI21_X1  g461(.A(new_n288_), .B1(new_n645_), .B2(KEYINPUT44), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n652_), .B1(new_n645_), .B2(KEYINPUT44), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n649_), .A2(KEYINPUT104), .A3(new_n650_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n664_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  OAI211_X1 g466(.A(new_n662_), .B(KEYINPUT46), .C1(new_n667_), .C2(new_n415_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT46), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n666_), .A2(new_n665_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n415_), .B1(new_n670_), .B2(new_n663_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n661_), .B(KEYINPUT45), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n669_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n668_), .A2(new_n673_), .ZN(G1329gat));
  AOI21_X1  g473(.A(G43gat), .B1(new_n627_), .B2(new_n403_), .ZN(new_n675_));
  AOI211_X1 g474(.A(new_n358_), .B(new_n377_), .C1(new_n645_), .C2(KEYINPUT44), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n670_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT47), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n677_), .B(new_n678_), .ZN(G1330gat));
  AOI21_X1  g478(.A(G50gat), .B1(new_n627_), .B2(new_n402_), .ZN(new_n680_));
  AOI211_X1 g479(.A(new_n339_), .B(new_n356_), .C1(new_n645_), .C2(KEYINPUT44), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n670_), .B2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT107), .ZN(G1331gat));
  NOR2_X1   g482(.A1(new_n405_), .A2(new_n591_), .ZN(new_n684_));
  AND4_X1   g483(.A1(new_n636_), .A2(new_n684_), .A3(new_n478_), .A4(new_n541_), .ZN(new_n685_));
  AOI21_X1  g484(.A(G57gat), .B1(new_n685_), .B2(new_n585_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT108), .ZN(new_n687_));
  INV_X1    g486(.A(new_n581_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n479_), .A2(new_n540_), .A3(new_n591_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n642_), .A2(new_n688_), .A3(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT109), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n326_), .A2(G57gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n687_), .B1(new_n691_), .B2(new_n692_), .ZN(G1332gat));
  INV_X1    g492(.A(G64gat), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n685_), .A2(new_n694_), .A3(new_n660_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n691_), .A2(new_n660_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(G64gat), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n697_), .A2(KEYINPUT48), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n697_), .A2(KEYINPUT48), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n695_), .B1(new_n698_), .B2(new_n699_), .ZN(G1333gat));
  INV_X1    g499(.A(G71gat), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n685_), .A2(new_n701_), .A3(new_n403_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n691_), .A2(new_n403_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(G71gat), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n704_), .A2(KEYINPUT49), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(KEYINPUT49), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n702_), .B1(new_n705_), .B2(new_n706_), .ZN(G1334gat));
  INV_X1    g506(.A(G78gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n685_), .A2(new_n708_), .A3(new_n402_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n691_), .B2(new_n402_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n710_), .A2(new_n711_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n709_), .B1(new_n712_), .B2(new_n713_), .ZN(G1335gat));
  NAND3_X1  g513(.A1(new_n479_), .A2(new_n541_), .A3(new_n452_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n637_), .B2(new_n644_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G85gat), .B1(new_n717_), .B2(new_n639_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n625_), .A2(new_n540_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n684_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(new_n488_), .A3(new_n585_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n718_), .A2(new_n721_), .ZN(G1336gat));
  INV_X1    g521(.A(new_n660_), .ZN(new_n723_));
  OAI21_X1  g522(.A(G92gat), .B1(new_n717_), .B2(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n720_), .A2(new_n489_), .A3(new_n600_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(G1337gat));
  NAND4_X1  g525(.A1(new_n720_), .A2(new_n378_), .A3(new_n484_), .A4(new_n486_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT111), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n716_), .A2(new_n403_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(G99gat), .ZN(new_n730_));
  AOI211_X1 g529(.A(KEYINPUT111), .B(new_n496_), .C1(new_n716_), .C2(new_n403_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND2_X1  g532(.A1(new_n716_), .A2(new_n402_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(G106gat), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT52), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n684_), .A2(new_n485_), .A3(new_n402_), .A4(new_n719_), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n737_), .A2(KEYINPUT112), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(KEYINPUT112), .ZN(new_n739_));
  AOI22_X1  g538(.A1(new_n735_), .A2(new_n736_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n734_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n741_));
  XNOR2_X1  g540(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n740_), .A2(new_n741_), .A3(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1339gat));
  NAND3_X1  g544(.A1(new_n585_), .A2(new_n378_), .A3(new_n356_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n746_), .A2(new_n600_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n450_), .A2(new_n451_), .A3(new_n534_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT55), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n526_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n461_), .ZN(new_n752_));
  AOI21_X1  g551(.A(KEYINPUT12), .B1(new_n508_), .B2(new_n752_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n753_), .A2(new_n528_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n754_), .A2(KEYINPUT55), .A3(new_n517_), .A4(new_n514_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n514_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n525_), .A2(new_n518_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n516_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n751_), .A2(new_n755_), .A3(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n533_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT56), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n533_), .A2(new_n762_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n759_), .A2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n749_), .B1(new_n763_), .B2(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n443_), .A2(new_n447_), .A3(new_n410_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n445_), .A2(new_n446_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n438_), .A2(new_n442_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT114), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n438_), .A2(KEYINPUT114), .A3(new_n442_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n768_), .B1(new_n773_), .B2(new_n446_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n767_), .B1(new_n774_), .B2(new_n410_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n775_), .A2(new_n537_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n688_), .B1(new_n766_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT57), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n688_), .B(KEYINPUT57), .C1(new_n766_), .C2(new_n776_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n534_), .B(new_n767_), .C1(new_n774_), .C2(new_n410_), .ZN(new_n781_));
  AOI21_X1  g580(.A(KEYINPUT56), .B1(new_n759_), .B2(new_n760_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(new_n759_), .B2(new_n764_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n759_), .A2(new_n783_), .A3(new_n764_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n781_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n582_), .B1(new_n787_), .B2(KEYINPUT58), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n765_), .A2(KEYINPUT115), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n763_), .A2(new_n789_), .A3(new_n786_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n781_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT58), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n779_), .B(new_n780_), .C1(new_n788_), .C2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT116), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n787_), .A2(KEYINPUT58), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n792_), .A2(new_n793_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(new_n799_), .A3(new_n582_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n800_), .A2(KEYINPUT116), .A3(new_n780_), .A4(new_n779_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n797_), .A2(new_n479_), .A3(new_n801_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n636_), .A2(new_n478_), .A3(new_n452_), .A4(new_n540_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(KEYINPUT54), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n748_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(G113gat), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n806_), .A3(new_n591_), .ZN(new_n807_));
  XOR2_X1   g606(.A(new_n803_), .B(KEYINPUT54), .Z(new_n808_));
  OAI21_X1  g607(.A(new_n779_), .B1(new_n788_), .B2(new_n794_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n800_), .A2(KEYINPUT117), .A3(new_n779_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(new_n780_), .A3(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n808_), .B1(new_n813_), .B2(new_n479_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n748_), .A2(KEYINPUT59), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(KEYINPUT118), .B1(new_n814_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n818_));
  INV_X1    g617(.A(new_n780_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT58), .B1(new_n790_), .B2(new_n791_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n820_), .A2(new_n636_), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n821_), .A2(new_n798_), .B1(new_n778_), .B2(new_n777_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n819_), .B1(new_n822_), .B2(KEYINPUT117), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n478_), .B1(new_n823_), .B2(new_n811_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n818_), .B(new_n815_), .C1(new_n824_), .C2(new_n808_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n817_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n802_), .A2(new_n804_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n747_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT59), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n826_), .A2(new_n591_), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n807_), .B1(new_n831_), .B2(new_n806_), .ZN(G1340gat));
  INV_X1    g631(.A(KEYINPUT121), .ZN(new_n833_));
  XNOR2_X1  g632(.A(KEYINPUT119), .B(G120gat), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n540_), .B1(new_n828_), .B2(KEYINPUT59), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n826_), .B2(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n540_), .A2(KEYINPUT60), .ZN(new_n837_));
  MUX2_X1   g636(.A(KEYINPUT60), .B(new_n837_), .S(new_n834_), .Z(new_n838_));
  NAND3_X1  g637(.A1(new_n827_), .A2(new_n747_), .A3(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n839_), .B(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n833_), .B1(new_n836_), .B2(new_n841_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n839_), .B(KEYINPUT120), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n541_), .B1(new_n805_), .B2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n845_), .B1(new_n817_), .B2(new_n825_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n843_), .B(KEYINPUT121), .C1(new_n846_), .C2(new_n834_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n842_), .A2(new_n847_), .ZN(G1341gat));
  AOI21_X1  g647(.A(G127gat), .B1(new_n805_), .B2(new_n478_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n826_), .A2(new_n829_), .ZN(new_n850_));
  INV_X1    g649(.A(G127gat), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n851_), .B1(new_n478_), .B2(KEYINPUT122), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(KEYINPUT122), .B2(new_n851_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n849_), .B1(new_n850_), .B2(new_n853_), .ZN(G1342gat));
  INV_X1    g653(.A(G134gat), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n805_), .A2(new_n855_), .A3(new_n581_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n826_), .A2(new_n582_), .A3(new_n829_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n856_), .B1(new_n858_), .B2(new_n855_), .ZN(G1343gat));
  AOI21_X1  g658(.A(new_n383_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n860_), .A2(new_n585_), .A3(new_n723_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(new_n452_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT123), .B(G141gat), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(G1344gat));
  NOR2_X1   g663(.A1(new_n861_), .A2(new_n540_), .ZN(new_n865_));
  XOR2_X1   g664(.A(KEYINPUT124), .B(G148gat), .Z(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1345gat));
  NOR2_X1   g666(.A1(new_n861_), .A2(new_n479_), .ZN(new_n868_));
  XOR2_X1   g667(.A(KEYINPUT61), .B(G155gat), .Z(new_n869_));
  XNOR2_X1  g668(.A(new_n868_), .B(new_n869_), .ZN(G1346gat));
  OAI21_X1  g669(.A(G162gat), .B1(new_n861_), .B2(new_n636_), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n688_), .A2(G162gat), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n861_), .B2(new_n872_), .ZN(G1347gat));
  INV_X1    g672(.A(G169gat), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n585_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n660_), .A2(new_n356_), .A3(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n814_), .A2(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n874_), .B1(new_n877_), .B2(new_n591_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n879_), .A2(KEYINPUT125), .A3(new_n880_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n452_), .A2(new_n251_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(KEYINPUT126), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n877_), .A2(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n879_), .A2(KEYINPUT125), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT125), .ZN(new_n886_));
  OAI21_X1  g685(.A(KEYINPUT62), .B1(new_n878_), .B2(new_n886_), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n881_), .B(new_n884_), .C1(new_n885_), .C2(new_n887_), .ZN(G1348gat));
  AOI21_X1  g687(.A(G176gat), .B1(new_n877_), .B2(new_n541_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n402_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n890_));
  AND4_X1   g689(.A1(G176gat), .A2(new_n660_), .A3(new_n541_), .A4(new_n875_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n889_), .B1(new_n890_), .B2(new_n891_), .ZN(G1349gat));
  INV_X1    g691(.A(new_n877_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n893_), .A2(new_n221_), .A3(new_n479_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n890_), .A2(new_n478_), .A3(new_n660_), .A4(new_n875_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT127), .ZN(new_n896_));
  OR2_X1    g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  AOI21_X1  g696(.A(G183gat), .B1(new_n895_), .B2(new_n896_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n894_), .B1(new_n897_), .B2(new_n898_), .ZN(G1350gat));
  OAI21_X1  g698(.A(G190gat), .B1(new_n893_), .B2(new_n636_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n877_), .A2(new_n218_), .A3(new_n581_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(G1351gat));
  NAND3_X1  g701(.A1(new_n860_), .A2(new_n639_), .A3(new_n660_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n903_), .A2(new_n452_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(new_n203_), .ZN(G1352gat));
  NOR2_X1   g704(.A1(new_n903_), .A2(new_n540_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(new_n205_), .ZN(G1353gat));
  NOR2_X1   g706(.A1(new_n903_), .A2(new_n479_), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n908_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n909_));
  XOR2_X1   g708(.A(KEYINPUT63), .B(G211gat), .Z(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(new_n908_), .B2(new_n910_), .ZN(G1354gat));
  OAI21_X1  g710(.A(G218gat), .B1(new_n903_), .B2(new_n636_), .ZN(new_n912_));
  OR2_X1    g711(.A1(new_n688_), .A2(G218gat), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n903_), .B2(new_n913_), .ZN(G1355gat));
endmodule


