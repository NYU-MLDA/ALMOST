//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 1 0 0 0 0 1 1 0 1 0 0 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n646_, new_n647_, new_n648_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n808_, new_n809_, new_n810_, new_n812_, new_n813_, new_n814_,
    new_n816_, new_n817_, new_n818_, new_n820_, new_n821_, new_n823_,
    new_n824_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n856_, new_n857_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_;
  XNOR2_X1  g000(.A(G85gat), .B(G92gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT69), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT6), .ZN(new_n205_));
  OR3_X1    g004(.A1(KEYINPUT67), .A2(G99gat), .A3(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT7), .ZN(new_n207_));
  OR4_X1    g006(.A1(KEYINPUT67), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n205_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n203_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT70), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT8), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n211_), .B1(new_n210_), .B2(KEYINPUT68), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT10), .B(G99gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT66), .ZN(new_n216_));
  INV_X1    g015(.A(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT9), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n202_), .A2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(G85gat), .A3(G92gat), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n218_), .A2(new_n205_), .A3(new_n220_), .A4(new_n221_), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n214_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G57gat), .B(G64gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT11), .ZN(new_n225_));
  XOR2_X1   g024(.A(G71gat), .B(G78gat), .Z(new_n226_));
  OR2_X1    g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n224_), .A2(KEYINPUT11), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n225_), .A2(new_n226_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n227_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n223_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n223_), .A2(new_n230_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT71), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT12), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n232_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G230gat), .A2(G233gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT12), .B1(new_n233_), .B2(new_n234_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n237_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n240_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n243_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G120gat), .B(G148gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G176gat), .B(G204gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(KEYINPUT72), .B(KEYINPUT5), .Z(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT73), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n245_), .A2(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n242_), .A2(new_n244_), .A3(new_n250_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT74), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT74), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n252_), .A2(new_n256_), .A3(new_n253_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT13), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n258_), .A2(KEYINPUT13), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT27), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G8gat), .B(G36gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT18), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G64gat), .B(G92gat), .ZN(new_n267_));
  XOR2_X1   g066(.A(new_n266_), .B(new_n267_), .Z(new_n268_));
  INV_X1    g067(.A(G218gat), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n269_), .A2(G211gat), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n269_), .A2(G211gat), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT92), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G211gat), .B(G218gat), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT92), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n272_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT93), .ZN(new_n277_));
  OR2_X1    g076(.A1(G197gat), .A2(G204gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G197gat), .A2(G204gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT21), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n278_), .A2(KEYINPUT21), .A3(new_n279_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NOR3_X1   g083(.A1(new_n276_), .A2(new_n277_), .A3(new_n284_), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n282_), .A2(new_n283_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n272_), .A2(new_n275_), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT93), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  OAI22_X1  g087(.A1(new_n285_), .A2(new_n288_), .B1(new_n287_), .B2(new_n283_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G183gat), .A2(G190gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT23), .ZN(new_n291_));
  OR2_X1    g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(G176gat), .ZN(new_n296_));
  INV_X1    g095(.A(G169gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT83), .B1(new_n297_), .B2(KEYINPUT22), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT22), .B(G169gat), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n296_), .B(new_n298_), .C1(new_n299_), .C2(KEYINPUT83), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n295_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n297_), .A2(new_n296_), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n302_), .A2(KEYINPUT24), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n302_), .A2(KEYINPUT24), .A3(new_n294_), .ZN(new_n304_));
  AND3_X1   g103(.A1(new_n291_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT26), .B(G190gat), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT82), .ZN(new_n307_));
  INV_X1    g106(.A(G183gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT25), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT25), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n310_), .A2(KEYINPUT82), .A3(G183gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n306_), .A2(new_n309_), .A3(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n305_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n301_), .A2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT20), .B1(new_n289_), .B2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT96), .B(KEYINPUT24), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n316_), .A2(new_n297_), .A3(new_n296_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n291_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  XOR2_X1   g118(.A(KEYINPUT26), .B(G190gat), .Z(new_n320_));
  INV_X1    g119(.A(KEYINPUT95), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n310_), .A2(G183gat), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n308_), .A2(KEYINPUT25), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n321_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n308_), .A2(KEYINPUT25), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n310_), .A2(G183gat), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n325_), .A2(new_n326_), .A3(KEYINPUT95), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n320_), .B1(new_n324_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT97), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n302_), .A2(new_n294_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n330_), .A2(new_n316_), .ZN(new_n331_));
  NOR3_X1   g130(.A1(new_n328_), .A2(new_n329_), .A3(new_n331_), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n325_), .A2(new_n326_), .A3(KEYINPUT95), .ZN(new_n333_));
  AOI21_X1  g132(.A(KEYINPUT95), .B1(new_n325_), .B2(new_n326_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n306_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n331_), .ZN(new_n336_));
  AOI21_X1  g135(.A(KEYINPUT97), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n319_), .B1(new_n332_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT98), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  OAI211_X1 g139(.A(KEYINPUT98), .B(new_n319_), .C1(new_n332_), .C2(new_n337_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n299_), .A2(new_n296_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n293_), .A2(new_n294_), .A3(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n340_), .A2(new_n341_), .A3(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n315_), .B1(new_n344_), .B2(new_n289_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G226gat), .A2(G233gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT19), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT99), .B1(new_n345_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT99), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n287_), .A2(new_n283_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n277_), .B1(new_n276_), .B2(new_n284_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n286_), .A2(KEYINPUT93), .A3(new_n287_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n351_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n343_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n329_), .B1(new_n328_), .B2(new_n331_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n335_), .A2(new_n336_), .A3(KEYINPUT97), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n318_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n355_), .B1(new_n358_), .B2(KEYINPUT98), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n354_), .B1(new_n359_), .B2(new_n340_), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n350_), .B(new_n347_), .C1(new_n360_), .C2(new_n315_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n349_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n289_), .A2(KEYINPUT100), .A3(new_n314_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT100), .ZN(new_n364_));
  AOI22_X1  g163(.A1(new_n295_), .A2(new_n300_), .B1(new_n312_), .B2(new_n305_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n364_), .B1(new_n354_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n363_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n359_), .A2(new_n354_), .A3(new_n340_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT20), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n347_), .A2(new_n369_), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n367_), .A2(new_n368_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n268_), .B1(new_n362_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n268_), .ZN(new_n374_));
  AOI211_X1 g173(.A(new_n374_), .B(new_n371_), .C1(new_n349_), .C2(new_n361_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n264_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n362_), .A2(new_n268_), .A3(new_n372_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n289_), .A2(new_n355_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(new_n338_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n367_), .A2(new_n379_), .A3(KEYINPUT20), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n347_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n341_), .A2(new_n343_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n358_), .A2(KEYINPUT98), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n289_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n369_), .B1(new_n354_), .B2(new_n365_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n381_), .B1(new_n347_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n374_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n377_), .A2(new_n388_), .A3(KEYINPUT27), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n376_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(KEYINPUT84), .B(KEYINPUT30), .Z(new_n392_));
  XNOR2_X1  g191(.A(new_n314_), .B(new_n392_), .ZN(new_n393_));
  XOR2_X1   g192(.A(G71gat), .B(G99gat), .Z(new_n394_));
  NAND2_X1  g193(.A1(G227gat), .A2(G233gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G15gat), .B(G43gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT85), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n396_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n393_), .B(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n400_), .A2(KEYINPUT87), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G127gat), .B(G134gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G113gat), .B(G120gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  XOR2_X1   g203(.A(KEYINPUT86), .B(KEYINPUT31), .Z(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n401_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n400_), .A2(KEYINPUT87), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n400_), .A2(KEYINPUT87), .A3(new_n406_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G225gat), .A2(G233gat), .ZN(new_n412_));
  XOR2_X1   g211(.A(G141gat), .B(G148gat), .Z(new_n413_));
  NAND2_X1  g212(.A1(G155gat), .A2(G162gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT89), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT89), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n416_), .A2(G155gat), .A3(G162gat), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT1), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n415_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  OR3_X1    g218(.A1(KEYINPUT88), .A2(G155gat), .A3(G162gat), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT88), .B1(G155gat), .B2(G162gat), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n419_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n418_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n413_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  OR3_X1    g223(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G141gat), .A2(G148gat), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT2), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n425_), .A2(new_n428_), .A3(new_n429_), .A4(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n415_), .A2(new_n417_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n431_), .A2(new_n432_), .A3(new_n420_), .A4(new_n421_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n424_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT90), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT101), .ZN(new_n437_));
  INV_X1    g236(.A(new_n404_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n424_), .A2(KEYINPUT90), .A3(new_n433_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .A4(new_n439_), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n424_), .A2(KEYINPUT90), .A3(new_n433_), .ZN(new_n441_));
  AOI21_X1  g240(.A(KEYINPUT90), .B1(new_n424_), .B2(new_n433_), .ZN(new_n442_));
  NOR3_X1   g241(.A1(new_n441_), .A2(new_n442_), .A3(new_n404_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n437_), .B1(new_n434_), .B2(new_n438_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  OAI211_X1 g244(.A(KEYINPUT4), .B(new_n440_), .C1(new_n443_), .C2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n436_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n447_), .A2(KEYINPUT4), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n412_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  XOR2_X1   g248(.A(G1gat), .B(G29gat), .Z(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT0), .ZN(new_n451_));
  XOR2_X1   g250(.A(new_n451_), .B(KEYINPUT102), .Z(new_n452_));
  XNOR2_X1  g251(.A(G57gat), .B(G85gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n412_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n447_), .A2(new_n444_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n455_), .B1(new_n456_), .B2(new_n440_), .ZN(new_n457_));
  OR3_X1    g256(.A1(new_n449_), .A2(new_n454_), .A3(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n454_), .B1(new_n449_), .B2(new_n457_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n411_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT94), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT29), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n463_), .B1(new_n424_), .B2(new_n433_), .ZN(new_n464_));
  OAI211_X1 g263(.A(G228gat), .B(G233gat), .C1(new_n354_), .C2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G78gat), .B(G106gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NOR3_X1   g266(.A1(new_n441_), .A2(new_n442_), .A3(new_n463_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G228gat), .A2(G233gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n289_), .A2(new_n469_), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n465_), .B(new_n467_), .C1(new_n468_), .C2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n436_), .A2(KEYINPUT29), .A3(new_n439_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(new_n469_), .A3(new_n289_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n467_), .B1(new_n474_), .B2(new_n465_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n462_), .B1(new_n472_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n465_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(new_n466_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(KEYINPUT94), .A3(new_n471_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n463_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n480_));
  XOR2_X1   g279(.A(G22gat), .B(G50gat), .Z(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n463_), .B(new_n481_), .C1(new_n441_), .C2(new_n442_), .ZN(new_n484_));
  XOR2_X1   g283(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  AND3_X1   g285(.A1(new_n483_), .A2(new_n484_), .A3(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n486_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n476_), .A2(new_n479_), .A3(new_n489_), .ZN(new_n490_));
  OAI221_X1 g289(.A(new_n462_), .B1(new_n487_), .B2(new_n488_), .C1(new_n472_), .C2(new_n475_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n391_), .A2(new_n461_), .A3(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(new_n493_), .B(KEYINPUT107), .Z(new_n494_));
  NOR2_X1   g293(.A1(new_n492_), .A2(new_n460_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n376_), .A2(new_n495_), .A3(new_n389_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT105), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n376_), .A2(new_n495_), .A3(KEYINPUT105), .A4(new_n389_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n492_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n459_), .A2(KEYINPUT33), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT33), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n502_), .B(new_n454_), .C1(new_n449_), .C2(new_n457_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n350_), .B1(new_n386_), .B2(new_n347_), .ZN(new_n505_));
  AOI211_X1 g304(.A(KEYINPUT99), .B(new_n348_), .C1(new_n384_), .C2(new_n385_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n372_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(new_n374_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n446_), .A2(new_n412_), .A3(new_n448_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n454_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT103), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n456_), .A2(new_n455_), .A3(new_n440_), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n511_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n509_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n504_), .A2(new_n508_), .A3(new_n377_), .A4(new_n515_), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n268_), .A2(KEYINPUT32), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n387_), .A2(new_n517_), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n460_), .B(new_n518_), .C1(new_n517_), .C2(new_n507_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n500_), .B1(new_n516_), .B2(new_n519_), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n498_), .B(new_n499_), .C1(KEYINPUT104), .C2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(KEYINPUT104), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n411_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT106), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  OAI211_X1 g325(.A(KEYINPUT106), .B(new_n411_), .C1(new_n521_), .C2(new_n523_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n494_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G29gat), .B(G36gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G43gat), .B(G50gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(KEYINPUT75), .B(KEYINPUT15), .Z(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(G1gat), .ZN(new_n534_));
  INV_X1    g333(.A(G8gat), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT14), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(G22gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(G15gat), .ZN(new_n538_));
  INV_X1    g337(.A(G15gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(G22gat), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n536_), .A2(new_n538_), .A3(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT80), .ZN(new_n542_));
  XOR2_X1   g341(.A(G1gat), .B(G8gat), .Z(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(new_n544_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  MUX2_X1   g346(.A(new_n533_), .B(new_n531_), .S(new_n547_), .Z(new_n548_));
  NAND2_X1  g347(.A1(G229gat), .A2(G233gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n547_), .B(new_n531_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n550_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G113gat), .B(G141gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G169gat), .B(G197gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n552_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n552_), .A2(new_n556_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n559_), .B(KEYINPUT81), .Z(new_n560_));
  NOR3_X1   g359(.A1(new_n263_), .A2(new_n528_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n223_), .A2(new_n531_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT76), .ZN(new_n563_));
  INV_X1    g362(.A(new_n223_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT35), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G232gat), .A2(G233gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT34), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  AOI22_X1  g367(.A1(new_n564_), .A2(new_n533_), .B1(new_n565_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n563_), .A2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n568_), .A2(new_n565_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n570_), .A2(new_n571_), .ZN(new_n573_));
  XOR2_X1   g372(.A(G190gat), .B(G218gat), .Z(new_n574_));
  XNOR2_X1  g373(.A(G134gat), .B(G162gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT36), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT77), .ZN(new_n579_));
  OR3_X1    g378(.A1(new_n572_), .A2(new_n573_), .A3(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n576_), .B(new_n577_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT79), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n582_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n580_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT37), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT78), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n585_), .B1(new_n583_), .B2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n584_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n547_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G231gat), .A2(G233gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n230_), .B(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n590_), .B(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT17), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G127gat), .B(G155gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT16), .ZN(new_n597_));
  XOR2_X1   g396(.A(G183gat), .B(G211gat), .Z(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n594_), .B1(new_n595_), .B2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n595_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n593_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n589_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n561_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT108), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n561_), .A2(KEYINPUT108), .A3(new_n605_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n460_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n611_), .A2(G1gat), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n584_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n528_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n559_), .ZN(new_n616_));
  NOR4_X1   g415(.A1(new_n260_), .A2(new_n261_), .A3(new_n604_), .A4(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(G1gat), .B1(new_n618_), .B2(new_n611_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n619_), .A2(KEYINPUT38), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n608_), .A2(KEYINPUT38), .A3(new_n609_), .A4(new_n612_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT109), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n621_), .A2(new_n622_), .ZN(new_n624_));
  OAI22_X1  g423(.A1(new_n613_), .A2(new_n620_), .B1(new_n623_), .B2(new_n624_), .ZN(G1324gat));
  NAND3_X1  g424(.A1(new_n615_), .A2(new_n390_), .A3(new_n617_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(G8gat), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT110), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT110), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n626_), .A2(new_n629_), .A3(G8gat), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n628_), .A2(KEYINPUT39), .A3(new_n630_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n608_), .A2(new_n535_), .A3(new_n390_), .A4(new_n609_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n633_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT40), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n633_), .A2(new_n635_), .A3(KEYINPUT40), .A4(new_n634_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(G1325gat));
  INV_X1    g439(.A(new_n411_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n610_), .A2(new_n539_), .A3(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G15gat), .B1(new_n618_), .B2(new_n411_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT41), .Z(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(G1326gat));
  NAND3_X1  g444(.A1(new_n610_), .A2(new_n537_), .A3(new_n500_), .ZN(new_n646_));
  OAI21_X1  g445(.A(G22gat), .B1(new_n618_), .B2(new_n492_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT42), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(G1327gat));
  NOR2_X1   g448(.A1(new_n584_), .A2(new_n603_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n561_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(G29gat), .B1(new_n652_), .B2(new_n460_), .ZN(new_n653_));
  OAI21_X1  g452(.A(KEYINPUT43), .B1(new_n528_), .B2(new_n588_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n493_), .B(KEYINPUT107), .ZN(new_n655_));
  INV_X1    g454(.A(new_n527_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n516_), .A2(new_n519_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(new_n492_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT104), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n660_), .A2(new_n522_), .A3(new_n498_), .A4(new_n499_), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT106), .B1(new_n661_), .B2(new_n411_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n655_), .B1(new_n656_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n663_), .A2(new_n664_), .A3(new_n589_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n654_), .A2(new_n665_), .ZN(new_n666_));
  NOR4_X1   g465(.A1(new_n260_), .A2(new_n261_), .A3(new_n603_), .A4(new_n616_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n666_), .A2(KEYINPUT44), .A3(new_n667_), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n668_), .A2(G29gat), .A3(new_n460_), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n528_), .A2(KEYINPUT43), .A3(new_n588_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n664_), .B1(new_n663_), .B2(new_n589_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n667_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n653_), .B1(new_n669_), .B2(new_n674_), .ZN(G1328gat));
  INV_X1    g474(.A(G36gat), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n668_), .A2(new_n390_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n677_), .B2(new_n674_), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n391_), .A2(KEYINPUT111), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n391_), .A2(KEYINPUT111), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n561_), .A2(new_n676_), .A3(new_n650_), .A4(new_n681_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT45), .Z(new_n683_));
  NOR2_X1   g482(.A1(new_n678_), .A2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT46), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT46), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n686_), .B1(new_n678_), .B2(new_n683_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(G1329gat));
  XOR2_X1   g487(.A(KEYINPUT113), .B(KEYINPUT47), .Z(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(G43gat), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n411_), .A2(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n674_), .A2(new_n668_), .A3(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT112), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT112), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n674_), .A2(new_n695_), .A3(new_n668_), .A4(new_n692_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n561_), .A2(new_n641_), .A3(new_n650_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(new_n691_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n690_), .B1(new_n697_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n699_), .ZN(new_n701_));
  AOI211_X1 g500(.A(new_n701_), .B(new_n689_), .C1(new_n694_), .C2(new_n696_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n700_), .A2(new_n702_), .ZN(G1330gat));
  OR3_X1    g502(.A1(new_n651_), .A2(G50gat), .A3(new_n492_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n674_), .A2(new_n500_), .A3(new_n668_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT114), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n705_), .A2(new_n706_), .A3(G50gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n705_), .B2(G50gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n704_), .B1(new_n707_), .B2(new_n708_), .ZN(G1331gat));
  NOR3_X1   g508(.A1(new_n528_), .A2(new_n262_), .A3(new_n559_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(new_n605_), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT115), .Z(new_n712_));
  AOI21_X1  g511(.A(G57gat), .B1(new_n712_), .B2(new_n460_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n560_), .A2(new_n603_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n262_), .A2(new_n714_), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n615_), .A2(new_n715_), .A3(G57gat), .A4(new_n460_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT116), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n713_), .A2(new_n717_), .ZN(G1332gat));
  INV_X1    g517(.A(G64gat), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n712_), .A2(new_n719_), .A3(new_n681_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n615_), .A2(new_n715_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n681_), .ZN(new_n722_));
  OAI21_X1  g521(.A(G64gat), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT48), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n720_), .A2(new_n724_), .ZN(G1333gat));
  INV_X1    g524(.A(G71gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n712_), .A2(new_n726_), .A3(new_n641_), .ZN(new_n727_));
  OAI21_X1  g526(.A(G71gat), .B1(new_n721_), .B2(new_n411_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT49), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1334gat));
  INV_X1    g529(.A(G78gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n712_), .A2(new_n731_), .A3(new_n500_), .ZN(new_n732_));
  OAI21_X1  g531(.A(G78gat), .B1(new_n721_), .B2(new_n492_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT50), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(G1335gat));
  NOR3_X1   g534(.A1(new_n262_), .A2(new_n603_), .A3(new_n559_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n666_), .A2(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(G85gat), .B1(new_n737_), .B2(new_n611_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n710_), .A2(new_n650_), .ZN(new_n739_));
  INV_X1    g538(.A(G85gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(new_n740_), .A3(new_n460_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n738_), .A2(new_n741_), .ZN(G1336gat));
  OAI21_X1  g541(.A(G92gat), .B1(new_n737_), .B2(new_n722_), .ZN(new_n743_));
  INV_X1    g542(.A(G92gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n739_), .A2(new_n744_), .A3(new_n390_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1337gat));
  NAND3_X1  g545(.A1(new_n739_), .A2(new_n216_), .A3(new_n641_), .ZN(new_n747_));
  OAI21_X1  g546(.A(G99gat), .B1(new_n737_), .B2(new_n411_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g549(.A1(new_n739_), .A2(new_n217_), .A3(new_n500_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n666_), .A2(new_n500_), .A3(new_n736_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n752_), .A2(new_n753_), .A3(G106gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n752_), .B2(G106gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT53), .ZN(G1339gat));
  AND2_X1   g556(.A1(new_n237_), .A2(new_n241_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(KEYINPUT55), .A3(new_n240_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT55), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n242_), .A2(new_n760_), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n759_), .B(new_n761_), .C1(new_n240_), .C2(new_n758_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n251_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT56), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n762_), .A2(KEYINPUT56), .A3(new_n251_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n253_), .A2(new_n559_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT118), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n551_), .A2(new_n549_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n771_), .B(new_n555_), .C1(new_n548_), .C2(new_n549_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n558_), .B1(new_n772_), .B2(KEYINPUT119), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n773_), .B1(KEYINPUT119), .B2(new_n772_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n255_), .A2(new_n257_), .A3(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n614_), .B1(new_n770_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n253_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n777_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT58), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n589_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n778_), .A2(KEYINPUT58), .ZN(new_n781_));
  OAI22_X1  g580(.A1(new_n776_), .A2(KEYINPUT57), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n776_), .A2(KEYINPUT57), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n604_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n785_));
  XOR2_X1   g584(.A(new_n714_), .B(KEYINPUT117), .Z(new_n786_));
  NAND3_X1  g585(.A1(new_n262_), .A2(new_n588_), .A3(new_n786_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT54), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n785_), .A2(new_n788_), .ZN(new_n789_));
  NOR4_X1   g588(.A1(new_n390_), .A2(new_n411_), .A3(new_n500_), .A4(new_n611_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(G113gat), .B1(new_n792_), .B2(new_n559_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT59), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n791_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n789_), .A2(KEYINPUT59), .A3(new_n790_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  XOR2_X1   g596(.A(KEYINPUT120), .B(G113gat), .Z(new_n798_));
  NOR2_X1   g597(.A1(new_n560_), .A2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n793_), .B1(new_n797_), .B2(new_n799_), .ZN(G1340gat));
  INV_X1    g599(.A(KEYINPUT60), .ZN(new_n801_));
  INV_X1    g600(.A(G120gat), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n263_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n803_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n792_), .A2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n262_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(new_n802_), .ZN(G1341gat));
  INV_X1    g606(.A(G127gat), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n792_), .A2(new_n808_), .A3(new_n603_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n604_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(new_n808_), .ZN(G1342gat));
  INV_X1    g610(.A(G134gat), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n792_), .A2(new_n812_), .A3(new_n614_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n588_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(new_n812_), .ZN(G1343gat));
  NAND4_X1  g614(.A1(new_n722_), .A2(new_n411_), .A3(new_n500_), .A4(new_n460_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n816_), .B1(new_n785_), .B2(new_n788_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n559_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n263_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(KEYINPUT121), .B(G148gat), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n820_), .B(new_n821_), .ZN(G1345gat));
  NAND2_X1  g621(.A1(new_n817_), .A2(new_n603_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(KEYINPUT61), .B(G155gat), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n823_), .B(new_n824_), .ZN(G1346gat));
  INV_X1    g624(.A(G162gat), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n817_), .A2(new_n826_), .A3(new_n614_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n826_), .B1(new_n817_), .B2(new_n589_), .ZN(new_n829_));
  OAI21_X1  g628(.A(KEYINPUT122), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT122), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n817_), .A2(new_n589_), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n831_), .B(new_n827_), .C1(new_n832_), .C2(new_n826_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n830_), .A2(new_n833_), .ZN(G1347gat));
  INV_X1    g633(.A(KEYINPUT62), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n681_), .A2(new_n492_), .A3(new_n461_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n789_), .A2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n838_), .A2(new_n616_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n835_), .B1(new_n839_), .B2(new_n297_), .ZN(new_n840_));
  OAI211_X1 g639(.A(KEYINPUT62), .B(G169gat), .C1(new_n838_), .C2(new_n616_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n299_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n840_), .A2(new_n841_), .A3(new_n842_), .ZN(G1348gat));
  NOR2_X1   g642(.A1(new_n838_), .A2(new_n262_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(new_n296_), .ZN(G1349gat));
  NAND2_X1  g644(.A1(new_n324_), .A2(new_n327_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n789_), .A2(new_n603_), .A3(new_n846_), .A4(new_n837_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT123), .ZN(new_n848_));
  AOI211_X1 g647(.A(new_n604_), .B(new_n836_), .C1(new_n785_), .C2(new_n788_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n847_), .B(new_n848_), .C1(new_n849_), .C2(new_n308_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n789_), .A2(new_n603_), .A3(new_n837_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(G183gat), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n848_), .B1(new_n853_), .B2(new_n847_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n851_), .A2(new_n854_), .ZN(G1350gat));
  OAI21_X1  g654(.A(G190gat), .B1(new_n838_), .B2(new_n588_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n614_), .A2(new_n306_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n838_), .B2(new_n857_), .ZN(G1351gat));
  NAND2_X1  g657(.A1(new_n411_), .A2(new_n495_), .ZN(new_n859_));
  XOR2_X1   g658(.A(new_n859_), .B(KEYINPUT124), .Z(new_n860_));
  NAND2_X1  g659(.A1(new_n681_), .A2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n861_), .B1(new_n785_), .B2(new_n788_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n559_), .ZN(new_n863_));
  XOR2_X1   g662(.A(KEYINPUT125), .B(G197gat), .Z(new_n864_));
  XNOR2_X1  g663(.A(new_n863_), .B(new_n864_), .ZN(G1352gat));
  NAND2_X1  g664(.A1(new_n862_), .A2(new_n263_), .ZN(new_n866_));
  INV_X1    g665(.A(G204gat), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(KEYINPUT126), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n866_), .B(new_n868_), .ZN(G1353gat));
  INV_X1    g668(.A(new_n862_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n870_), .A2(new_n604_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n872_));
  AND2_X1   g671(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n871_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n874_), .B1(new_n871_), .B2(new_n872_), .ZN(G1354gat));
  INV_X1    g674(.A(KEYINPUT127), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n862_), .A2(new_n269_), .A3(new_n614_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n269_), .B1(new_n862_), .B2(new_n589_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n876_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n879_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n881_), .A2(KEYINPUT127), .A3(new_n877_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(G1355gat));
endmodule


