//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 1 1 1 1 0 1 0 1 0 0 0 1 0 1 1 1 0 1 1 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n894_, new_n896_, new_n897_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT65), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G85gat), .B(G92gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT9), .ZN(new_n206_));
  XOR2_X1   g005(.A(KEYINPUT10), .B(G99gat), .Z(new_n207_));
  INV_X1    g006(.A(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT9), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(G85gat), .A3(G92gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT6), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n206_), .A2(new_n209_), .A3(new_n211_), .A4(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  NOR3_X1   g018(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  AOI211_X1 g020(.A(KEYINPUT8), .B(new_n204_), .C1(new_n221_), .C2(new_n216_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT8), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT7), .ZN(new_n224_));
  INV_X1    g023(.A(G99gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(new_n225_), .A3(new_n208_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n214_), .B1(G99gat), .B2(G106gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n228_));
  OAI211_X1 g027(.A(new_n218_), .B(new_n226_), .C1(new_n227_), .C2(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n223_), .B1(new_n229_), .B2(new_n205_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n217_), .B1(new_n222_), .B2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G57gat), .B(G64gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT11), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT11), .ZN(new_n234_));
  INV_X1    g033(.A(G57gat), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n235_), .A2(G64gat), .ZN(new_n236_));
  INV_X1    g035(.A(G64gat), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n237_), .A2(G57gat), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n234_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n233_), .A2(new_n239_), .ZN(new_n240_));
  AND2_X1   g039(.A1(KEYINPUT64), .A2(G71gat), .ZN(new_n241_));
  NOR2_X1   g040(.A1(KEYINPUT64), .A2(G71gat), .ZN(new_n242_));
  NOR3_X1   g041(.A1(new_n241_), .A2(new_n242_), .A3(G78gat), .ZN(new_n243_));
  INV_X1    g042(.A(G78gat), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT64), .ZN(new_n245_));
  INV_X1    g044(.A(G71gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(KEYINPUT64), .A2(G71gat), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n244_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n243_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n240_), .A2(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(G78gat), .B1(new_n241_), .B2(new_n242_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n247_), .A2(new_n244_), .A3(new_n248_), .ZN(new_n253_));
  AOI22_X1  g052(.A1(new_n252_), .A2(new_n253_), .B1(new_n232_), .B2(KEYINPUT11), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n251_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n231_), .A2(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n254_), .B1(new_n240_), .B2(new_n250_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n258_), .B(new_n217_), .C1(new_n230_), .C2(new_n222_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n257_), .A2(KEYINPUT12), .A3(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT12), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n231_), .A2(new_n261_), .A3(new_n256_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G230gat), .A2(G233gat), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n203_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n264_), .ZN(new_n266_));
  AOI211_X1 g065(.A(KEYINPUT65), .B(new_n266_), .C1(new_n260_), .C2(new_n262_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n264_), .B1(new_n257_), .B2(new_n259_), .ZN(new_n268_));
  NOR3_X1   g067(.A1(new_n265_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT66), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G120gat), .B(G148gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT5), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G176gat), .B(G204gat), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n272_), .B(new_n273_), .Z(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NOR3_X1   g074(.A1(new_n269_), .A2(new_n270_), .A3(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n263_), .A2(new_n264_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT65), .ZN(new_n278_));
  INV_X1    g077(.A(new_n268_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n266_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(new_n203_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n278_), .A2(new_n279_), .A3(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT66), .B1(new_n282_), .B2(new_n274_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n276_), .A2(new_n283_), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n278_), .A2(new_n279_), .A3(new_n281_), .A4(new_n275_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT67), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n265_), .A2(new_n267_), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n288_), .A2(KEYINPUT67), .A3(new_n279_), .A4(new_n275_), .ZN(new_n289_));
  AND2_X1   g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n202_), .B1(new_n284_), .B2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n270_), .B1(new_n269_), .B2(new_n275_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n282_), .A2(KEYINPUT66), .A3(new_n274_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n287_), .A2(new_n289_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(KEYINPUT13), .A3(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n291_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G29gat), .B(G36gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G43gat), .B(G50gat), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n299_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT74), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G15gat), .B(G22gat), .ZN(new_n305_));
  INV_X1    g104(.A(G1gat), .ZN(new_n306_));
  INV_X1    g105(.A(G8gat), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT14), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n305_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G1gat), .B(G8gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n304_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT75), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n304_), .A2(new_n312_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n316_), .A2(G229gat), .A3(G233gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n302_), .B(KEYINPUT15), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(new_n311_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G229gat), .A2(G233gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT76), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n313_), .A2(new_n319_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n317_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G113gat), .B(G141gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G169gat), .B(G197gat), .ZN(new_n325_));
  XOR2_X1   g124(.A(new_n324_), .B(new_n325_), .Z(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n323_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n317_), .A2(new_n322_), .A3(new_n326_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n297_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G227gat), .A2(G233gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(G71gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(new_n225_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G15gat), .B(G43gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT82), .B(KEYINPUT83), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n336_), .B(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT81), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT77), .ZN(new_n342_));
  INV_X1    g141(.A(G190gat), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n342_), .B1(new_n343_), .B2(KEYINPUT26), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT25), .B(G183gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT26), .B(G190gat), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n344_), .B(new_n345_), .C1(new_n346_), .C2(new_n342_), .ZN(new_n347_));
  INV_X1    g146(.A(G169gat), .ZN(new_n348_));
  INV_X1    g147(.A(G176gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n350_), .A2(KEYINPUT24), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n347_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G169gat), .A2(G176gat), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n350_), .A2(KEYINPUT24), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n350_), .A2(KEYINPUT78), .A3(KEYINPUT24), .A4(new_n353_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT23), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n359_), .B1(G183gat), .B2(G190gat), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n359_), .A2(G183gat), .A3(G190gat), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT79), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n359_), .A2(KEYINPUT79), .A3(G183gat), .A4(G190gat), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n360_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NOR3_X1   g164(.A1(new_n352_), .A2(new_n358_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n348_), .A2(KEYINPUT22), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT22), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(G169gat), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n367_), .A2(new_n369_), .A3(new_n349_), .ZN(new_n370_));
  AND3_X1   g169(.A1(new_n370_), .A2(KEYINPUT80), .A3(new_n353_), .ZN(new_n371_));
  AOI21_X1  g170(.A(KEYINPUT80), .B1(new_n370_), .B2(new_n353_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(G183gat), .A2(G190gat), .ZN(new_n373_));
  INV_X1    g172(.A(G183gat), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT23), .B1(new_n374_), .B2(new_n343_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n373_), .B1(new_n375_), .B2(new_n361_), .ZN(new_n376_));
  NOR3_X1   g175(.A1(new_n371_), .A2(new_n372_), .A3(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n341_), .B1(new_n366_), .B2(new_n377_), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n356_), .A2(new_n357_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n365_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n379_), .A2(new_n380_), .A3(new_n351_), .A4(new_n347_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n372_), .A2(new_n376_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n371_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n381_), .A2(new_n384_), .A3(KEYINPUT81), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n378_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT30), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n340_), .B1(new_n387_), .B2(KEYINPUT84), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(KEYINPUT84), .ZN(new_n389_));
  XOR2_X1   g188(.A(new_n388_), .B(new_n389_), .Z(new_n390_));
  XNOR2_X1  g189(.A(G127gat), .B(G134gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G113gat), .B(G120gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT85), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT31), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  OR2_X1    g195(.A1(new_n390_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n390_), .A2(new_n396_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G228gat), .A2(G233gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(new_n244_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(new_n208_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G22gat), .B(G50gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  OR2_X1    g205(.A1(G197gat), .A2(G204gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G197gat), .A2(G204gat), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(KEYINPUT21), .A3(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G211gat), .B(G218gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT90), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n407_), .A2(new_n408_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT21), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n411_), .B1(new_n412_), .B2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n413_), .A2(KEYINPUT90), .A3(new_n414_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n409_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n410_), .ZN(new_n419_));
  AOI22_X1  g218(.A1(new_n416_), .A2(new_n417_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G155gat), .A2(G162gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT87), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT87), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n424_), .A2(G155gat), .A3(G162gat), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(G155gat), .ZN(new_n428_));
  INV_X1    g227(.A(G162gat), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(new_n429_), .A3(KEYINPUT86), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT86), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n431_), .B1(G155gat), .B2(G162gat), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  OR3_X1    g232(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT2), .ZN(new_n435_));
  INV_X1    g234(.A(G141gat), .ZN(new_n436_));
  INV_X1    g235(.A(G148gat), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n435_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n434_), .A2(new_n438_), .A3(new_n439_), .A4(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n427_), .A2(new_n433_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT88), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT1), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n444_), .B(new_n433_), .C1(new_n426_), .C2(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n445_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n430_), .A2(new_n432_), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT88), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n426_), .A2(new_n445_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n446_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  XOR2_X1   g250(.A(G141gat), .B(G148gat), .Z(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT89), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT89), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n451_), .A2(new_n455_), .A3(new_n452_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n443_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT29), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n421_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n451_), .A2(new_n455_), .A3(new_n452_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n455_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n442_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT28), .B1(new_n462_), .B2(KEYINPUT29), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT28), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n457_), .A2(new_n464_), .A3(new_n458_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n459_), .A2(new_n463_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n459_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n406_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n463_), .A2(new_n465_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n459_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n472_), .A2(new_n466_), .A3(new_n405_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n469_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT96), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT93), .B1(new_n457_), .B2(new_n394_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n457_), .A2(new_n393_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT93), .ZN(new_n478_));
  INV_X1    g277(.A(new_n394_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n462_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n476_), .A2(KEYINPUT4), .A3(new_n477_), .A4(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G225gat), .A2(G233gat), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n457_), .A2(new_n394_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT4), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n483_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n481_), .A2(new_n486_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n476_), .A2(new_n483_), .A3(new_n477_), .A4(new_n480_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G1gat), .B(G29gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(G85gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT0), .B(G57gat), .ZN(new_n491_));
  XOR2_X1   g290(.A(new_n490_), .B(new_n491_), .Z(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n488_), .A2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n475_), .B1(new_n487_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n481_), .A2(new_n486_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n496_), .A2(KEYINPUT96), .A3(new_n493_), .A4(new_n488_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n378_), .A2(new_n385_), .A3(new_n420_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT20), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n353_), .B(new_n370_), .C1(new_n365_), .C2(new_n373_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n346_), .A2(new_n345_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n375_), .A2(new_n361_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n501_), .A2(new_n502_), .A3(new_n351_), .A4(new_n354_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n500_), .A2(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n499_), .B1(new_n421_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n498_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G226gat), .A2(G233gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT19), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  NOR3_X1   g308(.A1(new_n366_), .A2(new_n341_), .A3(new_n377_), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT81), .B1(new_n381_), .B2(new_n384_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n421_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n415_), .A2(new_n412_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n513_), .A2(new_n417_), .A3(new_n409_), .A4(new_n410_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n418_), .A2(new_n419_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n514_), .A2(new_n500_), .A3(new_n515_), .A4(new_n503_), .ZN(new_n516_));
  AOI211_X1 g315(.A(new_n499_), .B(new_n508_), .C1(new_n516_), .C2(KEYINPUT91), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT91), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n420_), .A2(new_n518_), .A3(new_n500_), .A4(new_n503_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n512_), .A2(new_n517_), .A3(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G8gat), .B(G36gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT18), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G64gat), .B(G92gat), .ZN(new_n523_));
  XOR2_X1   g322(.A(new_n522_), .B(new_n523_), .Z(new_n524_));
  NAND3_X1  g323(.A1(new_n509_), .A2(new_n520_), .A3(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n524_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n516_), .A2(KEYINPUT91), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n508_), .A2(new_n499_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n519_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n420_), .B1(new_n378_), .B2(new_n385_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n508_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n532_), .B1(new_n498_), .B2(new_n505_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n526_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n525_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT92), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT92), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n525_), .A2(new_n534_), .A3(new_n537_), .ZN(new_n538_));
  AOI22_X1  g337(.A1(new_n495_), .A2(new_n497_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n482_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n481_), .A2(new_n540_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n476_), .A2(new_n482_), .A3(new_n477_), .A4(new_n480_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n541_), .A2(new_n542_), .A3(new_n492_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT95), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT33), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n541_), .A2(KEYINPUT95), .A3(new_n542_), .A4(new_n492_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n545_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n493_), .A2(new_n546_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n541_), .A2(new_n542_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT94), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n541_), .A2(KEYINPUT94), .A3(new_n542_), .A4(new_n549_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n539_), .A2(new_n548_), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n492_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(new_n543_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n524_), .A2(KEYINPUT32), .ZN(new_n559_));
  NOR3_X1   g358(.A1(new_n531_), .A2(new_n533_), .A3(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n516_), .A2(KEYINPUT97), .A3(KEYINPUT20), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n516_), .A2(KEYINPUT20), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT97), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n512_), .A2(new_n561_), .A3(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(new_n508_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n566_), .B1(new_n508_), .B2(new_n506_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n560_), .B1(new_n567_), .B2(new_n559_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n558_), .A2(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n474_), .B1(new_n555_), .B2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n524_), .B(KEYINPUT98), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n567_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n525_), .A2(KEYINPUT27), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT27), .ZN(new_n577_));
  AOI21_X1  g376(.A(KEYINPUT99), .B1(new_n535_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT99), .ZN(new_n579_));
  AOI211_X1 g378(.A(new_n579_), .B(KEYINPUT27), .C1(new_n525_), .C2(new_n534_), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n474_), .B(new_n576_), .C1(new_n578_), .C2(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(KEYINPUT100), .B1(new_n581_), .B2(new_n558_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n574_), .B1(new_n567_), .B2(new_n572_), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n531_), .A2(new_n533_), .A3(new_n526_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n524_), .B1(new_n509_), .B2(new_n520_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n577_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(new_n579_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n535_), .A2(KEYINPUT99), .A3(new_n577_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n583_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT100), .ZN(new_n590_));
  INV_X1    g389(.A(new_n543_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n591_), .A2(new_n556_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n589_), .A2(new_n590_), .A3(new_n592_), .A4(new_n474_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n582_), .A2(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n400_), .B1(new_n570_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n474_), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n399_), .A2(new_n592_), .A3(new_n596_), .A4(new_n589_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n333_), .B1(new_n595_), .B2(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n231_), .B1(new_n301_), .B2(new_n300_), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n599_), .A2(KEYINPUT70), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(KEYINPUT70), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n318_), .A2(new_n231_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n600_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(KEYINPUT69), .B(KEYINPUT35), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G232gat), .A2(G233gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  OR3_X1    g407(.A1(new_n603_), .A2(KEYINPUT71), .A3(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G190gat), .B(G218gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G134gat), .B(G162gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  AOI22_X1  g411(.A1(new_n603_), .A2(new_n604_), .B1(KEYINPUT36), .B2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n608_), .B1(new_n603_), .B2(KEYINPUT71), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n609_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n612_), .A2(KEYINPUT36), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n616_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n609_), .A2(new_n613_), .A3(new_n618_), .A4(new_n614_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT37), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n617_), .A2(KEYINPUT37), .A3(new_n619_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n258_), .B(new_n311_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(G231gat), .A2(G233gat), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT72), .Z(new_n627_));
  XNOR2_X1  g426(.A(new_n625_), .B(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(G127gat), .B(G155gat), .Z(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT16), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G183gat), .B(G211gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT17), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT73), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n632_), .A2(new_n635_), .A3(new_n633_), .ZN(new_n636_));
  OR3_X1    g435(.A1(new_n628_), .A2(new_n634_), .A3(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n628_), .A2(new_n636_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n624_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n598_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n643_), .A2(new_n306_), .A3(new_n558_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT38), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n620_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n647_), .B1(new_n595_), .B2(new_n597_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n648_), .A2(new_n639_), .A3(new_n332_), .ZN(new_n649_));
  OAI21_X1  g448(.A(G1gat), .B1(new_n649_), .B2(new_n592_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n644_), .A2(new_n645_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n646_), .A2(new_n650_), .A3(new_n651_), .ZN(G1324gat));
  OAI21_X1  g451(.A(G8gat), .B1(new_n649_), .B2(new_n589_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT39), .ZN(new_n654_));
  INV_X1    g453(.A(new_n589_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n643_), .A2(new_n307_), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n657_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g457(.A(G15gat), .B1(new_n649_), .B2(new_n400_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(KEYINPUT101), .B(KEYINPUT41), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n660_), .ZN(new_n662_));
  OR3_X1    g461(.A1(new_n642_), .A2(G15gat), .A3(new_n400_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n661_), .A2(new_n662_), .A3(new_n663_), .ZN(G1326gat));
  OAI21_X1  g463(.A(G22gat), .B1(new_n649_), .B2(new_n596_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n596_), .A2(G22gat), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n667_), .B1(new_n642_), .B2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT103), .ZN(G1327gat));
  NOR2_X1   g469(.A1(new_n620_), .A2(new_n639_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n598_), .A2(new_n671_), .ZN(new_n672_));
  OR3_X1    g471(.A1(new_n672_), .A2(G29gat), .A3(new_n592_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n333_), .A2(new_n639_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n595_), .A2(new_n597_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n624_), .B(KEYINPUT104), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n675_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n624_), .A2(new_n675_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n679_), .B1(new_n595_), .B2(new_n597_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n674_), .B1(new_n678_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  OAI211_X1 g482(.A(KEYINPUT44), .B(new_n674_), .C1(new_n678_), .C2(new_n680_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n686_), .A2(new_n687_), .A3(new_n558_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(G29gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n687_), .B1(new_n686_), .B2(new_n558_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n673_), .B1(new_n689_), .B2(new_n690_), .ZN(G1328gat));
  INV_X1    g490(.A(KEYINPUT108), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n683_), .A2(new_n655_), .A3(new_n684_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(G36gat), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n589_), .A2(G36gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n598_), .A2(new_n671_), .A3(new_n695_), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT45), .Z(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n694_), .A2(KEYINPUT106), .A3(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT107), .ZN(new_n700_));
  AOI21_X1  g499(.A(KEYINPUT46), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n697_), .B1(new_n693_), .B2(G36gat), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n703_), .B1(new_n700_), .B2(KEYINPUT46), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n702_), .A2(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n692_), .B1(new_n701_), .B2(new_n705_), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n702_), .A2(new_n704_), .ZN(new_n707_));
  AOI21_X1  g506(.A(KEYINPUT107), .B1(new_n702_), .B2(KEYINPUT106), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n707_), .B(KEYINPUT108), .C1(new_n708_), .C2(KEYINPUT46), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n706_), .A2(new_n709_), .ZN(G1329gat));
  NAND3_X1  g509(.A1(new_n686_), .A2(G43gat), .A3(new_n399_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n672_), .A2(new_n400_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n711_), .B1(G43gat), .B2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g513(.A(new_n672_), .ZN(new_n715_));
  AOI21_X1  g514(.A(G50gat), .B1(new_n715_), .B2(new_n474_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n474_), .A2(G50gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n686_), .B2(new_n717_), .ZN(G1331gat));
  NOR2_X1   g517(.A1(new_n330_), .A2(new_n640_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n648_), .A2(new_n297_), .A3(new_n719_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n720_), .A2(new_n235_), .A3(new_n592_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n294_), .A2(KEYINPUT13), .A3(new_n295_), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT13), .B1(new_n294_), .B2(new_n295_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  AOI211_X1 g523(.A(new_n330_), .B(new_n724_), .C1(new_n595_), .C2(new_n597_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n641_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n727_), .A2(KEYINPUT109), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(KEYINPUT109), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n728_), .A2(new_n558_), .A3(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n721_), .B1(new_n730_), .B2(new_n235_), .ZN(G1332gat));
  OAI21_X1  g530(.A(G64gat), .B1(new_n720_), .B2(new_n589_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT48), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n727_), .A2(new_n237_), .A3(new_n655_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1333gat));
  OAI21_X1  g534(.A(G71gat), .B1(new_n720_), .B2(new_n400_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT49), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n727_), .A2(new_n246_), .A3(new_n399_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1334gat));
  OAI21_X1  g538(.A(G78gat), .B1(new_n720_), .B2(new_n596_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT50), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n727_), .A2(new_n244_), .A3(new_n474_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1335gat));
  AND2_X1   g542(.A1(new_n725_), .A2(new_n671_), .ZN(new_n744_));
  AOI21_X1  g543(.A(G85gat), .B1(new_n744_), .B2(new_n558_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT110), .Z(new_n746_));
  OR2_X1    g545(.A1(new_n678_), .A2(new_n680_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n724_), .A2(new_n639_), .A3(new_n330_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n558_), .A2(G85gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n746_), .B1(new_n750_), .B2(new_n751_), .ZN(G1336gat));
  AOI21_X1  g551(.A(G92gat), .B1(new_n744_), .B2(new_n655_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT111), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n750_), .A2(G92gat), .A3(new_n655_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT112), .Z(G1337gat));
  NAND3_X1  g556(.A1(new_n744_), .A2(new_n207_), .A3(new_n399_), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT113), .Z(new_n759_));
  OAI21_X1  g558(.A(G99gat), .B1(new_n749_), .B2(new_n400_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT51), .ZN(G1338gat));
  AOI21_X1  g561(.A(new_n208_), .B1(new_n750_), .B2(new_n474_), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n763_), .A2(KEYINPUT52), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(KEYINPUT52), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n744_), .A2(new_n208_), .A3(new_n474_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT114), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n764_), .A2(new_n765_), .A3(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT53), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n764_), .A2(new_n770_), .A3(new_n765_), .A4(new_n767_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(G1339gat));
  INV_X1    g571(.A(new_n624_), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT115), .B1(new_n724_), .B2(new_n719_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n291_), .A2(new_n719_), .A3(KEYINPUT115), .A4(new_n296_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n773_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT116), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n291_), .A2(new_n296_), .A3(new_n719_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT115), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n775_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(new_n783_), .A3(new_n773_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n778_), .A2(KEYINPUT54), .A3(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT54), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n783_), .B1(new_n782_), .B2(new_n773_), .ZN(new_n787_));
  AOI211_X1 g586(.A(KEYINPUT116), .B(new_n624_), .C1(new_n781_), .C2(new_n775_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n786_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n785_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT118), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n278_), .A2(new_n792_), .A3(new_n281_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT117), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n288_), .A2(KEYINPUT117), .A3(new_n792_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n280_), .A2(KEYINPUT55), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n798_), .B1(new_n264_), .B2(new_n263_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n791_), .B1(new_n797_), .B2(new_n800_), .ZN(new_n801_));
  AOI211_X1 g600(.A(KEYINPUT118), .B(new_n799_), .C1(new_n795_), .C2(new_n796_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n274_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT119), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(KEYINPUT56), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT117), .B1(new_n288_), .B2(new_n792_), .ZN(new_n807_));
  NOR4_X1   g606(.A1(new_n265_), .A2(new_n267_), .A3(new_n794_), .A4(KEYINPUT55), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n800_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT118), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n797_), .A2(new_n791_), .A3(new_n800_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT56), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n812_), .A2(KEYINPUT119), .A3(new_n813_), .A4(new_n274_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n331_), .A2(new_n290_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n805_), .A2(new_n806_), .A3(new_n814_), .A4(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n326_), .B1(new_n316_), .B2(new_n321_), .ZN(new_n817_));
  OR2_X1    g616(.A1(new_n817_), .A2(KEYINPUT120), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(KEYINPUT120), .ZN(new_n819_));
  INV_X1    g618(.A(new_n321_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n313_), .A2(new_n319_), .A3(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n818_), .A2(new_n819_), .A3(new_n821_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n822_), .B(new_n329_), .C1(new_n284_), .C2(new_n290_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n647_), .B1(new_n816_), .B2(new_n823_), .ZN(new_n824_));
  OR2_X1    g623(.A1(new_n824_), .A2(KEYINPUT57), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826_));
  AOI211_X1 g625(.A(new_n826_), .B(new_n647_), .C1(new_n816_), .C2(new_n823_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT58), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n822_), .A2(new_n329_), .A3(new_n295_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(new_n803_), .B2(KEYINPUT56), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n275_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n832_), .A2(new_n813_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n829_), .B1(new_n831_), .B2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n813_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n806_), .A2(new_n835_), .A3(KEYINPUT58), .A4(new_n830_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n834_), .A2(new_n624_), .A3(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n825_), .A2(new_n828_), .A3(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n790_), .B1(new_n838_), .B2(new_n640_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(new_n592_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n400_), .A2(new_n474_), .A3(new_n655_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(G113gat), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(new_n844_), .A3(new_n330_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n839_), .A2(KEYINPUT121), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n846_), .A2(KEYINPUT59), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n842_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n840_), .B(new_n841_), .C1(new_n846_), .C2(KEYINPUT59), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n331_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n845_), .B1(new_n850_), .B2(new_n844_), .ZN(G1340gat));
  INV_X1    g650(.A(G120gat), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n852_), .B1(new_n724_), .B2(KEYINPUT60), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n843_), .B(new_n853_), .C1(KEYINPUT60), .C2(new_n852_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n724_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n852_), .ZN(G1341gat));
  AOI21_X1  g655(.A(G127gat), .B1(new_n843_), .B2(new_n639_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n848_), .A2(new_n849_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n639_), .A2(G127gat), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(KEYINPUT122), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n857_), .B1(new_n858_), .B2(new_n860_), .ZN(G1342gat));
  INV_X1    g660(.A(G134gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n843_), .A2(new_n862_), .A3(new_n647_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n773_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(new_n862_), .ZN(G1343gat));
  NOR3_X1   g664(.A1(new_n399_), .A2(new_n596_), .A3(new_n655_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n840_), .A2(new_n866_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(new_n331_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(new_n436_), .ZN(G1344gat));
  NOR2_X1   g668(.A1(new_n867_), .A2(new_n724_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(new_n437_), .ZN(G1345gat));
  NOR2_X1   g670(.A1(new_n867_), .A2(new_n640_), .ZN(new_n872_));
  XOR2_X1   g671(.A(KEYINPUT61), .B(G155gat), .Z(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1346gat));
  INV_X1    g673(.A(new_n867_), .ZN(new_n875_));
  AOI21_X1  g674(.A(G162gat), .B1(new_n875_), .B2(new_n647_), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n677_), .A2(G162gat), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n876_), .B1(new_n875_), .B2(new_n877_), .ZN(G1347gat));
  AND2_X1   g677(.A1(new_n785_), .A2(new_n789_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n837_), .B1(new_n824_), .B2(KEYINPUT57), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n640_), .B1(new_n880_), .B2(new_n827_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n399_), .A2(new_n592_), .A3(new_n655_), .ZN(new_n883_));
  XOR2_X1   g682(.A(new_n883_), .B(KEYINPUT123), .Z(new_n884_));
  NAND4_X1  g683(.A1(new_n882_), .A2(new_n473_), .A3(new_n469_), .A4(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n331_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n886_), .A2(new_n348_), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n887_), .A2(KEYINPUT62), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n886_), .A2(new_n367_), .A3(new_n369_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(KEYINPUT62), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n888_), .A2(new_n889_), .A3(new_n890_), .ZN(G1348gat));
  NOR2_X1   g690(.A1(new_n885_), .A2(new_n724_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(new_n349_), .ZN(G1349gat));
  NOR2_X1   g692(.A1(new_n885_), .A2(new_n640_), .ZN(new_n894_));
  MUX2_X1   g693(.A(G183gat), .B(new_n345_), .S(new_n894_), .Z(G1350gat));
  OAI21_X1  g694(.A(G190gat), .B1(new_n885_), .B2(new_n773_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n647_), .A2(new_n346_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n885_), .B2(new_n897_), .ZN(G1351gat));
  NOR2_X1   g697(.A1(new_n399_), .A2(new_n596_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n899_), .A2(new_n592_), .A3(new_n655_), .ZN(new_n900_));
  OAI21_X1  g699(.A(KEYINPUT124), .B1(new_n839_), .B2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n902_));
  INV_X1    g701(.A(new_n900_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n882_), .A2(new_n902_), .A3(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n331_), .B1(new_n901_), .B2(new_n904_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(KEYINPUT125), .B(G197gat), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n905_), .B(new_n906_), .ZN(G1352gat));
  AOI21_X1  g706(.A(new_n724_), .B1(new_n901_), .B2(new_n904_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT126), .ZN(new_n909_));
  AND2_X1   g708(.A1(new_n909_), .A2(G204gat), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n909_), .A2(G204gat), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n908_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n912_), .B1(new_n908_), .B2(new_n911_), .ZN(G1353gat));
  AOI21_X1  g712(.A(new_n640_), .B1(new_n901_), .B2(new_n904_), .ZN(new_n914_));
  OR2_X1    g713(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n915_));
  NAND2_X1  g714(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n914_), .A2(new_n915_), .A3(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n917_), .B1(new_n914_), .B2(new_n915_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(G1354gat));
  INV_X1    g718(.A(KEYINPUT127), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n620_), .A2(G218gat), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n902_), .B1(new_n882_), .B2(new_n903_), .ZN(new_n922_));
  AOI211_X1 g721(.A(KEYINPUT124), .B(new_n900_), .C1(new_n879_), .C2(new_n881_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n921_), .B1(new_n922_), .B2(new_n923_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n773_), .B1(new_n901_), .B2(new_n904_), .ZN(new_n925_));
  INV_X1    g724(.A(G218gat), .ZN(new_n926_));
  OAI211_X1 g725(.A(new_n920_), .B(new_n924_), .C1(new_n925_), .C2(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n624_), .B1(new_n922_), .B2(new_n923_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(G218gat), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n920_), .B1(new_n930_), .B2(new_n924_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n928_), .A2(new_n931_), .ZN(G1355gat));
endmodule


