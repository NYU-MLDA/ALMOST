//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 1 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n855_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_;
  XOR2_X1   g000(.A(G1gat), .B(G29gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT100), .B(KEYINPUT0), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT92), .ZN(new_n208_));
  OR2_X1    g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT90), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT1), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT91), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n209_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT90), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n210_), .B(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT1), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n218_), .A2(KEYINPUT91), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n208_), .B1(new_n214_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(KEYINPUT91), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n212_), .A2(new_n213_), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n221_), .A2(new_n222_), .A3(KEYINPUT92), .A4(new_n209_), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n220_), .B(new_n223_), .C1(KEYINPUT1), .C2(new_n211_), .ZN(new_n224_));
  XOR2_X1   g023(.A(G141gat), .B(G148gat), .Z(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  OR3_X1    g025(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G141gat), .A2(G148gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT2), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n227_), .A2(new_n230_), .A3(new_n231_), .A4(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n233_), .A2(new_n211_), .A3(new_n209_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n226_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G127gat), .B(G134gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G113gat), .B(G120gat), .ZN(new_n237_));
  XOR2_X1   g036(.A(new_n236_), .B(new_n237_), .Z(new_n238_));
  NAND2_X1  g037(.A1(new_n235_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n234_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n240_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n238_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n239_), .A2(KEYINPUT4), .A3(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G225gat), .A2(G233gat), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n242_), .B1(new_n226_), .B2(new_n234_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT4), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n245_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n244_), .A2(KEYINPUT99), .A3(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n239_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(KEYINPUT99), .B1(new_n244_), .B2(new_n248_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n207_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT99), .ZN(new_n254_));
  AOI211_X1 g053(.A(new_n238_), .B(new_n240_), .C1(new_n224_), .C2(new_n225_), .ZN(new_n255_));
  NOR3_X1   g054(.A1(new_n246_), .A2(new_n255_), .A3(new_n247_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n235_), .A2(new_n247_), .A3(new_n238_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n245_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n254_), .B1(new_n256_), .B2(new_n259_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n260_), .A2(new_n206_), .A3(new_n250_), .A4(new_n249_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n253_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT25), .B(G183gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT95), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT26), .B(G190gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G183gat), .A2(G190gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT87), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n267_), .B1(new_n269_), .B2(KEYINPUT23), .ZN(new_n270_));
  NOR3_X1   g069(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G169gat), .A2(G176gat), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n271_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n266_), .A2(new_n270_), .A3(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT96), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT96), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n266_), .A2(new_n278_), .A3(new_n270_), .A4(new_n275_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(KEYINPUT22), .B(G169gat), .Z(new_n281_));
  OAI21_X1  g080(.A(new_n274_), .B1(new_n281_), .B2(G176gat), .ZN(new_n282_));
  MUX2_X1   g081(.A(new_n269_), .B(new_n268_), .S(KEYINPUT23), .Z(new_n283_));
  INV_X1    g082(.A(G183gat), .ZN(new_n284_));
  INV_X1    g083(.A(G190gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n282_), .B1(new_n283_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n280_), .A2(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(G197gat), .B(G204gat), .Z(new_n290_));
  OR2_X1    g089(.A1(new_n290_), .A2(KEYINPUT21), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(KEYINPUT21), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G211gat), .B(G218gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n291_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n292_), .A2(new_n293_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT86), .B(G183gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n285_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n270_), .A2(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT88), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(G169gat), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n301_), .A2(G169gat), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n299_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT25), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n284_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n306_), .B1(new_n297_), .B2(new_n305_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n265_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n283_), .A2(new_n275_), .A3(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n304_), .A2(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT20), .B1(new_n310_), .B2(new_n296_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT94), .ZN(new_n312_));
  AOI22_X1  g111(.A1(new_n289_), .A2(new_n296_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G226gat), .A2(G233gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT19), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n311_), .A2(new_n312_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n313_), .A2(new_n316_), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT20), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n320_), .B1(new_n310_), .B2(new_n296_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n296_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n288_), .A2(new_n322_), .A3(new_n276_), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n319_), .B1(new_n316_), .B2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G8gat), .B(G36gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT18), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G64gat), .B(G92gat), .ZN(new_n328_));
  XOR2_X1   g127(.A(new_n327_), .B(new_n328_), .Z(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT32), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n325_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n311_), .A2(new_n312_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n287_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n333_), .B1(new_n322_), .B2(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n315_), .B1(new_n335_), .B2(new_n317_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n322_), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n337_), .A2(KEYINPUT97), .A3(new_n316_), .A4(new_n321_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT97), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n321_), .A2(new_n316_), .ZN(new_n340_));
  AOI211_X1 g139(.A(new_n296_), .B(new_n287_), .C1(new_n277_), .C2(new_n279_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n339_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n336_), .A2(new_n338_), .A3(new_n342_), .A4(new_n330_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n332_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n262_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT101), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT29), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n296_), .B1(new_n241_), .B2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n350_), .A2(G228gat), .A3(G233gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G228gat), .A2(G233gat), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n352_), .B(new_n296_), .C1(new_n241_), .C2(new_n349_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G78gat), .B(G106gat), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT93), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n354_), .A2(new_n355_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n241_), .A2(new_n349_), .ZN(new_n360_));
  XOR2_X1   g159(.A(G22gat), .B(G50gat), .Z(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT28), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n360_), .B(new_n362_), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n357_), .A2(new_n358_), .A3(new_n359_), .A4(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n359_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n358_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n363_), .ZN(new_n367_));
  OAI22_X1  g166(.A1(new_n365_), .A2(new_n356_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n364_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n329_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n316_), .B1(new_n313_), .B2(new_n318_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n342_), .A2(new_n338_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n370_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n336_), .A2(new_n329_), .A3(new_n338_), .A4(new_n342_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT98), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT98), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n373_), .A2(new_n374_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n249_), .A2(new_n250_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n380_), .A2(KEYINPUT33), .A3(new_n206_), .A4(new_n260_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT33), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n261_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n244_), .A2(new_n245_), .A3(new_n257_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n239_), .A2(new_n243_), .A3(new_n258_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n384_), .A2(new_n207_), .A3(new_n385_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n379_), .A2(new_n381_), .A3(new_n383_), .A4(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n262_), .A2(KEYINPUT101), .A3(new_n345_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n348_), .A2(new_n369_), .A3(new_n387_), .A4(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G71gat), .B(G99gat), .ZN(new_n390_));
  INV_X1    g189(.A(G43gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n310_), .B(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G227gat), .A2(G233gat), .ZN(new_n394_));
  INV_X1    g193(.A(G15gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT30), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT31), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n393_), .B(new_n398_), .ZN(new_n399_));
  XOR2_X1   g198(.A(new_n399_), .B(KEYINPUT89), .Z(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(new_n238_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT102), .B(KEYINPUT27), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n375_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n325_), .A2(new_n370_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n404_), .A2(KEYINPUT27), .A3(new_n374_), .ZN(new_n405_));
  AND4_X1   g204(.A1(new_n253_), .A2(new_n403_), .A3(new_n261_), .A4(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n401_), .B1(new_n406_), .B2(new_n369_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n389_), .A2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n400_), .B(new_n242_), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n406_), .A2(new_n369_), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n409_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT81), .B(G15gat), .ZN(new_n414_));
  INV_X1    g213(.A(G22gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(G1gat), .ZN(new_n417_));
  INV_X1    g216(.A(G8gat), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT14), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n416_), .A2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G1gat), .B(G8gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT82), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n420_), .B(new_n422_), .ZN(new_n423_));
  XOR2_X1   g222(.A(G29gat), .B(G36gat), .Z(new_n424_));
  XOR2_X1   g223(.A(G43gat), .B(G50gat), .Z(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT84), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n423_), .B(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT85), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(G229gat), .A3(G233gat), .ZN(new_n431_));
  INV_X1    g230(.A(new_n423_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n426_), .B(KEYINPUT15), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G229gat), .A2(G233gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n423_), .A2(new_n428_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n434_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n431_), .A2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G113gat), .B(G141gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G169gat), .B(G197gat), .ZN(new_n440_));
  XOR2_X1   g239(.A(new_n439_), .B(new_n440_), .Z(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n438_), .A2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n431_), .A2(new_n437_), .A3(new_n441_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n413_), .A2(new_n445_), .ZN(new_n446_));
  XOR2_X1   g245(.A(KEYINPUT64), .B(G85gat), .Z(new_n447_));
  INV_X1    g246(.A(G92gat), .ZN(new_n448_));
  OR3_X1    g247(.A1(new_n447_), .A2(KEYINPUT9), .A3(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G85gat), .B(G92gat), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT9), .ZN(new_n452_));
  XOR2_X1   g251(.A(KEYINPUT10), .B(G99gat), .Z(new_n453_));
  INV_X1    g252(.A(G106gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(G99gat), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT6), .B1(new_n456_), .B2(new_n454_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT6), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n458_), .A2(G99gat), .A3(G106gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n449_), .A2(new_n452_), .A3(new_n455_), .A4(new_n460_), .ZN(new_n461_));
  XOR2_X1   g260(.A(new_n450_), .B(KEYINPUT66), .Z(new_n462_));
  INV_X1    g261(.A(KEYINPUT8), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n456_), .A2(new_n454_), .A3(KEYINPUT65), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT7), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT65), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n466_), .A2(G99gat), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT7), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n467_), .A2(new_n468_), .A3(new_n454_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n460_), .A2(new_n465_), .A3(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n462_), .A2(new_n463_), .A3(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n468_), .B1(new_n467_), .B2(new_n454_), .ZN(new_n472_));
  NOR4_X1   g271(.A1(new_n466_), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT69), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT69), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n469_), .A2(new_n465_), .A3(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n460_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n477_), .A2(new_n457_), .A3(new_n459_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n474_), .A2(new_n476_), .A3(new_n479_), .A4(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n463_), .B1(new_n481_), .B2(new_n462_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT70), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n471_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  AOI211_X1 g283(.A(KEYINPUT70), .B(new_n463_), .C1(new_n481_), .C2(new_n462_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n461_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT72), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  OAI211_X1 g287(.A(KEYINPUT72), .B(new_n461_), .C1(new_n484_), .C2(new_n485_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(new_n433_), .A3(new_n489_), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n426_), .B(new_n461_), .C1(new_n484_), .C2(new_n485_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT76), .B(KEYINPUT34), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G232gat), .A2(G233gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT35), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n491_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n490_), .A2(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n495_), .A2(new_n496_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(G190gat), .B(G218gat), .Z(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT77), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G134gat), .B(G162gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n505_), .A2(KEYINPUT36), .ZN(new_n506_));
  INV_X1    g305(.A(new_n500_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n490_), .A2(new_n507_), .A3(new_n498_), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n501_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n505_), .B(KEYINPUT36), .Z(new_n510_));
  XOR2_X1   g309(.A(new_n510_), .B(KEYINPUT78), .Z(new_n511_));
  AOI21_X1  g310(.A(new_n511_), .B1(new_n501_), .B2(new_n508_), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT37), .B1(new_n509_), .B2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT79), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT80), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n490_), .A2(new_n507_), .A3(new_n498_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n507_), .B1(new_n490_), .B2(new_n498_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n515_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n501_), .A2(KEYINPUT80), .A3(new_n508_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n511_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n501_), .A2(new_n506_), .A3(new_n508_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n523_), .A2(KEYINPUT37), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n514_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G127gat), .B(G155gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT16), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G183gat), .B(G211gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(KEYINPUT83), .B1(new_n529_), .B2(KEYINPUT17), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G231gat), .A2(G233gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G57gat), .B(G64gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G71gat), .B(G78gat), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n533_), .A2(new_n534_), .A3(KEYINPUT11), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n533_), .A2(KEYINPUT11), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n536_), .A2(new_n534_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n533_), .A2(KEYINPUT11), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n535_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n532_), .B(new_n539_), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n540_), .A2(new_n423_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n529_), .A2(KEYINPUT17), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n542_), .B1(new_n540_), .B2(new_n423_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT75), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n545_), .A2(KEYINPUT13), .ZN(new_n546_));
  INV_X1    g345(.A(new_n539_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT12), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n488_), .A2(new_n489_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT73), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n486_), .A2(new_n547_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT12), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n488_), .A2(KEYINPUT73), .A3(new_n489_), .A4(new_n549_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n461_), .B(new_n539_), .C1(new_n484_), .C2(new_n485_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  AND2_X1   g357(.A1(G230gat), .A2(G233gat), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n552_), .A2(new_n555_), .A3(new_n556_), .A4(new_n560_), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n557_), .A2(KEYINPUT71), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n557_), .A2(KEYINPUT71), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n562_), .A2(new_n553_), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(new_n559_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n561_), .A2(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(G120gat), .B(G148gat), .Z(new_n567_));
  XNOR2_X1  g366(.A(G176gat), .B(G204gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT74), .B(KEYINPUT5), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n566_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n566_), .A2(new_n571_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n546_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT75), .B(KEYINPUT13), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n572_), .A2(new_n573_), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n525_), .A2(new_n544_), .A3(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n446_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n262_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n582_), .A2(KEYINPUT103), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(KEYINPUT103), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n581_), .A2(new_n417_), .A3(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT38), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT105), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n523_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n521_), .A2(KEYINPUT105), .A3(new_n522_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n387_), .A2(new_n369_), .ZN(new_n593_));
  AOI21_X1  g392(.A(KEYINPUT101), .B1(new_n262_), .B2(new_n345_), .ZN(new_n594_));
  AOI211_X1 g393(.A(new_n347_), .B(new_n344_), .C1(new_n253_), .C2(new_n261_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n407_), .B1(new_n593_), .B2(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n592_), .B1(new_n597_), .B2(new_n411_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n578_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n599_), .A2(new_n574_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n445_), .ZN(new_n601_));
  OAI21_X1  g400(.A(KEYINPUT104), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT104), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n579_), .A2(new_n603_), .A3(new_n445_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n602_), .A2(new_n604_), .A3(new_n544_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n598_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(G1gat), .B1(new_n607_), .B2(new_n582_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n587_), .A2(new_n608_), .ZN(G1324gat));
  XNOR2_X1  g408(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n411_), .B1(new_n389_), .B2(new_n408_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n611_), .A2(new_n591_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n603_), .B1(new_n579_), .B2(new_n445_), .ZN(new_n613_));
  AOI211_X1 g412(.A(KEYINPUT104), .B(new_n601_), .C1(new_n575_), .C2(new_n578_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n403_), .A2(new_n405_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n612_), .A2(new_n615_), .A3(new_n617_), .A4(new_n544_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT106), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n606_), .A2(KEYINPUT106), .A3(new_n617_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n620_), .A2(new_n621_), .A3(G8gat), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT107), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n623_), .A2(KEYINPUT39), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n616_), .A2(G8gat), .ZN(new_n625_));
  AOI22_X1  g424(.A1(new_n622_), .A2(new_n624_), .B1(new_n581_), .B2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT107), .B(KEYINPUT39), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n620_), .A2(new_n621_), .A3(G8gat), .A4(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n610_), .B1(new_n626_), .B2(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(G8gat), .B1(new_n618_), .B2(new_n619_), .ZN(new_n630_));
  AOI21_X1  g429(.A(KEYINPUT106), .B1(new_n606_), .B2(new_n617_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n624_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n581_), .A2(new_n625_), .ZN(new_n633_));
  AND4_X1   g432(.A1(new_n628_), .A2(new_n632_), .A3(new_n633_), .A4(new_n610_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n629_), .A2(new_n634_), .ZN(G1325gat));
  NAND2_X1  g434(.A1(new_n606_), .A2(new_n410_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(G15gat), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(KEYINPUT41), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT41), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n636_), .A2(new_n639_), .A3(G15gat), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT109), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n581_), .A2(new_n395_), .A3(new_n410_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT110), .Z(new_n645_));
  NAND3_X1  g444(.A1(new_n638_), .A2(KEYINPUT109), .A3(new_n640_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n643_), .A2(new_n645_), .A3(new_n646_), .ZN(G1326gat));
  INV_X1    g446(.A(new_n369_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n415_), .B1(new_n606_), .B2(new_n648_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT42), .Z(new_n650_));
  NAND3_X1  g449(.A1(new_n581_), .A2(new_n415_), .A3(new_n648_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1327gat));
  INV_X1    g451(.A(KEYINPUT43), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n653_), .B1(new_n611_), .B2(new_n525_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n525_), .ZN(new_n655_));
  OAI211_X1 g454(.A(KEYINPUT43), .B(new_n655_), .C1(new_n597_), .C2(new_n411_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n544_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n654_), .A2(new_n656_), .A3(new_n657_), .A4(new_n615_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT44), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n655_), .B1(new_n597_), .B2(new_n411_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n544_), .B1(new_n661_), .B2(new_n653_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n662_), .A2(KEYINPUT44), .A3(new_n615_), .A4(new_n656_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n660_), .A2(new_n663_), .A3(G29gat), .A4(new_n585_), .ZN(new_n664_));
  INV_X1    g463(.A(G29gat), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT111), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n591_), .A2(new_n657_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n667_), .A2(new_n600_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n666_), .B1(new_n446_), .B2(new_n669_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n413_), .A2(KEYINPUT111), .A3(new_n445_), .A4(new_n668_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n665_), .B1(new_n672_), .B2(new_n582_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n664_), .A2(new_n673_), .ZN(G1328gat));
  NAND3_X1  g473(.A1(new_n660_), .A2(new_n663_), .A3(new_n617_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(G36gat), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n616_), .A2(G36gat), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n670_), .A2(new_n671_), .A3(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT45), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT45), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n670_), .A2(new_n680_), .A3(new_n671_), .A4(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n676_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT46), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n676_), .A2(new_n682_), .A3(KEYINPUT46), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1329gat));
  NAND4_X1  g486(.A1(new_n660_), .A2(new_n663_), .A3(G43gat), .A4(new_n410_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n391_), .B1(new_n672_), .B2(new_n401_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g490(.A1(new_n660_), .A2(new_n663_), .A3(G50gat), .A4(new_n648_), .ZN(new_n692_));
  INV_X1    g491(.A(G50gat), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n693_), .B1(new_n672_), .B2(new_n369_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n692_), .A2(new_n694_), .ZN(G1331gat));
  NOR2_X1   g494(.A1(new_n611_), .A2(new_n445_), .ZN(new_n696_));
  AND4_X1   g495(.A1(new_n544_), .A2(new_n696_), .A3(new_n600_), .A4(new_n525_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(new_n585_), .ZN(new_n698_));
  INV_X1    g497(.A(G57gat), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n700_), .A2(KEYINPUT112), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(KEYINPUT112), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n612_), .A2(new_n544_), .A3(new_n601_), .A4(new_n600_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT113), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n582_), .A2(new_n699_), .ZN(new_n705_));
  AOI22_X1  g504(.A1(new_n701_), .A2(new_n702_), .B1(new_n704_), .B2(new_n705_), .ZN(G1332gat));
  INV_X1    g505(.A(G64gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n697_), .A2(new_n707_), .A3(new_n617_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT48), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n704_), .A2(new_n617_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n710_), .B2(G64gat), .ZN(new_n711_));
  AOI211_X1 g510(.A(KEYINPUT48), .B(new_n707_), .C1(new_n704_), .C2(new_n617_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n708_), .B1(new_n711_), .B2(new_n712_), .ZN(G1333gat));
  INV_X1    g512(.A(G71gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n697_), .A2(new_n714_), .A3(new_n410_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT49), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n704_), .A2(new_n410_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n717_), .B2(G71gat), .ZN(new_n718_));
  AOI211_X1 g517(.A(KEYINPUT49), .B(new_n714_), .C1(new_n704_), .C2(new_n410_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n715_), .B1(new_n718_), .B2(new_n719_), .ZN(G1334gat));
  INV_X1    g519(.A(G78gat), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n697_), .A2(new_n721_), .A3(new_n648_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT50), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n704_), .A2(new_n648_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n723_), .B1(new_n724_), .B2(G78gat), .ZN(new_n725_));
  AOI211_X1 g524(.A(KEYINPUT50), .B(new_n721_), .C1(new_n704_), .C2(new_n648_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n722_), .B1(new_n725_), .B2(new_n726_), .ZN(G1335gat));
  NOR2_X1   g526(.A1(new_n667_), .A2(new_n579_), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n696_), .A2(KEYINPUT114), .A3(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(KEYINPUT114), .B1(new_n696_), .B2(new_n728_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(G85gat), .B1(new_n732_), .B2(new_n585_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n579_), .A2(new_n445_), .ZN(new_n734_));
  NAND4_X1  g533(.A1(new_n654_), .A2(new_n656_), .A3(new_n657_), .A4(new_n734_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n735_), .A2(new_n582_), .A3(new_n447_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n733_), .A2(new_n736_), .ZN(G1336gat));
  OAI21_X1  g536(.A(G92gat), .B1(new_n735_), .B2(new_n616_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n617_), .A2(new_n448_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n731_), .B2(new_n739_), .ZN(G1337gat));
  OAI21_X1  g539(.A(G99gat), .B1(new_n735_), .B2(new_n401_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n410_), .A2(new_n453_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n741_), .B1(new_n731_), .B2(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n743_), .B(new_n744_), .Z(G1338gat));
  OAI211_X1 g544(.A(new_n454_), .B(new_n648_), .C1(new_n729_), .C2(new_n730_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT52), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n747_), .B(G106gat), .C1(new_n735_), .C2(new_n369_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n662_), .A2(new_n648_), .A3(new_n656_), .A4(new_n734_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n747_), .B1(new_n750_), .B2(G106gat), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n746_), .B1(new_n749_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT53), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT53), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n746_), .B(new_n754_), .C1(new_n749_), .C2(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1339gat));
  XNOR2_X1  g555(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n583_), .A2(new_n584_), .A3(new_n617_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n648_), .A2(new_n401_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n757_), .B1(new_n760_), .B2(KEYINPUT119), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n572_), .A2(new_n445_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n552_), .A2(new_n555_), .A3(new_n556_), .A4(new_n557_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n559_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n561_), .A2(new_n765_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n556_), .A2(new_n555_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n767_), .A2(KEYINPUT55), .A3(new_n552_), .A4(new_n560_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n764_), .A2(new_n766_), .A3(new_n768_), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n769_), .A2(KEYINPUT56), .A3(new_n571_), .ZN(new_n770_));
  AOI21_X1  g569(.A(KEYINPUT56), .B1(new_n769_), .B2(new_n571_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n762_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n572_), .A2(new_n573_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n430_), .A2(new_n435_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n435_), .B1(new_n423_), .B2(new_n428_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n441_), .B1(new_n434_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n444_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n773_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n772_), .A2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT57), .B1(new_n780_), .B2(new_n592_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT57), .ZN(new_n782_));
  AOI211_X1 g581(.A(new_n782_), .B(new_n591_), .C1(new_n772_), .C2(new_n779_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n572_), .A2(new_n778_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n769_), .A2(new_n571_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT56), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n769_), .A2(KEYINPUT56), .A3(new_n571_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n785_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT116), .ZN(new_n791_));
  OAI21_X1  g590(.A(KEYINPUT58), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n572_), .A2(new_n778_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n793_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT58), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n794_), .A2(KEYINPUT116), .A3(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n792_), .A2(new_n655_), .A3(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n544_), .B1(new_n784_), .B2(new_n797_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n525_), .A2(new_n579_), .A3(new_n544_), .A4(new_n601_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n799_), .B(new_n800_), .ZN(new_n801_));
  OAI221_X1 g600(.A(new_n761_), .B1(KEYINPUT119), .B2(new_n760_), .C1(new_n798_), .C2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT117), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n797_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n794_), .A2(KEYINPUT116), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n525_), .B1(new_n805_), .B2(KEYINPUT58), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(KEYINPUT117), .A3(new_n796_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n804_), .A2(new_n784_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n657_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n801_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n760_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT59), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n445_), .B(new_n802_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(G113gat), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n809_), .A2(new_n810_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n760_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  OR3_X1    g616(.A1(new_n817_), .A2(G113gat), .A3(new_n601_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n814_), .A2(new_n818_), .ZN(G1340gat));
  OAI211_X1 g618(.A(new_n600_), .B(new_n802_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(G120gat), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n579_), .A2(KEYINPUT60), .ZN(new_n822_));
  MUX2_X1   g621(.A(new_n822_), .B(KEYINPUT60), .S(G120gat), .Z(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT117), .B1(new_n806_), .B2(new_n796_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n572_), .A2(new_n445_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n825_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n779_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n592_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n782_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n780_), .A2(KEYINPUT57), .A3(new_n592_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n824_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n544_), .B1(new_n832_), .B2(new_n807_), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n816_), .B(new_n823_), .C1(new_n833_), .C2(new_n801_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(KEYINPUT120), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT120), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n811_), .A2(new_n836_), .A3(new_n823_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n821_), .A2(new_n838_), .ZN(G1341gat));
  INV_X1    g638(.A(G127gat), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n817_), .B2(new_n657_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n544_), .A2(G127gat), .ZN(new_n842_));
  XOR2_X1   g641(.A(new_n842_), .B(KEYINPUT121), .Z(new_n843_));
  OAI211_X1 g642(.A(new_n802_), .B(new_n843_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n841_), .A2(new_n844_), .ZN(G1342gat));
  OAI211_X1 g644(.A(new_n655_), .B(new_n802_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(G134gat), .ZN(new_n847_));
  OR3_X1    g646(.A1(new_n817_), .A2(G134gat), .A3(new_n592_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(G1343gat));
  NOR2_X1   g648(.A1(new_n410_), .A2(new_n369_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n758_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n815_), .A2(new_n445_), .A3(new_n852_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g653(.A1(new_n815_), .A2(new_n600_), .A3(new_n852_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(G148gat), .ZN(G1345gat));
  AOI21_X1  g655(.A(new_n801_), .B1(new_n808_), .B2(new_n657_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n857_), .A2(new_n657_), .A3(new_n851_), .ZN(new_n858_));
  XOR2_X1   g657(.A(KEYINPUT61), .B(G155gat), .Z(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(G1346gat));
  INV_X1    g659(.A(G162gat), .ZN(new_n861_));
  NOR4_X1   g660(.A1(new_n857_), .A2(new_n861_), .A3(new_n525_), .A4(new_n851_), .ZN(new_n862_));
  NOR3_X1   g661(.A1(new_n857_), .A2(new_n592_), .A3(new_n851_), .ZN(new_n863_));
  OAI21_X1  g662(.A(KEYINPUT122), .B1(new_n863_), .B2(G162gat), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n815_), .A2(new_n591_), .A3(new_n852_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n866_), .A3(new_n861_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n862_), .B1(new_n864_), .B2(new_n867_), .ZN(G1347gat));
  NOR3_X1   g667(.A1(new_n585_), .A2(new_n616_), .A3(new_n401_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n369_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n871_), .B1(new_n798_), .B2(new_n801_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(KEYINPUT124), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT124), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n874_), .B(new_n871_), .C1(new_n798_), .C2(new_n801_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n601_), .A2(new_n281_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  XOR2_X1   g677(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n879_));
  OAI211_X1 g678(.A(new_n445_), .B(new_n871_), .C1(new_n798_), .C2(new_n801_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(G169gat), .ZN(new_n881_));
  AND3_X1   g680(.A1(new_n880_), .A2(G169gat), .A3(new_n879_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n878_), .B1(new_n881_), .B2(new_n882_), .ZN(G1348gat));
  AOI21_X1  g682(.A(G176gat), .B1(new_n876_), .B2(new_n600_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n869_), .A2(G176gat), .A3(new_n600_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n857_), .A2(new_n648_), .A3(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n884_), .A2(new_n886_), .ZN(G1349gat));
  NOR2_X1   g686(.A1(new_n657_), .A2(new_n264_), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n815_), .A2(new_n369_), .A3(new_n544_), .A4(new_n869_), .ZN(new_n889_));
  AOI22_X1  g688(.A1(new_n876_), .A2(new_n888_), .B1(new_n889_), .B2(new_n297_), .ZN(G1350gat));
  NAND2_X1  g689(.A1(new_n591_), .A2(new_n265_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(KEYINPUT125), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n876_), .A2(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n525_), .B1(new_n873_), .B2(new_n875_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n285_), .B2(new_n894_), .ZN(G1351gat));
  NOR4_X1   g694(.A1(new_n410_), .A2(new_n369_), .A3(new_n616_), .A4(new_n262_), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n815_), .A2(new_n896_), .ZN(new_n897_));
  AOI21_X1  g696(.A(G197gat), .B1(new_n897_), .B2(new_n445_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n815_), .A2(new_n896_), .ZN(new_n899_));
  INV_X1    g698(.A(G197gat), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n899_), .A2(new_n900_), .A3(new_n601_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n898_), .A2(new_n901_), .ZN(G1352gat));
  NAND3_X1  g701(.A1(new_n815_), .A2(new_n600_), .A3(new_n896_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g703(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(KEYINPUT126), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n657_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n897_), .B2(new_n907_), .ZN(new_n908_));
  AND4_X1   g707(.A1(new_n815_), .A2(new_n896_), .A3(new_n906_), .A4(new_n907_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n908_), .A2(new_n909_), .ZN(G1354gat));
  OR3_X1    g709(.A1(new_n899_), .A2(G218gat), .A3(new_n592_), .ZN(new_n911_));
  OAI21_X1  g710(.A(G218gat), .B1(new_n899_), .B2(new_n525_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1355gat));
endmodule


