//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 1 1 0 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 1 0 0 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n766_, new_n767_, new_n768_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n901_, new_n903_, new_n904_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n946_, new_n947_, new_n949_,
    new_n950_, new_n951_, new_n953_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n960_, new_n961_, new_n962_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT84), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G113gat), .B(G120gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT31), .ZN(new_n207_));
  XOR2_X1   g006(.A(G15gat), .B(G43gat), .Z(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT24), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n210_), .B1(G169gat), .B2(G176gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT81), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n211_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT23), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n219_), .A2(G183gat), .A3(G190gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n216_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT25), .B(G183gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT26), .B(G190gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT80), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n214_), .A2(new_n215_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(new_n210_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n223_), .A2(new_n224_), .A3(KEYINPUT80), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n222_), .A2(new_n227_), .A3(new_n229_), .A4(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(G183gat), .A2(G190gat), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n232_), .B1(new_n218_), .B2(new_n220_), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n233_), .A2(KEYINPUT82), .ZN(new_n234_));
  OR3_X1    g033(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n233_), .A2(KEYINPUT82), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n234_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n231_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G227gat), .A2(G233gat), .ZN(new_n241_));
  XOR2_X1   g040(.A(new_n241_), .B(KEYINPUT83), .Z(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT30), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n240_), .B(new_n243_), .ZN(new_n244_));
  XOR2_X1   g043(.A(G71gat), .B(G99gat), .Z(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n209_), .B(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G228gat), .A2(G233gat), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT29), .ZN(new_n251_));
  XOR2_X1   g050(.A(G141gat), .B(G148gat), .Z(new_n252_));
  INV_X1    g051(.A(G155gat), .ZN(new_n253_));
  INV_X1    g052(.A(G162gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n253_), .A2(new_n254_), .A3(KEYINPUT85), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT85), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n256_), .B1(G155gat), .B2(G162gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT86), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G155gat), .A2(G162gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT1), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n258_), .A2(new_n259_), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n260_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT1), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  AOI22_X1  g065(.A1(new_n255_), .A2(new_n257_), .B1(KEYINPUT1), .B2(new_n260_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n267_), .A2(new_n259_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n252_), .B1(new_n266_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n258_), .A2(new_n260_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NOR3_X1   g071(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n273_));
  AOI21_X1  g072(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n274_));
  NOR3_X1   g073(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT87), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n270_), .B1(new_n275_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n251_), .B1(new_n269_), .B2(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(G197gat), .B(G204gat), .Z(new_n281_));
  XOR2_X1   g080(.A(G211gat), .B(G218gat), .Z(new_n282_));
  NAND3_X1  g081(.A1(new_n281_), .A2(new_n282_), .A3(KEYINPUT21), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT90), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT90), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n281_), .A2(new_n282_), .A3(new_n285_), .A4(KEYINPUT21), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G197gat), .B(G204gat), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT89), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n282_), .B1(new_n289_), .B2(KEYINPUT21), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT21), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n287_), .A2(new_n288_), .A3(new_n291_), .ZN(new_n292_));
  AOI22_X1  g091(.A1(new_n284_), .A2(new_n286_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n250_), .B1(new_n280_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n284_), .A2(new_n286_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n290_), .A2(new_n292_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n258_), .A2(new_n261_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT86), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n299_), .A2(new_n262_), .A3(new_n265_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n278_), .B1(new_n300_), .B2(new_n252_), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n249_), .B(new_n297_), .C1(new_n301_), .C2(new_n251_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G78gat), .B(G106gat), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n303_), .B(KEYINPUT91), .Z(new_n304_));
  NAND3_X1  g103(.A1(new_n294_), .A2(new_n302_), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT93), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(G22gat), .B(G50gat), .Z(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n269_), .A2(new_n251_), .A3(new_n279_), .ZN(new_n310_));
  XOR2_X1   g109(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n311_));
  NOR2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n311_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n313_), .B1(new_n301_), .B2(new_n251_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n309_), .B1(new_n312_), .B2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n310_), .A2(new_n311_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n301_), .A2(new_n251_), .A3(new_n313_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n316_), .A2(new_n317_), .A3(new_n308_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n315_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n294_), .A2(new_n302_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n304_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n294_), .A2(new_n302_), .A3(KEYINPUT93), .A4(new_n304_), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n307_), .A2(new_n319_), .A3(new_n322_), .A4(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT94), .ZN(new_n325_));
  AOI22_X1  g124(.A1(new_n318_), .A2(new_n315_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT94), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n326_), .A2(new_n327_), .A3(new_n323_), .A4(new_n307_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n322_), .A2(new_n305_), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n315_), .A2(new_n318_), .ZN(new_n330_));
  AND3_X1   g129(.A1(new_n329_), .A2(KEYINPUT92), .A3(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(KEYINPUT92), .B1(new_n329_), .B2(new_n330_), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n325_), .B(new_n328_), .C1(new_n331_), .C2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT95), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n329_), .A2(new_n330_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT92), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n329_), .A2(new_n330_), .A3(KEYINPUT92), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n340_), .A2(KEYINPUT95), .A3(new_n328_), .A4(new_n325_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n335_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n204_), .A2(new_n205_), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n204_), .A2(new_n205_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n301_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n269_), .A2(new_n279_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(new_n206_), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G225gat), .A2(G233gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n345_), .A2(new_n347_), .A3(KEYINPUT4), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT4), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n346_), .A2(new_n206_), .A3(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n349_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n351_), .A2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G1gat), .B(G29gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(G85gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT0), .B(G57gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n358_), .B(new_n359_), .Z(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n356_), .A2(new_n361_), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n351_), .A2(new_n355_), .A3(new_n360_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT27), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G8gat), .B(G36gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT18), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G64gat), .B(G92gat), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n367_), .B(new_n368_), .Z(new_n369_));
  NAND2_X1  g168(.A1(G226gat), .A2(G233gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT19), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n293_), .A2(new_n231_), .A3(new_n239_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT20), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n212_), .A2(new_n210_), .ZN(new_n374_));
  AND4_X1   g173(.A1(new_n216_), .A2(new_n225_), .A3(new_n221_), .A4(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n233_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT97), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n376_), .A2(new_n237_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n235_), .A2(new_n236_), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT97), .B1(new_n233_), .B2(new_n379_), .ZN(new_n380_));
  AOI22_X1  g179(.A1(new_n375_), .A2(KEYINPUT96), .B1(new_n378_), .B2(new_n380_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n225_), .A2(new_n216_), .A3(new_n221_), .A4(new_n374_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT96), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n293_), .B1(new_n381_), .B2(new_n384_), .ZN(new_n385_));
  OAI211_X1 g184(.A(KEYINPUT98), .B(new_n371_), .C1(new_n373_), .C2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n378_), .A2(new_n380_), .ZN(new_n388_));
  AOI22_X1  g187(.A1(new_n223_), .A2(new_n224_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n389_), .A2(KEYINPUT96), .A3(new_n216_), .A4(new_n221_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n388_), .A2(new_n384_), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n297_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n392_), .A2(KEYINPUT20), .A3(new_n372_), .ZN(new_n393_));
  AOI21_X1  g192(.A(KEYINPUT98), .B1(new_n393_), .B2(new_n371_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n387_), .A2(new_n394_), .ZN(new_n395_));
  OR3_X1    g194(.A1(new_n391_), .A2(new_n297_), .A3(KEYINPUT99), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT99), .B1(new_n391_), .B2(new_n297_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n371_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT20), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n399_), .B1(new_n240_), .B2(new_n297_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n396_), .A2(new_n397_), .A3(new_n398_), .A4(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n369_), .B1(new_n395_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT98), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n373_), .A2(new_n385_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n403_), .B1(new_n404_), .B2(new_n398_), .ZN(new_n405_));
  AND4_X1   g204(.A1(new_n369_), .A2(new_n405_), .A3(new_n401_), .A4(new_n386_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n365_), .B1(new_n402_), .B2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n395_), .A2(new_n369_), .A3(new_n401_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n382_), .B1(new_n233_), .B2(new_n379_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n400_), .B1(new_n297_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(new_n371_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n411_), .B1(new_n371_), .B2(new_n393_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n369_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n365_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n408_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n407_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n342_), .A2(new_n364_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT100), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n419_), .A2(KEYINPUT33), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n360_), .B(new_n420_), .C1(new_n351_), .C2(new_n355_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(KEYINPUT33), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n348_), .A2(new_n350_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n352_), .A2(new_n349_), .A3(new_n354_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n424_), .A2(new_n425_), .A3(new_n361_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n405_), .A2(new_n401_), .A3(new_n386_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n413_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n423_), .A2(new_n426_), .A3(new_n428_), .A4(new_n408_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n421_), .A2(new_n422_), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n369_), .A2(KEYINPUT32), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n412_), .A2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n432_), .B1(new_n427_), .B2(new_n431_), .ZN(new_n433_));
  OAI22_X1  g232(.A1(new_n429_), .A2(new_n430_), .B1(new_n364_), .B2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n434_), .A2(new_n335_), .A3(new_n341_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n248_), .B1(new_n418_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n364_), .ZN(new_n437_));
  NOR4_X1   g236(.A1(new_n342_), .A2(new_n437_), .A3(new_n416_), .A4(new_n247_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT68), .ZN(new_n440_));
  AND2_X1   g239(.A1(G85gat), .A2(G92gat), .ZN(new_n441_));
  NOR2_X1   g240(.A1(G85gat), .A2(G92gat), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT8), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT67), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NOR3_X1   g247(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n446_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  OR3_X1    g249(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n451_), .A2(KEYINPUT67), .A3(new_n447_), .ZN(new_n452_));
  AND2_X1   g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G99gat), .A2(G106gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT6), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT6), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n456_), .A2(G99gat), .A3(G106gat), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT66), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n455_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n458_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n445_), .B1(new_n453_), .B2(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n448_), .A2(new_n449_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n455_), .A2(new_n457_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n443_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n466_), .B1(G85gat), .B2(G92gat), .ZN(new_n467_));
  AND2_X1   g266(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n468_));
  NOR2_X1   g267(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n469_));
  OAI21_X1  g268(.A(G85gat), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  AND2_X1   g269(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n471_));
  NOR2_X1   g270(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n467_), .B1(new_n470_), .B2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT10), .B(G99gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n464_), .B1(new_n475_), .B2(G106gat), .ZN(new_n476_));
  OAI22_X1  g275(.A1(new_n465_), .A2(KEYINPUT8), .B1(new_n474_), .B2(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n440_), .B1(new_n462_), .B2(new_n477_), .ZN(new_n478_));
  XOR2_X1   g277(.A(G71gat), .B(G78gat), .Z(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G57gat), .B(G64gat), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT69), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(G57gat), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n484_), .A2(G64gat), .ZN(new_n485_));
  INV_X1    g284(.A(G64gat), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n486_), .A2(G57gat), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT69), .B1(new_n485_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n483_), .A2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n480_), .B1(new_n489_), .B2(KEYINPUT11), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT11), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n483_), .A2(new_n488_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  AOI211_X1 g292(.A(new_n491_), .B(new_n479_), .C1(new_n483_), .C2(new_n488_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n464_), .A2(KEYINPUT66), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n455_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n497_), .A2(new_n450_), .A3(new_n452_), .A4(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT8), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n443_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n464_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n451_), .A2(new_n447_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n444_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(new_n500_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n475_), .ZN(new_n507_));
  INV_X1    g306(.A(G106gat), .ZN(new_n508_));
  AOI22_X1  g307(.A1(new_n507_), .A2(new_n508_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n470_), .A2(new_n473_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n467_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n509_), .A2(new_n512_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n502_), .A2(new_n506_), .A3(KEYINPUT68), .A4(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n478_), .A2(new_n496_), .A3(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n494_), .B1(new_n492_), .B2(new_n490_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n502_), .A2(new_n513_), .A3(new_n506_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n516_), .A2(new_n517_), .A3(KEYINPUT12), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n496_), .B1(new_n478_), .B2(new_n514_), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n515_), .B(new_n518_), .C1(new_n519_), .C2(KEYINPUT12), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G230gat), .A2(G233gat), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n478_), .A2(new_n514_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(new_n516_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n521_), .B1(new_n525_), .B2(new_n515_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n523_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G120gat), .B(G148gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT5), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G176gat), .B(G204gat), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n529_), .B(new_n530_), .Z(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n527_), .A2(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n531_), .B1(new_n523_), .B2(new_n526_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT13), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G29gat), .B(G36gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT70), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G43gat), .B(G50gat), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n538_), .A2(KEYINPUT70), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n538_), .A2(KEYINPUT70), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(new_n544_), .A3(new_n540_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n542_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G15gat), .B(G22gat), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G1gat), .A2(G8gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT14), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G1gat), .B(G8gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n546_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n542_), .A2(new_n545_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n555_), .A2(new_n552_), .ZN(new_n556_));
  OAI211_X1 g355(.A(G229gat), .B(G233gat), .C1(new_n554_), .C2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT71), .B(KEYINPUT15), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n555_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n542_), .A2(new_n545_), .A3(new_n558_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n560_), .A2(new_n552_), .A3(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G229gat), .A2(G233gat), .ZN(new_n563_));
  INV_X1    g362(.A(new_n556_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n562_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G113gat), .B(G141gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G169gat), .B(G197gat), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n566_), .B(new_n567_), .Z(new_n568_));
  AND3_X1   g367(.A1(new_n557_), .A2(new_n565_), .A3(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n568_), .B1(new_n557_), .B2(new_n565_), .ZN(new_n570_));
  OAI21_X1  g369(.A(KEYINPUT79), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n557_), .A2(new_n565_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n568_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT79), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n557_), .A2(new_n565_), .A3(new_n568_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n574_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n571_), .A2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n533_), .A2(KEYINPUT13), .A3(new_n534_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n537_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n439_), .A2(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(KEYINPUT72), .B1(new_n524_), .B2(new_n555_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT34), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n584_), .A2(KEYINPUT35), .ZN(new_n585_));
  INV_X1    g384(.A(new_n561_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n558_), .B1(new_n542_), .B2(new_n545_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n585_), .B1(new_n588_), .B2(new_n517_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT72), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n478_), .A2(new_n590_), .A3(new_n546_), .A4(new_n514_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n582_), .A2(new_n589_), .A3(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n592_), .A2(KEYINPUT35), .A3(new_n584_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G190gat), .B(G218gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT73), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G134gat), .B(G162gat), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n595_), .B(new_n596_), .Z(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n598_), .A2(KEYINPUT36), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n584_), .A2(KEYINPUT35), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n589_), .A2(new_n582_), .A3(new_n600_), .A4(new_n591_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n593_), .A2(new_n599_), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT74), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT74), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n593_), .A2(new_n604_), .A3(new_n599_), .A4(new_n601_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n593_), .A2(new_n601_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n597_), .B(KEYINPUT36), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n606_), .A2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(KEYINPUT75), .B(KEYINPUT37), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n606_), .A2(new_n609_), .A3(new_n611_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n516_), .B(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT76), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n619_), .A2(new_n552_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n617_), .B(KEYINPUT76), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n621_), .A2(new_n553_), .ZN(new_n622_));
  OAI21_X1  g421(.A(KEYINPUT77), .B1(new_n620_), .B2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n553_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n619_), .A2(new_n552_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT77), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n624_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(G127gat), .B(G155gat), .Z(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT16), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G183gat), .B(G211gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT17), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n623_), .A2(new_n627_), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT78), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n635_), .B1(new_n620_), .B2(new_n622_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n624_), .A2(new_n625_), .A3(KEYINPUT78), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n631_), .B(KEYINPUT17), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n636_), .A2(new_n637_), .A3(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n634_), .A2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n615_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n581_), .A2(new_n641_), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n642_), .A2(G1gat), .A3(new_n364_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT38), .Z(new_n644_));
  INV_X1    g443(.A(new_n610_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n439_), .A2(new_n640_), .A3(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n580_), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n647_), .A2(KEYINPUT101), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(KEYINPUT101), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n646_), .A2(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(G1gat), .B1(new_n651_), .B2(new_n364_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n644_), .A2(new_n652_), .ZN(G1324gat));
  OAI21_X1  g452(.A(G8gat), .B1(new_n651_), .B2(new_n417_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT39), .Z(new_n655_));
  NOR3_X1   g454(.A1(new_n642_), .A2(G8gat), .A3(new_n417_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT40), .ZN(G1325gat));
  OAI21_X1  g457(.A(G15gat), .B1(new_n651_), .B2(new_n247_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT41), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n642_), .A2(G15gat), .A3(new_n247_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT102), .ZN(G1326gat));
  INV_X1    g462(.A(new_n342_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G22gat), .B1(new_n651_), .B2(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT42), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n664_), .A2(G22gat), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n666_), .B1(new_n642_), .B2(new_n667_), .ZN(G1327gat));
  INV_X1    g467(.A(new_n640_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n669_), .A2(new_n610_), .ZN(new_n670_));
  OAI211_X1 g469(.A(new_n647_), .B(new_n670_), .C1(new_n436_), .C2(new_n438_), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n671_), .A2(KEYINPUT106), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(KEYINPUT106), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(G29gat), .B1(new_n674_), .B2(new_n437_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n676_));
  INV_X1    g475(.A(new_n615_), .ZN(new_n677_));
  AOI211_X1 g476(.A(new_n437_), .B(new_n416_), .C1(new_n335_), .C2(new_n341_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n434_), .A2(new_n335_), .A3(new_n341_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n247_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n438_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n677_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT104), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n676_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n615_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n686_), .A2(KEYINPUT104), .A3(KEYINPUT43), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n684_), .A2(new_n685_), .A3(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n669_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(KEYINPUT105), .B1(new_n690_), .B2(new_n691_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n688_), .A2(new_n689_), .A3(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n689_), .B1(new_n688_), .B2(new_n694_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n437_), .A2(G29gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n675_), .B1(new_n698_), .B2(new_n699_), .ZN(G1328gat));
  INV_X1    g499(.A(G36gat), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n417_), .A2(KEYINPUT107), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n417_), .A2(KEYINPUT107), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n672_), .A2(new_n701_), .A3(new_n673_), .A4(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT45), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n705_), .B(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n416_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n708_), .B2(G36gat), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT46), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n710_), .A2(KEYINPUT108), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(KEYINPUT108), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT109), .Z(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n709_), .A2(new_n711_), .A3(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n705_), .B(KEYINPUT45), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n686_), .A2(KEYINPUT104), .A3(KEYINPUT43), .ZN(new_n717_));
  AOI21_X1  g516(.A(KEYINPUT43), .B1(new_n686_), .B2(KEYINPUT104), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n717_), .A2(new_n718_), .A3(KEYINPUT105), .ZN(new_n719_));
  INV_X1    g518(.A(new_n694_), .ZN(new_n720_));
  OAI21_X1  g519(.A(KEYINPUT44), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n688_), .A2(new_n689_), .A3(new_n694_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n417_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n716_), .B1(new_n723_), .B2(new_n701_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n711_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n713_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n715_), .A2(new_n726_), .ZN(G1329gat));
  AOI21_X1  g526(.A(G43gat), .B1(new_n674_), .B2(new_n248_), .ZN(new_n728_));
  XOR2_X1   g527(.A(new_n728_), .B(KEYINPUT110), .Z(new_n729_));
  NAND2_X1  g528(.A1(new_n248_), .A2(G43gat), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n697_), .A2(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(KEYINPUT47), .B1(new_n729_), .B2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n728_), .B(KEYINPUT110), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT47), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n733_), .B(new_n734_), .C1(new_n697_), .C2(new_n730_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n732_), .A2(new_n735_), .ZN(G1330gat));
  INV_X1    g535(.A(G50gat), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n674_), .A2(new_n737_), .A3(new_n342_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n342_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n739_), .A2(new_n740_), .A3(G50gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n740_), .B1(new_n739_), .B2(G50gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n738_), .B1(new_n741_), .B2(new_n742_), .ZN(G1331gat));
  NAND2_X1  g542(.A1(new_n537_), .A2(new_n579_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  NOR3_X1   g544(.A1(new_n439_), .A2(new_n578_), .A3(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(new_n641_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n484_), .B1(new_n747_), .B2(new_n364_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n578_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n646_), .A2(new_n749_), .A3(new_n744_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT112), .ZN(new_n751_));
  OAI21_X1  g550(.A(G57gat), .B1(new_n364_), .B2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n752_), .B1(new_n751_), .B2(G57gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n748_), .B1(new_n750_), .B2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT113), .ZN(G1332gat));
  INV_X1    g554(.A(new_n704_), .ZN(new_n756_));
  OAI21_X1  g555(.A(G64gat), .B1(new_n750_), .B2(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT48), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n704_), .A2(new_n486_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n758_), .B1(new_n747_), .B2(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT114), .ZN(G1333gat));
  OAI21_X1  g560(.A(G71gat), .B1(new_n750_), .B2(new_n247_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT49), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n247_), .A2(G71gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n747_), .B2(new_n764_), .ZN(G1334gat));
  OAI21_X1  g564(.A(G78gat), .B1(new_n750_), .B2(new_n664_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT50), .ZN(new_n767_));
  OR2_X1    g566(.A1(new_n664_), .A2(G78gat), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n747_), .B2(new_n768_), .ZN(G1335gat));
  INV_X1    g568(.A(G85gat), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n746_), .A2(new_n670_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(new_n364_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT115), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n684_), .A2(new_n687_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n669_), .A2(new_n745_), .A3(new_n578_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n776_), .A2(new_n770_), .A3(new_n364_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n773_), .A2(new_n777_), .ZN(G1336gat));
  NOR2_X1   g577(.A1(new_n468_), .A2(new_n469_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n776_), .A2(new_n779_), .A3(new_n756_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n771_), .ZN(new_n781_));
  AOI21_X1  g580(.A(G92gat), .B1(new_n781_), .B2(new_n416_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n780_), .A2(new_n782_), .ZN(G1337gat));
  NOR2_X1   g582(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n784_));
  OAI21_X1  g583(.A(G99gat), .B1(new_n776_), .B2(new_n247_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n781_), .A2(new_n507_), .A3(new_n248_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n784_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(KEYINPUT116), .A2(KEYINPUT51), .ZN(new_n788_));
  XOR2_X1   g587(.A(new_n787_), .B(new_n788_), .Z(G1338gat));
  NAND3_X1  g588(.A1(new_n781_), .A2(new_n508_), .A3(new_n342_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n774_), .A2(new_n342_), .A3(new_n775_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n791_), .A2(new_n792_), .A3(G106gat), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n791_), .B2(G106gat), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n790_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n634_), .A2(new_n639_), .A3(new_n749_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(new_n799_), .A3(new_n745_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n634_), .A2(new_n639_), .A3(new_n749_), .ZN(new_n801_));
  OAI21_X1  g600(.A(KEYINPUT117), .B1(new_n801_), .B2(new_n744_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n797_), .B1(new_n803_), .B2(new_n677_), .ZN(new_n804_));
  AOI211_X1 g603(.A(KEYINPUT54), .B(new_n615_), .C1(new_n800_), .C2(new_n802_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  OR2_X1    g605(.A1(new_n554_), .A2(new_n556_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n568_), .B1(new_n807_), .B2(new_n563_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n562_), .A2(new_n564_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n808_), .B1(new_n563_), .B2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n576_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n527_), .B2(new_n532_), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT12), .B1(new_n524_), .B2(new_n516_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n515_), .A2(new_n518_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n522_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT118), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT118), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n520_), .A2(new_n819_), .A3(new_n522_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT12), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n525_), .A2(new_n821_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n515_), .A2(new_n518_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n822_), .A2(new_n823_), .A3(KEYINPUT55), .A4(new_n521_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n816_), .A2(new_n818_), .A3(new_n820_), .A4(new_n824_), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n825_), .A2(KEYINPUT56), .A3(new_n531_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT56), .B1(new_n825_), .B2(new_n531_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n812_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT58), .ZN(new_n829_));
  OR2_X1    g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n829_), .ZN(new_n831_));
  AND3_X1   g630(.A1(new_n830_), .A2(new_n615_), .A3(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n811_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  NOR3_X1   g633(.A1(new_n826_), .A2(new_n827_), .A3(KEYINPUT119), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n825_), .A2(KEYINPUT119), .A3(KEYINPUT56), .A4(new_n531_), .ZN(new_n836_));
  AOI22_X1  g635(.A1(new_n571_), .A2(new_n577_), .B1(new_n527_), .B2(new_n532_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n834_), .B1(new_n835_), .B2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(KEYINPUT57), .A3(new_n610_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n825_), .A2(new_n531_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT56), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT119), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n825_), .A2(KEYINPUT56), .A3(new_n531_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n845_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n836_), .A2(new_n837_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n645_), .B1(new_n850_), .B2(new_n834_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n851_), .A2(KEYINPUT121), .A3(KEYINPUT57), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n832_), .B1(new_n842_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n833_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n645_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n853_), .A2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n806_), .B1(new_n857_), .B2(new_n640_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n342_), .A2(new_n247_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n859_), .A2(new_n437_), .A3(new_n417_), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n858_), .A2(KEYINPUT59), .A3(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT120), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n856_), .A2(new_n862_), .ZN(new_n863_));
  OAI211_X1 g662(.A(KEYINPUT120), .B(new_n854_), .C1(new_n855_), .C2(new_n645_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n669_), .B1(new_n853_), .B2(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(KEYINPUT122), .B1(new_n866_), .B2(new_n806_), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n863_), .A2(new_n864_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n830_), .A2(new_n615_), .A3(new_n831_), .ZN(new_n869_));
  AOI21_X1  g668(.A(KEYINPUT121), .B1(new_n851_), .B2(KEYINPUT57), .ZN(new_n870_));
  NOR4_X1   g669(.A1(new_n855_), .A2(new_n841_), .A3(new_n854_), .A4(new_n645_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n869_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n640_), .B1(new_n868_), .B2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n874_));
  INV_X1    g673(.A(new_n806_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n873_), .A2(new_n874_), .A3(new_n875_), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n867_), .A2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n860_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  AOI211_X1 g678(.A(new_n749_), .B(new_n861_), .C1(new_n879_), .C2(KEYINPUT59), .ZN(new_n880_));
  INV_X1    g679(.A(G113gat), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n578_), .A2(new_n881_), .ZN(new_n882_));
  OAI22_X1  g681(.A1(new_n880_), .A2(new_n881_), .B1(new_n879_), .B2(new_n882_), .ZN(G1340gat));
  INV_X1    g682(.A(new_n879_), .ZN(new_n884_));
  INV_X1    g683(.A(G120gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n885_), .B1(new_n745_), .B2(KEYINPUT60), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n884_), .B(new_n886_), .C1(KEYINPUT60), .C2(new_n885_), .ZN(new_n887_));
  AOI211_X1 g686(.A(new_n745_), .B(new_n861_), .C1(new_n879_), .C2(KEYINPUT59), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n888_), .B2(new_n885_), .ZN(G1341gat));
  INV_X1    g688(.A(G127gat), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n884_), .A2(new_n890_), .A3(new_n669_), .ZN(new_n891_));
  AOI211_X1 g690(.A(new_n640_), .B(new_n861_), .C1(new_n879_), .C2(KEYINPUT59), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(new_n890_), .ZN(G1342gat));
  INV_X1    g692(.A(G134gat), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n884_), .A2(new_n894_), .A3(new_n645_), .ZN(new_n895_));
  AOI211_X1 g694(.A(new_n677_), .B(new_n861_), .C1(new_n879_), .C2(KEYINPUT59), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n896_), .B2(new_n894_), .ZN(G1343gat));
  NOR4_X1   g696(.A1(new_n704_), .A2(new_n364_), .A3(new_n664_), .A4(new_n248_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n877_), .A2(new_n578_), .A3(new_n898_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g699(.A1(new_n877_), .A2(new_n744_), .A3(new_n898_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g701(.A1(new_n877_), .A2(new_n669_), .A3(new_n898_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(KEYINPUT61), .B(G155gat), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1346gat));
  NAND4_X1  g704(.A1(new_n877_), .A2(G162gat), .A3(new_n615_), .A4(new_n898_), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n867_), .A2(new_n876_), .A3(new_n645_), .A4(new_n898_), .ZN(new_n907_));
  AND3_X1   g706(.A1(new_n907_), .A2(KEYINPUT123), .A3(new_n254_), .ZN(new_n908_));
  AOI21_X1  g707(.A(KEYINPUT123), .B1(new_n907_), .B2(new_n254_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n906_), .B1(new_n908_), .B2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  OAI211_X1 g711(.A(KEYINPUT124), .B(new_n906_), .C1(new_n908_), .C2(new_n909_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1347gat));
  NOR2_X1   g713(.A1(new_n756_), .A2(new_n437_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n859_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n858_), .A2(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n578_), .ZN(new_n918_));
  XOR2_X1   g717(.A(KEYINPUT22), .B(G169gat), .Z(new_n919_));
  NOR2_X1   g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n918_), .A2(G169gat), .A3(new_n921_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n920_), .B1(new_n922_), .B2(new_n923_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n924_), .B1(new_n922_), .B2(new_n923_), .ZN(G1348gat));
  INV_X1    g724(.A(G176gat), .ZN(new_n926_));
  INV_X1    g725(.A(new_n917_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n927_), .B2(new_n745_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT126), .ZN(new_n929_));
  OR2_X1    g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n928_), .A2(new_n929_), .ZN(new_n931_));
  AND2_X1   g730(.A1(new_n877_), .A2(new_n664_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n915_), .A2(new_n248_), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n933_), .A2(new_n926_), .A3(new_n745_), .ZN(new_n934_));
  AOI22_X1  g733(.A1(new_n930_), .A2(new_n931_), .B1(new_n932_), .B2(new_n934_), .ZN(G1349gat));
  NOR2_X1   g734(.A1(new_n933_), .A2(new_n640_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n877_), .A2(new_n664_), .A3(new_n936_), .ZN(new_n937_));
  INV_X1    g736(.A(G183gat), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n937_), .A2(new_n938_), .ZN(new_n939_));
  OR3_X1    g738(.A1(new_n927_), .A2(new_n223_), .A3(new_n640_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT127), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n941_), .A2(new_n942_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n939_), .A2(new_n940_), .A3(KEYINPUT127), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n943_), .A2(new_n944_), .ZN(G1350gat));
  OAI21_X1  g744(.A(G190gat), .B1(new_n927_), .B2(new_n677_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n917_), .A2(new_n224_), .A3(new_n645_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n946_), .A2(new_n947_), .ZN(G1351gat));
  NOR4_X1   g747(.A1(new_n756_), .A2(new_n437_), .A3(new_n664_), .A4(new_n248_), .ZN(new_n949_));
  AND2_X1   g748(.A1(new_n877_), .A2(new_n949_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n950_), .A2(new_n578_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n951_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g751(.A1(new_n950_), .A2(new_n744_), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n953_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g753(.A1(new_n877_), .A2(new_n669_), .A3(new_n949_), .ZN(new_n955_));
  NOR2_X1   g754(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n956_));
  AND2_X1   g755(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n957_));
  NOR3_X1   g756(.A1(new_n955_), .A2(new_n956_), .A3(new_n957_), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n958_), .B1(new_n955_), .B2(new_n956_), .ZN(G1354gat));
  INV_X1    g758(.A(G218gat), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n950_), .A2(new_n960_), .A3(new_n645_), .ZN(new_n961_));
  AND2_X1   g760(.A1(new_n950_), .A2(new_n615_), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n961_), .B1(new_n962_), .B2(new_n960_), .ZN(G1355gat));
endmodule


