//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 0 0 1 0 0 1 1 0 1 0 0 1 1 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n776_, new_n777_, new_n778_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n813_, new_n814_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n918_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n944_, new_n945_, new_n947_, new_n948_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n955_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n978_, new_n979_;
  XOR2_X1   g000(.A(G1gat), .B(G29gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT99), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT0), .B(G57gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT84), .ZN(new_n208_));
  OR2_X1    g007(.A1(KEYINPUT82), .A2(KEYINPUT83), .ZN(new_n209_));
  NAND2_X1  g008(.A1(KEYINPUT82), .A2(KEYINPUT83), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(G127gat), .A2(G134gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G127gat), .A2(G134gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G127gat), .B(G134gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(G113gat), .B(G120gat), .ZN(new_n217_));
  AND3_X1   g016(.A1(new_n214_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n217_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n208_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n214_), .A2(new_n216_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n217_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n214_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(KEYINPUT84), .A3(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT86), .ZN(new_n226_));
  OAI22_X1  g025(.A1(new_n226_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G141gat), .A2(G148gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT2), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  AND3_X1   g030(.A1(new_n227_), .A2(new_n228_), .A3(new_n231_), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n226_), .A2(KEYINPUT3), .ZN(new_n233_));
  NOR2_X1   g032(.A1(G141gat), .A2(G148gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n226_), .A2(KEYINPUT3), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n233_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n232_), .A2(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(G155gat), .A2(G162gat), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G155gat), .A2(G162gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n237_), .A2(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n240_), .A2(KEYINPUT1), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n240_), .A2(KEYINPUT1), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(new_n239_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n229_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n247_), .A2(new_n234_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n243_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n220_), .A2(new_n225_), .A3(new_n250_), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n243_), .B(new_n249_), .C1(new_n218_), .C2(new_n219_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n251_), .A2(KEYINPUT4), .A3(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT4), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n220_), .A2(new_n225_), .A3(new_n254_), .A4(new_n250_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G225gat), .A2(G233gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT98), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n253_), .A2(new_n255_), .A3(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n251_), .A2(new_n252_), .A3(new_n256_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n207_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  AND3_X1   g060(.A1(new_n251_), .A2(KEYINPUT4), .A3(new_n252_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n255_), .A2(new_n257_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n259_), .B(new_n207_), .C1(new_n262_), .C2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n261_), .A2(new_n264_), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n220_), .A2(new_n225_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT31), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n266_), .A2(new_n267_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT25), .ZN(new_n272_));
  INV_X1    g071(.A(G183gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT78), .B(G183gat), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n274_), .B1(new_n275_), .B2(new_n272_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT26), .B(G190gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(G169gat), .ZN(new_n279_));
  INV_X1    g078(.A(G176gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n281_), .A2(KEYINPUT24), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT24), .ZN(new_n284_));
  NOR2_X1   g083(.A1(G169gat), .A2(G176gat), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT79), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT79), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n281_), .A2(new_n287_), .A3(KEYINPUT24), .A4(new_n283_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n282_), .B1(new_n286_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G183gat), .A2(G190gat), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT23), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(KEYINPUT80), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT80), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n294_), .A2(G183gat), .A3(G190gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n292_), .B1(new_n296_), .B2(new_n291_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n278_), .A2(new_n289_), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT81), .ZN(new_n299_));
  INV_X1    g098(.A(new_n283_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT22), .B(G169gat), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n300_), .B1(new_n301_), .B2(new_n280_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n290_), .A2(KEYINPUT23), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n303_), .B1(new_n296_), .B2(KEYINPUT23), .ZN(new_n304_));
  INV_X1    g103(.A(G190gat), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n275_), .A2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n302_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n298_), .A2(new_n299_), .A3(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n299_), .B1(new_n298_), .B2(new_n307_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(G15gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n298_), .A2(new_n307_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT81), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n298_), .A2(new_n299_), .A3(new_n307_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(G15gat), .ZN(new_n317_));
  XOR2_X1   g116(.A(G71gat), .B(G99gat), .Z(new_n318_));
  NAND2_X1  g117(.A1(G227gat), .A2(G233gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT30), .B(G43gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n312_), .A2(new_n317_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT85), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n322_), .B1(new_n312_), .B2(new_n317_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n271_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n312_), .A2(new_n317_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n322_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n330_), .A2(new_n324_), .A3(new_n323_), .A4(new_n270_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n327_), .A2(new_n331_), .ZN(new_n332_));
  OR3_X1    g131(.A1(new_n250_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT28), .B1(new_n250_), .B2(KEYINPUT29), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G22gat), .B(G50gat), .ZN(new_n335_));
  AND3_X1   g134(.A1(new_n333_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n335_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n249_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n241_), .B1(new_n232_), .B2(new_n236_), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT29), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G211gat), .B(G218gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT89), .ZN(new_n343_));
  INV_X1    g142(.A(G197gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(KEYINPUT89), .A2(G197gat), .ZN(new_n346_));
  AOI21_X1  g145(.A(G204gat), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(G204gat), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT21), .B1(new_n344_), .B2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n342_), .B1(new_n347_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n346_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(KEYINPUT89), .A2(G197gat), .ZN(new_n352_));
  OAI21_X1  g151(.A(G204gat), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT21), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n344_), .A2(G204gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n353_), .A2(new_n354_), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT90), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n345_), .A2(new_n346_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n355_), .B1(new_n359_), .B2(G204gat), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT90), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(new_n361_), .A3(new_n354_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n350_), .B1(new_n358_), .B2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n353_), .A2(KEYINPUT91), .A3(new_n356_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n342_), .A2(new_n354_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n360_), .A2(KEYINPUT91), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n341_), .B1(new_n363_), .B2(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT87), .B(G228gat), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT88), .B(G233gat), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n369_), .A2(new_n374_), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n341_), .B(new_n373_), .C1(new_n363_), .C2(new_n368_), .ZN(new_n376_));
  XOR2_X1   g175(.A(G78gat), .B(G106gat), .Z(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT92), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT92), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n375_), .A2(new_n380_), .A3(new_n376_), .A4(new_n377_), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT93), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n375_), .A2(new_n376_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n377_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n383_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  AOI211_X1 g185(.A(KEYINPUT93), .B(new_n377_), .C1(new_n375_), .C2(new_n376_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n338_), .B1(new_n382_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n358_), .A2(new_n362_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n350_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  OR2_X1    g191(.A1(new_n366_), .A2(new_n367_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n373_), .B1(new_n394_), .B2(new_n341_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n376_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n385_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n338_), .A2(new_n378_), .A3(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n332_), .B1(new_n389_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n397_), .A2(KEYINPUT93), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n384_), .A2(new_n383_), .A3(new_n385_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n401_), .A2(new_n379_), .A3(new_n381_), .A4(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n338_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n405_), .A2(new_n398_), .A3(new_n331_), .A4(new_n327_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n265_), .B1(new_n400_), .B2(new_n406_), .ZN(new_n407_));
  XOR2_X1   g206(.A(KEYINPUT106), .B(KEYINPUT27), .Z(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n284_), .A2(new_n285_), .ZN(new_n410_));
  NOR3_X1   g209(.A1(new_n304_), .A2(new_n410_), .A3(new_n282_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n277_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT25), .B(G183gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT95), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n411_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n273_), .A2(new_n305_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n297_), .A2(new_n416_), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n417_), .A2(KEYINPUT96), .A3(new_n302_), .ZN(new_n418_));
  AOI21_X1  g217(.A(KEYINPUT96), .B1(new_n417_), .B2(new_n302_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n415_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n394_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n363_), .A2(new_n368_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n314_), .A2(new_n422_), .A3(new_n315_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(new_n423_), .A3(KEYINPUT20), .ZN(new_n424_));
  AND3_X1   g223(.A1(KEYINPUT19), .A2(G226gat), .A3(G233gat), .ZN(new_n425_));
  AOI21_X1  g224(.A(KEYINPUT19), .B1(G226gat), .B2(G233gat), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  XOR2_X1   g226(.A(new_n427_), .B(KEYINPUT94), .Z(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT20), .B1(new_n425_), .B2(new_n426_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n430_), .B1(new_n316_), .B2(new_n394_), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n420_), .A2(new_n394_), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n424_), .A2(new_n429_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G64gat), .B(G92gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G8gat), .B(G36gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  OR2_X1    g237(.A1(new_n433_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n424_), .A2(new_n429_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n431_), .A2(new_n432_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(new_n441_), .A3(new_n438_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n409_), .B1(new_n439_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(KEYINPUT27), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n421_), .A2(new_n423_), .A3(KEYINPUT20), .A4(new_n428_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT102), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT20), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n447_), .B1(new_n310_), .B2(new_n422_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT102), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n448_), .A2(new_n449_), .A3(new_n428_), .A4(new_n421_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n417_), .A2(new_n302_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n422_), .A2(new_n415_), .A3(new_n451_), .ZN(new_n452_));
  XOR2_X1   g251(.A(KEYINPUT101), .B(KEYINPUT20), .Z(new_n453_));
  OAI211_X1 g252(.A(new_n452_), .B(new_n453_), .C1(new_n310_), .C2(new_n422_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n427_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n446_), .A2(new_n450_), .A3(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(new_n438_), .B(KEYINPUT104), .Z(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n444_), .B1(new_n458_), .B2(KEYINPUT105), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT105), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n456_), .A2(new_n460_), .A3(new_n457_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n443_), .B1(new_n459_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT33), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n253_), .A2(new_n256_), .A3(new_n255_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n251_), .A2(new_n252_), .A3(new_n257_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n465_), .A2(new_n206_), .ZN(new_n466_));
  AOI22_X1  g265(.A1(new_n264_), .A2(new_n463_), .B1(new_n464_), .B2(new_n466_), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n251_), .A2(new_n252_), .A3(new_n256_), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n255_), .A2(new_n257_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n468_), .B1(new_n253_), .B2(new_n469_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n470_), .A2(KEYINPUT100), .A3(KEYINPUT33), .A4(new_n207_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n258_), .A2(KEYINPUT33), .A3(new_n259_), .A4(new_n207_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT100), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n467_), .A2(new_n471_), .A3(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n438_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n433_), .B(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT103), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n440_), .A2(new_n441_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n438_), .A2(KEYINPUT32), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n264_), .ZN(new_n483_));
  OAI22_X1  g282(.A1(new_n480_), .A2(new_n482_), .B1(new_n483_), .B2(new_n260_), .ZN(new_n484_));
  AOI22_X1  g283(.A1(new_n445_), .A2(KEYINPUT102), .B1(new_n454_), .B2(new_n427_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n481_), .B1(new_n485_), .B2(new_n450_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n479_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n456_), .A2(new_n482_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n433_), .A2(new_n481_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n488_), .A2(KEYINPUT103), .A3(new_n265_), .A4(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n478_), .A2(new_n487_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n405_), .A2(new_n398_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n332_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  AOI22_X1  g293(.A1(new_n407_), .A2(new_n462_), .B1(new_n491_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G230gat), .A2(G233gat), .ZN(new_n496_));
  XOR2_X1   g295(.A(new_n496_), .B(KEYINPUT64), .Z(new_n497_));
  XNOR2_X1  g296(.A(G57gat), .B(G64gat), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n498_), .A2(KEYINPUT11), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(KEYINPUT11), .ZN(new_n500_));
  XOR2_X1   g299(.A(G71gat), .B(G78gat), .Z(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n500_), .A2(new_n501_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT66), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NOR3_X1   g306(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n505_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G99gat), .A2(G106gat), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT6), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT7), .ZN(new_n515_));
  INV_X1    g314(.A(G99gat), .ZN(new_n516_));
  INV_X1    g315(.A(G106gat), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n515_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n518_), .A2(KEYINPUT66), .A3(new_n506_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n509_), .A2(new_n514_), .A3(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT8), .ZN(new_n521_));
  INV_X1    g320(.A(G92gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(G85gat), .ZN(new_n523_));
  INV_X1    g322(.A(G85gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(G92gat), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n521_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n520_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n523_), .A2(new_n525_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n518_), .A2(new_n506_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n512_), .A2(new_n513_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n528_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(new_n521_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n527_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT10), .B(G99gat), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n514_), .B1(G106gat), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT9), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n536_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n537_));
  NOR3_X1   g336(.A1(new_n524_), .A2(new_n522_), .A3(KEYINPUT9), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT65), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n524_), .A2(G92gat), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n522_), .A2(G85gat), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT9), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n538_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT65), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n535_), .B1(new_n539_), .B2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n504_), .B1(new_n533_), .B2(new_n546_), .ZN(new_n547_));
  AOI22_X1  g346(.A1(new_n520_), .A2(new_n526_), .B1(new_n531_), .B2(new_n521_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n534_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n530_), .B1(new_n549_), .B2(new_n517_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n544_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n551_));
  NOR3_X1   g350(.A1(new_n537_), .A2(KEYINPUT65), .A3(new_n538_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n550_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n502_), .A2(new_n503_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n548_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n547_), .A2(KEYINPUT12), .A3(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n548_), .A2(new_n553_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT12), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(new_n558_), .A3(new_n504_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n497_), .B1(new_n556_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n497_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n561_), .B1(new_n547_), .B2(new_n555_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G120gat), .B(G148gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(new_n348_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(KEYINPUT5), .B(G176gat), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n564_), .B(new_n565_), .Z(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n560_), .A2(new_n562_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n567_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT13), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n569_), .A2(KEYINPUT13), .A3(new_n570_), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G113gat), .B(G141gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G169gat), .B(G197gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G229gat), .A2(G233gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G15gat), .B(G22gat), .ZN(new_n581_));
  INV_X1    g380(.A(G1gat), .ZN(new_n582_));
  INV_X1    g381(.A(G8gat), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT14), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G1gat), .B(G8gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  XOR2_X1   g387(.A(G29gat), .B(G36gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(G43gat), .B(G50gat), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(G43gat), .B(G50gat), .Z(new_n592_));
  XNOR2_X1  g391(.A(G29gat), .B(G36gat), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n591_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n588_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n587_), .A2(new_n595_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT76), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n597_), .A2(KEYINPUT76), .A3(new_n598_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n580_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(KEYINPUT68), .B(KEYINPUT15), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n595_), .B(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(new_n587_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n606_), .A2(new_n580_), .A3(new_n597_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n579_), .B1(new_n603_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT77), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n603_), .A2(new_n607_), .A3(new_n579_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n609_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n611_), .ZN(new_n613_));
  AOI21_X1  g412(.A(KEYINPUT77), .B1(new_n613_), .B2(new_n608_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n495_), .A2(new_n576_), .A3(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(G127gat), .B(G155gat), .Z(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(G211gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT16), .B(G183gat), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n618_), .B(new_n619_), .Z(new_n620_));
  AND2_X1   g419(.A1(new_n620_), .A2(KEYINPUT17), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT74), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n622_), .B1(KEYINPUT17), .B2(new_n620_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n588_), .B(new_n554_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G231gat), .A2(G233gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT75), .ZN(new_n627_));
  OR2_X1    g426(.A1(KEYINPUT74), .A2(KEYINPUT17), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n627_), .B1(new_n620_), .B2(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n623_), .B1(new_n626_), .B2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n621_), .A2(new_n627_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n626_), .A2(new_n631_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(KEYINPUT67), .B(KEYINPUT34), .ZN(new_n634_));
  NAND2_X1  g433(.A1(G232gat), .A2(G233gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT35), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n605_), .A2(new_n557_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n638_), .B1(new_n639_), .B2(KEYINPUT69), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n605_), .A2(new_n557_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n548_), .A2(new_n553_), .A3(new_n596_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(new_n643_), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n641_), .A2(KEYINPUT69), .A3(new_n642_), .A4(new_n638_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n636_), .A2(new_n637_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n644_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(G190gat), .B(G218gat), .ZN(new_n648_));
  INV_X1    g447(.A(G162gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(KEYINPUT70), .B(G134gat), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n648_), .B(G162gat), .ZN(new_n653_));
  INV_X1    g452(.A(new_n651_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n652_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT36), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n647_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT71), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n652_), .A2(new_n655_), .A3(KEYINPUT36), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n658_), .A2(KEYINPUT72), .A3(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT72), .B1(new_n658_), .B2(new_n663_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n644_), .A2(new_n645_), .A3(new_n646_), .A4(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT73), .ZN(new_n668_));
  AOI22_X1  g467(.A1(new_n640_), .A2(new_n643_), .B1(new_n637_), .B2(new_n636_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT73), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n669_), .A2(new_n670_), .A3(new_n645_), .A4(new_n666_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n647_), .A2(KEYINPUT71), .A3(new_n659_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n662_), .A2(new_n668_), .A3(new_n671_), .A4(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT37), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n669_), .A2(new_n658_), .A3(new_n645_), .A4(new_n663_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT37), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n660_), .A2(new_n675_), .A3(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n633_), .B1(new_n674_), .B2(new_n678_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n616_), .A2(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n680_), .A2(new_n582_), .A3(new_n265_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(KEYINPUT107), .B(KEYINPUT38), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n682_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n660_), .A2(new_n675_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n495_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n613_), .A2(new_n608_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n575_), .A2(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n688_), .A2(new_n633_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n686_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n265_), .ZN(new_n691_));
  OAI21_X1  g490(.A(G1gat), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n683_), .A2(new_n684_), .A3(new_n692_), .ZN(G1324gat));
  INV_X1    g492(.A(new_n462_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n680_), .A2(new_n583_), .A3(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G8gat), .B1(new_n690_), .B2(new_n462_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT108), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n696_), .A2(new_n697_), .A3(KEYINPUT39), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n698_), .B1(KEYINPUT39), .B2(new_n696_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n697_), .B1(new_n696_), .B2(KEYINPUT39), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n695_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT40), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  OAI211_X1 g502(.A(KEYINPUT40), .B(new_n695_), .C1(new_n699_), .C2(new_n700_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1325gat));
  NAND3_X1  g504(.A1(new_n680_), .A2(new_n311_), .A3(new_n493_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT109), .ZN(new_n707_));
  INV_X1    g506(.A(new_n690_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n311_), .B1(new_n708_), .B2(new_n493_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT41), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n709_), .A2(new_n710_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n707_), .A2(new_n711_), .A3(new_n712_), .ZN(G1326gat));
  INV_X1    g512(.A(new_n492_), .ZN(new_n714_));
  OAI21_X1  g513(.A(G22gat), .B1(new_n690_), .B2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT42), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n714_), .A2(G22gat), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT110), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n680_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n716_), .A2(new_n719_), .ZN(G1327gat));
  NAND2_X1  g519(.A1(new_n633_), .A2(new_n685_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT112), .Z(new_n722_));
  AND2_X1   g521(.A1(new_n616_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(G29gat), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n265_), .A2(new_n724_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT113), .Z(new_n726_));
  NAND2_X1  g525(.A1(new_n723_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n668_), .A2(new_n671_), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT71), .B1(new_n647_), .B2(new_n659_), .ZN(new_n729_));
  AOI211_X1 g528(.A(new_n661_), .B(new_n658_), .C1(new_n669_), .C2(new_n645_), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n728_), .A2(new_n729_), .A3(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n678_), .B1(new_n731_), .B2(new_n676_), .ZN(new_n732_));
  OAI21_X1  g531(.A(KEYINPUT43), .B1(new_n495_), .B2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n400_), .A2(new_n406_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n462_), .A2(new_n734_), .A3(new_n691_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n491_), .A2(new_n494_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n677_), .B1(new_n673_), .B2(KEYINPUT37), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n737_), .A2(new_n738_), .A3(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n733_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n633_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n688_), .A2(new_n742_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n741_), .A2(new_n743_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n744_), .A2(KEYINPUT44), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n741_), .A2(new_n743_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n746_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n741_), .A2(KEYINPUT111), .A3(KEYINPUT44), .A4(new_n743_), .ZN(new_n750_));
  AOI211_X1 g549(.A(new_n691_), .B(new_n745_), .C1(new_n749_), .C2(new_n750_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n727_), .B1(new_n751_), .B2(new_n724_), .ZN(G1328gat));
  INV_X1    g551(.A(G36gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n723_), .A2(new_n753_), .A3(new_n694_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT45), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n694_), .B1(new_n744_), .B2(KEYINPUT44), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n757_));
  OAI211_X1 g556(.A(KEYINPUT46), .B(new_n755_), .C1(new_n757_), .C2(new_n753_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT46), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n749_), .A2(new_n750_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n462_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n753_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n754_), .B(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n759_), .B1(new_n762_), .B2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n758_), .A2(new_n765_), .ZN(G1329gat));
  OAI211_X1 g565(.A(G43gat), .B(new_n493_), .C1(new_n744_), .C2(KEYINPUT44), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n767_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n768_));
  AOI21_X1  g567(.A(G43gat), .B1(new_n723_), .B2(new_n493_), .ZN(new_n769_));
  OAI21_X1  g568(.A(KEYINPUT47), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n767_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n769_), .B1(new_n771_), .B2(new_n760_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT47), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n770_), .A2(new_n774_), .ZN(G1330gat));
  AOI21_X1  g574(.A(G50gat), .B1(new_n723_), .B2(new_n492_), .ZN(new_n776_));
  INV_X1    g575(.A(G50gat), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n745_), .A2(new_n777_), .A3(new_n714_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n776_), .B1(new_n778_), .B2(new_n760_), .ZN(G1331gat));
  NOR3_X1   g578(.A1(new_n495_), .A2(new_n575_), .A3(new_n687_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n780_), .A2(new_n679_), .ZN(new_n781_));
  AOI21_X1  g580(.A(G57gat), .B1(new_n781_), .B2(new_n265_), .ZN(new_n782_));
  AND4_X1   g581(.A1(new_n742_), .A2(new_n686_), .A3(new_n576_), .A4(new_n615_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n265_), .A2(G57gat), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n782_), .B1(new_n783_), .B2(new_n784_), .ZN(G1332gat));
  INV_X1    g584(.A(G64gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n786_), .B1(new_n783_), .B2(new_n694_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(KEYINPUT114), .B(KEYINPUT48), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n787_), .B(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n781_), .A2(new_n786_), .A3(new_n694_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(G1333gat));
  INV_X1    g590(.A(G71gat), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n792_), .B1(new_n783_), .B2(new_n493_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(KEYINPUT115), .B(KEYINPUT49), .ZN(new_n794_));
  OR2_X1    g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n794_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n332_), .A2(G71gat), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(KEYINPUT116), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n781_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n795_), .A2(new_n796_), .A3(new_n799_), .ZN(G1334gat));
  INV_X1    g599(.A(G78gat), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n783_), .B2(new_n492_), .ZN(new_n802_));
  XOR2_X1   g601(.A(new_n802_), .B(KEYINPUT50), .Z(new_n803_));
  NAND3_X1  g602(.A1(new_n781_), .A2(new_n801_), .A3(new_n492_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(G1335gat));
  NAND2_X1  g604(.A1(new_n780_), .A2(new_n722_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(G85gat), .B1(new_n807_), .B2(new_n265_), .ZN(new_n808_));
  NOR3_X1   g607(.A1(new_n575_), .A2(new_n742_), .A3(new_n687_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n741_), .A2(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n691_), .A2(new_n524_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n808_), .B1(new_n810_), .B2(new_n811_), .ZN(G1336gat));
  AOI21_X1  g611(.A(G92gat), .B1(new_n807_), .B2(new_n694_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n462_), .A2(new_n522_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n813_), .B1(new_n810_), .B2(new_n814_), .ZN(G1337gat));
  NAND3_X1  g614(.A1(new_n807_), .A2(new_n549_), .A3(new_n493_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n810_), .A2(new_n493_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n816_), .B1(new_n817_), .B2(new_n516_), .ZN(new_n818_));
  AND2_X1   g617(.A1(KEYINPUT117), .A2(KEYINPUT51), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n818_), .B(new_n819_), .ZN(G1338gat));
  NOR3_X1   g619(.A1(new_n806_), .A2(G106gat), .A3(new_n714_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT118), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n821_), .B(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n738_), .B1(new_n737_), .B2(new_n739_), .ZN(new_n825_));
  AOI211_X1 g624(.A(KEYINPUT43), .B(new_n732_), .C1(new_n735_), .C2(new_n736_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n492_), .B(new_n809_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT119), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n741_), .A2(KEYINPUT119), .A3(new_n492_), .A4(new_n809_), .ZN(new_n830_));
  AND4_X1   g629(.A1(new_n824_), .A2(new_n829_), .A3(G106gat), .A4(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n517_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n824_), .B1(new_n832_), .B2(new_n830_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n823_), .B1(new_n831_), .B2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(KEYINPUT53), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n823_), .B(new_n836_), .C1(new_n831_), .C2(new_n833_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n837_), .ZN(G1339gat));
  NAND3_X1  g637(.A1(new_n615_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n839_));
  NOR4_X1   g638(.A1(new_n739_), .A2(new_n839_), .A3(KEYINPUT54), .A4(new_n633_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n841_));
  INV_X1    g640(.A(new_n839_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n841_), .B1(new_n679_), .B2(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n840_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n560_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n556_), .A2(new_n497_), .A3(new_n559_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT120), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n846_), .A2(new_n847_), .A3(KEYINPUT55), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n847_), .B1(new_n846_), .B2(KEYINPUT55), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n845_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n846_), .A2(KEYINPUT55), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(KEYINPUT120), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n846_), .A2(new_n847_), .A3(KEYINPUT55), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(new_n560_), .A3(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n850_), .A2(new_n854_), .A3(new_n567_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(KEYINPUT56), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT56), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n850_), .A2(new_n854_), .A3(new_n857_), .A4(new_n567_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n856_), .A2(new_n569_), .A3(new_n687_), .A4(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n601_), .A2(new_n602_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n580_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n579_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n606_), .A2(new_n597_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n580_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n862_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n611_), .B1(new_n861_), .B2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n571_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n859_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n685_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n856_), .A2(new_n569_), .A3(new_n866_), .A4(new_n858_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT58), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n858_), .A2(new_n569_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n876_), .A2(KEYINPUT58), .A3(new_n866_), .A4(new_n856_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n875_), .A2(new_n877_), .A3(new_n739_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n868_), .A2(KEYINPUT57), .A3(new_n869_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n872_), .A2(new_n878_), .A3(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n844_), .B1(new_n880_), .B2(new_n633_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n691_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n694_), .A2(new_n406_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(G113gat), .B1(new_n884_), .B2(new_n687_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n880_), .A2(new_n633_), .ZN(new_n886_));
  OR2_X1    g685(.A1(new_n840_), .A2(new_n843_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n888_), .A2(KEYINPUT121), .A3(new_n265_), .A4(new_n883_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT59), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n882_), .A2(KEYINPUT121), .A3(KEYINPUT59), .A4(new_n883_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(G113gat), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n615_), .A2(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n885_), .B1(new_n893_), .B2(new_n895_), .ZN(G1340gat));
  AOI21_X1  g695(.A(new_n575_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n897_));
  INV_X1    g696(.A(G120gat), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(KEYINPUT60), .ZN(new_n899_));
  OR2_X1    g698(.A1(new_n575_), .A2(KEYINPUT60), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(new_n898_), .ZN(new_n901_));
  AOI21_X1  g700(.A(KEYINPUT122), .B1(new_n884_), .B2(new_n901_), .ZN(new_n902_));
  AND4_X1   g701(.A1(KEYINPUT122), .A2(new_n882_), .A3(new_n883_), .A4(new_n901_), .ZN(new_n903_));
  OAI22_X1  g702(.A1(new_n897_), .A2(new_n898_), .B1(new_n902_), .B2(new_n903_), .ZN(G1341gat));
  AOI21_X1  g703(.A(G127gat), .B1(new_n884_), .B2(new_n742_), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n742_), .A2(G127gat), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n905_), .B1(new_n893_), .B2(new_n906_), .ZN(G1342gat));
  AOI21_X1  g706(.A(G134gat), .B1(new_n884_), .B2(new_n685_), .ZN(new_n908_));
  AND2_X1   g707(.A1(new_n739_), .A2(G134gat), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n908_), .B1(new_n893_), .B2(new_n909_), .ZN(G1343gat));
  NOR2_X1   g709(.A1(new_n694_), .A2(new_n400_), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n882_), .A2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n687_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(G141gat), .ZN(new_n914_));
  INV_X1    g713(.A(G141gat), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n912_), .A2(new_n915_), .A3(new_n687_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n916_), .ZN(G1344gat));
  AND3_X1   g716(.A1(new_n882_), .A2(new_n576_), .A3(new_n911_), .ZN(new_n918_));
  XOR2_X1   g717(.A(new_n918_), .B(G148gat), .Z(G1345gat));
  NAND3_X1  g718(.A1(new_n882_), .A2(new_n742_), .A3(new_n911_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(KEYINPUT61), .B(G155gat), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n920_), .B(new_n921_), .ZN(G1346gat));
  AOI21_X1  g721(.A(G162gat), .B1(new_n912_), .B2(new_n685_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n732_), .A2(new_n649_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n923_), .B1(new_n912_), .B2(new_n924_), .ZN(G1347gat));
  NOR2_X1   g724(.A1(new_n881_), .A2(new_n492_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n694_), .A2(new_n691_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n927_), .A2(new_n332_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n926_), .A2(new_n687_), .A3(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n930_));
  AND3_X1   g729(.A1(new_n929_), .A2(new_n930_), .A3(G169gat), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n929_), .B2(G169gat), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n926_), .A2(new_n928_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n687_), .A2(new_n301_), .ZN(new_n934_));
  XOR2_X1   g733(.A(new_n934_), .B(KEYINPUT123), .Z(new_n935_));
  OAI22_X1  g734(.A1(new_n931_), .A2(new_n932_), .B1(new_n933_), .B2(new_n935_), .ZN(G1348gat));
  INV_X1    g735(.A(new_n933_), .ZN(new_n937_));
  AOI21_X1  g736(.A(G176gat), .B1(new_n937_), .B2(new_n576_), .ZN(new_n938_));
  OR3_X1    g737(.A1(new_n881_), .A2(KEYINPUT124), .A3(new_n492_), .ZN(new_n939_));
  OAI21_X1  g738(.A(KEYINPUT124), .B1(new_n881_), .B2(new_n492_), .ZN(new_n940_));
  AND3_X1   g739(.A1(new_n939_), .A2(new_n928_), .A3(new_n940_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n575_), .A2(new_n280_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n938_), .B1(new_n941_), .B2(new_n942_), .ZN(G1349gat));
  AND4_X1   g742(.A1(new_n742_), .A2(new_n926_), .A3(new_n414_), .A4(new_n928_), .ZN(new_n944_));
  NAND4_X1  g743(.A1(new_n939_), .A2(new_n742_), .A3(new_n928_), .A4(new_n940_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n944_), .B1(new_n945_), .B2(new_n275_), .ZN(G1350gat));
  OAI21_X1  g745(.A(G190gat), .B1(new_n933_), .B2(new_n732_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n685_), .A2(new_n277_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n933_), .B2(new_n948_), .ZN(G1351gat));
  NOR2_X1   g748(.A1(new_n927_), .A2(new_n400_), .ZN(new_n950_));
  INV_X1    g749(.A(new_n950_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n881_), .A2(new_n951_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n952_), .A2(new_n687_), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n953_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g753(.A1(new_n952_), .A2(new_n576_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n955_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g755(.A(new_n633_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n957_));
  AOI21_X1  g756(.A(KEYINPUT57), .B1(new_n868_), .B2(new_n869_), .ZN(new_n958_));
  AOI211_X1 g757(.A(new_n871_), .B(new_n685_), .C1(new_n859_), .C2(new_n867_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n958_), .A2(new_n959_), .ZN(new_n960_));
  AOI21_X1  g759(.A(new_n742_), .B1(new_n960_), .B2(new_n878_), .ZN(new_n961_));
  OAI211_X1 g760(.A(new_n950_), .B(new_n957_), .C1(new_n961_), .C2(new_n844_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n963_));
  XOR2_X1   g762(.A(new_n963_), .B(KEYINPUT125), .Z(new_n964_));
  INV_X1    g763(.A(new_n964_), .ZN(new_n965_));
  AOI21_X1  g764(.A(KEYINPUT126), .B1(new_n962_), .B2(new_n965_), .ZN(new_n966_));
  INV_X1    g765(.A(KEYINPUT127), .ZN(new_n967_));
  INV_X1    g766(.A(new_n957_), .ZN(new_n968_));
  NOR3_X1   g767(.A1(new_n881_), .A2(new_n951_), .A3(new_n968_), .ZN(new_n969_));
  AOI21_X1  g768(.A(new_n967_), .B1(new_n969_), .B2(new_n964_), .ZN(new_n970_));
  NOR3_X1   g769(.A1(new_n962_), .A2(KEYINPUT127), .A3(new_n965_), .ZN(new_n971_));
  OAI21_X1  g770(.A(new_n966_), .B1(new_n970_), .B2(new_n971_), .ZN(new_n972_));
  OAI21_X1  g771(.A(KEYINPUT127), .B1(new_n962_), .B2(new_n965_), .ZN(new_n973_));
  NAND4_X1  g772(.A1(new_n952_), .A2(new_n967_), .A3(new_n957_), .A4(new_n964_), .ZN(new_n974_));
  AOI21_X1  g773(.A(new_n964_), .B1(new_n952_), .B2(new_n957_), .ZN(new_n975_));
  OAI211_X1 g774(.A(new_n973_), .B(new_n974_), .C1(new_n975_), .C2(KEYINPUT126), .ZN(new_n976_));
  AND2_X1   g775(.A1(new_n972_), .A2(new_n976_), .ZN(G1354gat));
  AOI21_X1  g776(.A(G218gat), .B1(new_n952_), .B2(new_n685_), .ZN(new_n978_));
  AND2_X1   g777(.A1(new_n739_), .A2(G218gat), .ZN(new_n979_));
  AOI21_X1  g778(.A(new_n978_), .B1(new_n952_), .B2(new_n979_), .ZN(G1355gat));
endmodule


