//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 0 1 0 1 0 1 0 0 1 1 1 0 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n785_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n911_, new_n912_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_, new_n939_, new_n941_,
    new_n942_, new_n943_, new_n945_, new_n946_, new_n948_, new_n949_,
    new_n951_, new_n953_, new_n954_, new_n955_, new_n956_, new_n958_,
    new_n959_, new_n960_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(new_n202_), .A2(KEYINPUT73), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(KEYINPUT73), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G43gat), .B(G50gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n203_), .A2(new_n204_), .A3(new_n206_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT15), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G15gat), .B(G22gat), .ZN(new_n213_));
  INV_X1    g012(.A(G1gat), .ZN(new_n214_));
  INV_X1    g013(.A(G8gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT14), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G1gat), .B(G8gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n212_), .A2(new_n219_), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n210_), .A2(new_n219_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G229gat), .A2(G233gat), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n210_), .B(new_n219_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n222_), .ZN(new_n225_));
  AOI22_X1  g024(.A1(new_n220_), .A2(new_n223_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(G113gat), .B(G141gat), .Z(new_n227_));
  XNOR2_X1  g026(.A(G169gat), .B(G197gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n226_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n226_), .A2(new_n229_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(new_n232_), .B(KEYINPUT81), .Z(new_n233_));
  INV_X1    g032(.A(G169gat), .ZN(new_n234_));
  INV_X1    g033(.A(G176gat), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT24), .ZN(new_n237_));
  NOR2_X1   g036(.A1(G169gat), .A2(G176gat), .ZN(new_n238_));
  NOR3_X1   g037(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n239_), .A2(KEYINPUT82), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G183gat), .A2(G190gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT83), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT83), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n243_), .A2(G183gat), .A3(G190gat), .ZN(new_n244_));
  AOI21_X1  g043(.A(KEYINPUT23), .B1(new_n242_), .B2(new_n244_), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n241_), .A2(KEYINPUT23), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n239_), .A2(KEYINPUT82), .ZN(new_n248_));
  NOR3_X1   g047(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT25), .B(G183gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT26), .B(G190gat), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n249_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n240_), .A2(new_n247_), .A3(new_n248_), .A4(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT85), .B(KEYINPUT22), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT86), .B1(new_n254_), .B2(new_n234_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT86), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT22), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n257_), .A2(KEYINPUT85), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(KEYINPUT85), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n256_), .B(G169gat), .C1(new_n258_), .C2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT22), .B1(KEYINPUT84), .B2(G169gat), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(KEYINPUT84), .A2(G169gat), .ZN(new_n263_));
  AOI21_X1  g062(.A(G176gat), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n255_), .A2(new_n260_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n236_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(KEYINPUT87), .A3(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n242_), .A2(new_n244_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n268_), .B1(new_n269_), .B2(KEYINPUT23), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n270_), .B1(G183gat), .B2(G190gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n267_), .A2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(KEYINPUT87), .B1(new_n265_), .B2(new_n266_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n253_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G71gat), .B(G99gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(G43gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n274_), .B(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(G127gat), .B(G134gat), .Z(new_n278_));
  XOR2_X1   g077(.A(G113gat), .B(G120gat), .Z(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n277_), .B(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G227gat), .A2(G233gat), .ZN(new_n282_));
  INV_X1    g081(.A(G15gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT30), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT31), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n281_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n281_), .A2(new_n287_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G22gat), .B(G50gat), .ZN(new_n291_));
  XOR2_X1   g090(.A(new_n291_), .B(KEYINPUT92), .Z(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT28), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT3), .ZN(new_n295_));
  INV_X1    g094(.A(G141gat), .ZN(new_n296_));
  INV_X1    g095(.A(G148gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n295_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(KEYINPUT90), .B1(G141gat), .B2(G148gat), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT2), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n302_), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n300_), .A2(KEYINPUT91), .A3(new_n303_), .A4(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT88), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(KEYINPUT88), .A2(G155gat), .A3(G162gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n300_), .A2(new_n304_), .A3(new_n303_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT91), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n313_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT1), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n317_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT89), .B1(new_n318_), .B2(new_n311_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n308_), .A2(new_n317_), .A3(new_n309_), .ZN(new_n320_));
  AND3_X1   g119(.A1(KEYINPUT88), .A2(G155gat), .A3(G162gat), .ZN(new_n321_));
  AOI21_X1  g120(.A(KEYINPUT88), .B1(G155gat), .B2(G162gat), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT1), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT89), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n324_), .A3(new_n312_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n319_), .A2(new_n320_), .A3(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(G141gat), .B(G148gat), .Z(new_n327_));
  AOI22_X1  g126(.A1(new_n305_), .A2(new_n316_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT29), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n294_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n325_), .A2(new_n320_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n324_), .B1(new_n323_), .B2(new_n312_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n327_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n298_), .B(new_n299_), .C1(new_n302_), .C2(new_n301_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n304_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n315_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n336_), .A2(new_n305_), .A3(new_n312_), .A4(new_n310_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n333_), .A2(new_n337_), .A3(new_n329_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n338_), .A2(KEYINPUT28), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n293_), .B1(new_n330_), .B2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n328_), .A2(new_n294_), .A3(new_n329_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n338_), .A2(KEYINPUT28), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n341_), .A2(new_n342_), .A3(new_n292_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n340_), .A2(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n329_), .B1(new_n333_), .B2(new_n337_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G211gat), .B(G218gat), .ZN(new_n346_));
  AND2_X1   g145(.A1(G197gat), .A2(G204gat), .ZN(new_n347_));
  NOR2_X1   g146(.A1(G197gat), .A2(G204gat), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n346_), .B1(new_n349_), .B2(KEYINPUT93), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n350_), .A2(KEYINPUT21), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT21), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n347_), .A2(new_n348_), .ZN(new_n353_));
  XOR2_X1   g152(.A(G211gat), .B(G218gat), .Z(new_n354_));
  AOI21_X1  g153(.A(new_n352_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n351_), .B1(new_n350_), .B2(new_n355_), .ZN(new_n356_));
  OAI211_X1 g155(.A(G228gat), .B(G233gat), .C1(new_n345_), .C2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G228gat), .A2(G233gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n355_), .A2(new_n350_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n359_), .B1(KEYINPUT21), .B2(new_n350_), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n358_), .B(new_n360_), .C1(new_n328_), .C2(new_n329_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G78gat), .B(G106gat), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  AND3_X1   g162(.A1(new_n357_), .A2(new_n361_), .A3(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n363_), .B1(new_n357_), .B2(new_n361_), .ZN(new_n365_));
  NOR4_X1   g164(.A1(new_n344_), .A2(new_n364_), .A3(new_n365_), .A4(KEYINPUT94), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n340_), .A2(new_n343_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n357_), .A2(new_n361_), .A3(new_n363_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT94), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n357_), .A2(new_n361_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n362_), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n367_), .A2(new_n369_), .B1(new_n371_), .B2(new_n368_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n366_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT99), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n333_), .A2(new_n280_), .A3(new_n337_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n280_), .B1(new_n333_), .B2(new_n337_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT4), .ZN(new_n378_));
  NOR3_X1   g177(.A1(new_n376_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n333_), .A2(new_n337_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n280_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n380_), .A2(new_n378_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G225gat), .A2(G233gat), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n375_), .B1(new_n379_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n380_), .A2(new_n381_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n333_), .A2(new_n337_), .A3(new_n280_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n387_), .A2(KEYINPUT4), .A3(new_n388_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n389_), .A2(KEYINPUT99), .A3(new_n384_), .A4(new_n382_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G57gat), .B(G85gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT101), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(G1gat), .ZN(new_n393_));
  XOR2_X1   g192(.A(KEYINPUT100), .B(KEYINPUT0), .Z(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(G29gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n393_), .B(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n387_), .A2(new_n388_), .A3(new_n383_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n386_), .A2(new_n390_), .A3(new_n397_), .A4(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT33), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n253_), .B(new_n356_), .C1(new_n272_), .C2(new_n273_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT20), .ZN(new_n403_));
  OAI22_X1  g202(.A1(new_n245_), .A2(new_n246_), .B1(G183gat), .B2(G190gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n234_), .A2(KEYINPUT22), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n257_), .A2(G169gat), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(new_n406_), .A3(new_n235_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n266_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT96), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n407_), .A2(KEYINPUT96), .A3(new_n266_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n404_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT95), .ZN(new_n413_));
  INV_X1    g212(.A(G190gat), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n414_), .A2(KEYINPUT26), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n414_), .A2(KEYINPUT26), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n413_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n251_), .A2(KEYINPUT95), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n417_), .A2(new_n418_), .A3(new_n250_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n239_), .A2(new_n249_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(new_n420_), .A3(new_n270_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n412_), .A2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n403_), .B1(new_n422_), .B2(new_n360_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n402_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G226gat), .A2(G233gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT19), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT98), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n428_), .B(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G8gat), .B(G36gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G64gat), .B(G92gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n274_), .A2(new_n360_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n426_), .A2(new_n403_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n436_), .B1(new_n422_), .B2(new_n360_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n435_), .A2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n427_), .A2(new_n434_), .A3(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n434_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n426_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n442_), .B1(new_n402_), .B2(new_n423_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n437_), .B1(new_n274_), .B2(new_n360_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n441_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n387_), .A2(new_n388_), .A3(new_n384_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n382_), .A2(new_n383_), .ZN(new_n447_));
  OAI211_X1 g246(.A(new_n396_), .B(new_n446_), .C1(new_n379_), .C2(new_n447_), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n440_), .A2(new_n445_), .A3(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n396_), .A2(new_n400_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n386_), .A2(new_n390_), .A3(new_n398_), .A4(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n401_), .A2(new_n449_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT102), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n386_), .A2(new_n390_), .A3(new_n398_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n396_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n399_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n434_), .A2(KEYINPUT32), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n427_), .A2(new_n457_), .A3(new_n439_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT103), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n360_), .B1(new_n422_), .B2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n412_), .A2(new_n421_), .A3(KEYINPUT103), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n403_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n442_), .B1(new_n462_), .B2(new_n435_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n424_), .A2(new_n426_), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n457_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n458_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n452_), .A2(new_n453_), .B1(new_n456_), .B2(new_n467_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n401_), .A2(new_n449_), .A3(KEYINPUT102), .A4(new_n451_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n374_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n440_), .A2(new_n445_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT105), .B(KEYINPUT27), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  OR2_X1    g273(.A1(new_n434_), .A2(KEYINPUT104), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n434_), .A2(KEYINPUT104), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n475_), .B(new_n476_), .C1(new_n463_), .C2(new_n464_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT27), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n443_), .A2(new_n444_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n478_), .B1(new_n479_), .B2(new_n434_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n474_), .B(new_n481_), .C1(new_n366_), .C2(new_n372_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n482_), .A2(new_n456_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n290_), .B1(new_n470_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n290_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n456_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n481_), .A2(new_n474_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n485_), .A2(new_n373_), .A3(new_n486_), .A4(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n233_), .B1(new_n484_), .B2(new_n489_), .ZN(new_n490_));
  AND2_X1   g289(.A1(G231gat), .A2(G233gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n219_), .B(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G57gat), .B(G64gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G71gat), .B(G78gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(new_n494_), .A3(KEYINPUT11), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(KEYINPUT11), .ZN(new_n496_));
  INV_X1    g295(.A(new_n494_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n493_), .A2(KEYINPUT11), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n495_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT71), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n492_), .A2(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(G127gat), .B(G155gat), .Z(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G183gat), .B(G211gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT17), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n492_), .A2(new_n501_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n502_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT78), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n507_), .A2(new_n508_), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n500_), .B(KEYINPUT79), .Z(new_n515_));
  AOI211_X1 g314(.A(new_n509_), .B(new_n514_), .C1(new_n492_), .C2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n516_), .B1(new_n492_), .B2(new_n515_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n513_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT80), .ZN(new_n519_));
  AND2_X1   g318(.A1(G85gat), .A2(G92gat), .ZN(new_n520_));
  NOR2_X1   g319(.A1(G85gat), .A2(G92gat), .ZN(new_n521_));
  OAI21_X1  g320(.A(KEYINPUT67), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(G85gat), .ZN(new_n523_));
  INV_X1    g322(.A(G92gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT67), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G85gat), .A2(G92gat), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n525_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT8), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n522_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NOR3_X1   g331(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT66), .ZN(new_n535_));
  AND3_X1   g334(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n536_));
  AOI21_X1  g335(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n535_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G99gat), .A2(G106gat), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT6), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n541_), .A2(KEYINPUT66), .A3(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n534_), .A2(new_n538_), .A3(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n530_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT68), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n541_), .A2(KEYINPUT69), .A3(new_n542_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT69), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n549_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n534_), .A2(new_n548_), .A3(new_n550_), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n522_), .A2(new_n528_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT8), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n530_), .A2(new_n544_), .A3(KEYINPUT68), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n547_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(KEYINPUT10), .B(G99gat), .Z(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT64), .ZN(new_n558_));
  XNOR2_X1  g357(.A(KEYINPUT10), .B(G99gat), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT64), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(G106gat), .B1(new_n558_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n538_), .A2(new_n543_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT65), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT9), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n520_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT65), .B1(new_n525_), .B2(new_n527_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT9), .B1(new_n520_), .B2(new_n564_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n566_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NOR3_X1   g368(.A1(new_n562_), .A2(new_n563_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n556_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT70), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT70), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n556_), .A2(new_n571_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT71), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n500_), .B(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT12), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n573_), .A2(new_n575_), .A3(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G230gat), .A2(G233gat), .ZN(new_n581_));
  AOI21_X1  g380(.A(KEYINPUT68), .B1(new_n530_), .B2(new_n544_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n529_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n570_), .B1(new_n584_), .B2(new_n555_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n500_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n578_), .B1(new_n585_), .B2(new_n500_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n580_), .A2(new_n581_), .A3(new_n586_), .A4(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n586_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n585_), .A2(new_n500_), .ZN(new_n590_));
  OAI211_X1 g389(.A(G230gat), .B(G233gat), .C1(new_n589_), .C2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n588_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G120gat), .B(G148gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT5), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G176gat), .B(G204gat), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n594_), .B(new_n595_), .Z(new_n596_));
  NAND2_X1  g395(.A1(new_n592_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n596_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n588_), .A2(new_n591_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT13), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n597_), .B(new_n599_), .C1(KEYINPUT72), .C2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n602_));
  INV_X1    g401(.A(new_n599_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n598_), .B1(new_n588_), .B2(new_n591_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n602_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n601_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G190gat), .B(G218gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G134gat), .B(G162gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT36), .Z(new_n611_));
  NAND3_X1  g410(.A1(new_n573_), .A2(new_n212_), .A3(new_n575_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G232gat), .A2(G233gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT34), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT35), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n210_), .ZN(new_n619_));
  AOI22_X1  g418(.A1(new_n585_), .A2(new_n619_), .B1(new_n616_), .B2(new_n615_), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n612_), .A2(new_n618_), .A3(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n618_), .B1(new_n612_), .B2(new_n620_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n611_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n621_), .A2(new_n622_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n610_), .A2(KEYINPUT36), .ZN(new_n625_));
  AOI21_X1  g424(.A(KEYINPUT74), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n612_), .A2(new_n620_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n617_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n612_), .A2(new_n618_), .A3(new_n620_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n628_), .A2(KEYINPUT74), .A3(new_n629_), .A4(new_n625_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n623_), .B1(new_n626_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT76), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT75), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n623_), .A2(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n633_), .B1(new_n635_), .B2(KEYINPUT37), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT37), .ZN(new_n637_));
  AOI211_X1 g436(.A(KEYINPUT76), .B(new_n637_), .C1(new_n623_), .C2(new_n634_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n632_), .B1(new_n636_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n611_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n640_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n641_));
  OAI21_X1  g440(.A(KEYINPUT37), .B1(new_n641_), .B2(KEYINPUT75), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT76), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n628_), .A2(new_n629_), .A3(new_n625_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT74), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n641_), .B1(new_n646_), .B2(new_n630_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n635_), .A2(new_n633_), .A3(KEYINPUT37), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n643_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  AOI211_X1 g448(.A(new_n519_), .B(new_n607_), .C1(new_n639_), .C2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n490_), .A2(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT106), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n486_), .A2(KEYINPUT107), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n486_), .A2(KEYINPUT107), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n652_), .A2(new_n214_), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT38), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n647_), .B1(new_n484_), .B2(new_n489_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n232_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n607_), .A2(new_n660_), .A3(new_n518_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n659_), .A2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n214_), .B1(new_n662_), .B2(new_n456_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n658_), .A2(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n664_), .B1(new_n657_), .B2(new_n656_), .ZN(G1324gat));
  INV_X1    g464(.A(new_n662_), .ZN(new_n666_));
  OAI21_X1  g465(.A(G8gat), .B1(new_n666_), .B2(new_n488_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n667_), .A2(KEYINPUT39), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(KEYINPUT39), .ZN(new_n669_));
  INV_X1    g468(.A(new_n652_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n487_), .A2(new_n215_), .ZN(new_n671_));
  OAI22_X1  g470(.A1(new_n668_), .A2(new_n669_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(new_n675_));
  OAI221_X1 g474(.A(new_n673_), .B1(new_n670_), .B2(new_n671_), .C1(new_n668_), .C2(new_n669_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1325gat));
  AOI21_X1  g476(.A(new_n283_), .B1(new_n662_), .B2(new_n485_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT41), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n652_), .A2(new_n283_), .A3(new_n485_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1326gat));
  INV_X1    g480(.A(G22gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n662_), .B2(new_n374_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT42), .Z(new_n684_));
  NAND3_X1  g483(.A1(new_n652_), .A2(new_n682_), .A3(new_n374_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1327gat));
  NAND2_X1  g485(.A1(new_n519_), .A2(new_n647_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n687_), .A2(new_n607_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n490_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(G29gat), .B1(new_n690_), .B2(new_n456_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n519_), .A2(new_n232_), .A3(new_n606_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n639_), .A2(new_n649_), .ZN(new_n694_));
  AOI211_X1 g493(.A(KEYINPUT43), .B(new_n694_), .C1(new_n484_), .C2(new_n489_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT43), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n399_), .A2(new_n400_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n451_), .A2(new_n440_), .A3(new_n445_), .A4(new_n448_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n453_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n456_), .A2(new_n467_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(new_n469_), .A3(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n483_), .B1(new_n701_), .B2(new_n373_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n489_), .B1(new_n702_), .B2(new_n485_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n694_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n696_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  OAI211_X1 g504(.A(KEYINPUT44), .B(new_n693_), .C1(new_n695_), .C2(new_n705_), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n706_), .A2(G29gat), .A3(new_n655_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n693_), .B1(new_n695_), .B2(new_n705_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n691_), .B1(new_n707_), .B2(new_n710_), .ZN(G1328gat));
  INV_X1    g510(.A(new_n710_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n706_), .A2(new_n487_), .ZN(new_n713_));
  OAI21_X1  g512(.A(G36gat), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n488_), .A2(G36gat), .ZN(new_n716_));
  OR3_X1    g515(.A1(new_n689_), .A2(KEYINPUT45), .A3(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(KEYINPUT45), .B1(new_n689_), .B2(new_n716_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n715_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n714_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT110), .Z(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n720_), .B(new_n723_), .ZN(G1329gat));
  INV_X1    g523(.A(G43gat), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n725_), .B1(new_n689_), .B2(new_n290_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n290_), .A2(new_n725_), .ZN(new_n727_));
  AND4_X1   g526(.A1(KEYINPUT111), .A2(new_n710_), .A3(new_n706_), .A4(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n727_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n703_), .A2(new_n704_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT43), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n703_), .A2(new_n696_), .A3(new_n704_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n692_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n729_), .B1(new_n733_), .B2(KEYINPUT44), .ZN(new_n734_));
  AOI21_X1  g533(.A(KEYINPUT111), .B1(new_n734_), .B2(new_n710_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n726_), .B1(new_n728_), .B2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT47), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT47), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n738_), .B(new_n726_), .C1(new_n728_), .C2(new_n735_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(G1330gat));
  NAND2_X1  g539(.A1(new_n706_), .A2(new_n374_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G50gat), .B1(new_n712_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT112), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n742_), .B(new_n743_), .ZN(new_n744_));
  OR3_X1    g543(.A1(new_n689_), .A2(G50gat), .A3(new_n373_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1331gat));
  INV_X1    g545(.A(new_n233_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n747_), .A2(new_n606_), .A3(new_n519_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n659_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(G57gat), .B1(new_n750_), .B2(new_n486_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n232_), .B1(new_n484_), .B2(new_n489_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n519_), .ZN(new_n753_));
  AND4_X1   g552(.A1(new_n607_), .A2(new_n752_), .A3(new_n694_), .A4(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(G57gat), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n754_), .A2(new_n755_), .A3(new_n655_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n751_), .A2(new_n756_), .ZN(G1332gat));
  INV_X1    g556(.A(G64gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n749_), .B2(new_n487_), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT48), .Z(new_n760_));
  NAND3_X1  g559(.A1(new_n754_), .A2(new_n758_), .A3(new_n487_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(G1333gat));
  INV_X1    g561(.A(G71gat), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n763_), .B1(new_n749_), .B2(new_n485_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT49), .Z(new_n765_));
  NAND3_X1  g564(.A1(new_n754_), .A2(new_n763_), .A3(new_n485_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(G1334gat));
  INV_X1    g566(.A(G78gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n768_), .B1(new_n749_), .B2(new_n374_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT50), .Z(new_n770_));
  NAND3_X1  g569(.A1(new_n754_), .A2(new_n768_), .A3(new_n374_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(G1335gat));
  NOR2_X1   g571(.A1(new_n687_), .A2(new_n606_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n752_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n775_), .A2(new_n523_), .A3(new_n655_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n731_), .A2(new_n732_), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n753_), .A2(new_n232_), .A3(new_n606_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n456_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n776_), .B1(new_n781_), .B2(new_n523_), .ZN(G1336gat));
  NAND3_X1  g581(.A1(new_n775_), .A2(new_n524_), .A3(new_n487_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n779_), .A2(new_n487_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n783_), .B1(new_n785_), .B2(new_n524_), .ZN(G1337gat));
  AND2_X1   g585(.A1(new_n558_), .A2(new_n561_), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n774_), .A2(new_n290_), .A3(new_n787_), .ZN(new_n788_));
  XOR2_X1   g587(.A(new_n788_), .B(KEYINPUT113), .Z(new_n789_));
  NAND2_X1  g588(.A1(new_n779_), .A2(new_n485_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(G99gat), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n789_), .A2(new_n791_), .A3(new_n793_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(G1338gat));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n374_), .B(new_n778_), .C1(new_n695_), .C2(new_n705_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT116), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n799_), .A2(new_n800_), .A3(G106gat), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n799_), .B2(G106gat), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n798_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n799_), .A2(G106gat), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT116), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n799_), .A2(new_n800_), .A3(G106gat), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(KEYINPUT52), .A3(new_n806_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n774_), .A2(G106gat), .A3(new_n373_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT115), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n803_), .A2(new_n807_), .A3(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT53), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n803_), .A2(new_n807_), .A3(new_n812_), .A4(new_n809_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n813_), .ZN(G1339gat));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n694_), .A2(new_n233_), .A3(new_n606_), .A4(new_n753_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n815_), .B1(new_n816_), .B2(KEYINPUT54), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n650_), .A2(KEYINPUT117), .A3(new_n818_), .A4(new_n233_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n816_), .A2(KEYINPUT54), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n817_), .A2(new_n819_), .A3(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n660_), .A2(new_n603_), .ZN(new_n823_));
  XOR2_X1   g622(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n824_));
  NAND2_X1  g623(.A1(new_n588_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT119), .ZN(new_n826_));
  INV_X1    g625(.A(new_n575_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n574_), .B1(new_n556_), .B2(new_n571_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n501_), .A2(KEYINPUT12), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n827_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n587_), .A2(new_n586_), .ZN(new_n831_));
  OAI22_X1  g630(.A1(new_n830_), .A2(new_n831_), .B1(KEYINPUT120), .B2(new_n581_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n581_), .A2(KEYINPUT120), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n580_), .A2(new_n586_), .A3(new_n587_), .A4(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n581_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n832_), .A2(new_n834_), .A3(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT119), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n588_), .A2(new_n838_), .A3(new_n824_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n826_), .A2(new_n837_), .A3(new_n839_), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n840_), .A2(KEYINPUT56), .A3(new_n596_), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT56), .B1(new_n840_), .B2(new_n596_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n823_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n220_), .A2(new_n221_), .A3(new_n225_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n229_), .B1(new_n224_), .B2(new_n222_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n231_), .A2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n847_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n647_), .B1(new_n843_), .B2(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n822_), .B1(new_n850_), .B2(KEYINPUT121), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT121), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n840_), .A2(new_n596_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT56), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n840_), .A2(KEYINPUT56), .A3(new_n596_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n848_), .B1(new_n857_), .B2(new_n823_), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n852_), .B(KEYINPUT57), .C1(new_n858_), .C2(new_n647_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n603_), .A2(new_n847_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(KEYINPUT122), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n857_), .A2(KEYINPUT58), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n857_), .A2(new_n861_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT58), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n694_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  AOI22_X1  g664(.A1(new_n851_), .A2(new_n859_), .B1(new_n862_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n518_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n821_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n655_), .ZN(new_n869_));
  NOR4_X1   g668(.A1(new_n869_), .A2(new_n290_), .A3(new_n374_), .A4(new_n487_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(KEYINPUT59), .ZN(new_n872_));
  AND2_X1   g671(.A1(new_n870_), .A2(KEYINPUT123), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n870_), .A2(KEYINPUT123), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n873_), .A2(new_n874_), .A3(KEYINPUT59), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n851_), .A2(new_n859_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n865_), .A2(new_n862_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n753_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n817_), .A2(new_n819_), .A3(new_n820_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n875_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n821_), .B1(new_n866_), .B2(new_n753_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n883_), .A2(KEYINPUT124), .A3(new_n875_), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n872_), .A2(new_n882_), .A3(new_n747_), .A4(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(G113gat), .ZN(new_n886_));
  OR3_X1    g685(.A1(new_n871_), .A2(G113gat), .A3(new_n660_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1340gat));
  NAND4_X1  g687(.A1(new_n872_), .A2(new_n882_), .A3(new_n607_), .A4(new_n884_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(G120gat), .ZN(new_n890_));
  INV_X1    g689(.A(new_n871_), .ZN(new_n891_));
  INV_X1    g690(.A(G120gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n892_), .B1(new_n606_), .B2(KEYINPUT60), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n891_), .B(new_n893_), .C1(KEYINPUT60), .C2(new_n892_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n890_), .A2(new_n894_), .ZN(G1341gat));
  NAND4_X1  g694(.A1(new_n872_), .A2(new_n882_), .A3(new_n867_), .A4(new_n884_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(G127gat), .ZN(new_n897_));
  OR3_X1    g696(.A1(new_n871_), .A2(G127gat), .A3(new_n519_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1342gat));
  AOI21_X1  g698(.A(G134gat), .B1(new_n891_), .B2(new_n647_), .ZN(new_n900_));
  AND3_X1   g699(.A1(new_n872_), .A2(new_n882_), .A3(new_n884_), .ZN(new_n901_));
  XOR2_X1   g700(.A(KEYINPUT125), .B(G134gat), .Z(new_n902_));
  NOR2_X1   g701(.A1(new_n694_), .A2(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n900_), .B1(new_n901_), .B2(new_n903_), .ZN(G1343gat));
  AND2_X1   g703(.A1(new_n868_), .A2(new_n290_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n869_), .A2(new_n482_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  OAI21_X1  g706(.A(G141gat), .B1(new_n907_), .B2(new_n660_), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n905_), .A2(new_n296_), .A3(new_n232_), .A4(new_n906_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(G1344gat));
  OAI21_X1  g709(.A(G148gat), .B1(new_n907_), .B2(new_n606_), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n905_), .A2(new_n297_), .A3(new_n607_), .A4(new_n906_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1345gat));
  XNOR2_X1  g712(.A(KEYINPUT61), .B(G155gat), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n914_), .B1(new_n907_), .B2(new_n519_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n914_), .ZN(new_n916_));
  NAND4_X1  g715(.A1(new_n905_), .A2(new_n753_), .A3(new_n906_), .A4(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n915_), .A2(new_n917_), .ZN(G1346gat));
  INV_X1    g717(.A(new_n907_), .ZN(new_n919_));
  INV_X1    g718(.A(G162gat), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n694_), .A2(new_n920_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(KEYINPUT126), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n905_), .A2(new_n647_), .A3(new_n906_), .ZN(new_n923_));
  AOI22_X1  g722(.A1(new_n919_), .A2(new_n922_), .B1(new_n923_), .B2(new_n920_), .ZN(G1347gat));
  NOR2_X1   g723(.A1(new_n290_), .A2(new_n488_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n869_), .A2(new_n925_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n926_), .A2(new_n374_), .ZN(new_n927_));
  AND2_X1   g726(.A1(new_n883_), .A2(new_n927_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n232_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n929_));
  XOR2_X1   g728(.A(new_n929_), .B(KEYINPUT127), .Z(new_n930_));
  NAND2_X1  g729(.A1(new_n928_), .A2(new_n930_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n883_), .A2(new_n232_), .A3(new_n927_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT62), .ZN(new_n933_));
  AND3_X1   g732(.A1(new_n932_), .A2(new_n933_), .A3(G169gat), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n933_), .B1(new_n932_), .B2(G169gat), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n931_), .B1(new_n934_), .B2(new_n935_), .ZN(G1348gat));
  AOI21_X1  g735(.A(G176gat), .B1(new_n928_), .B2(new_n607_), .ZN(new_n937_));
  AND2_X1   g736(.A1(new_n868_), .A2(new_n373_), .ZN(new_n938_));
  NOR3_X1   g737(.A1(new_n926_), .A2(new_n235_), .A3(new_n606_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n937_), .B1(new_n938_), .B2(new_n939_), .ZN(G1349gat));
  NAND4_X1  g739(.A1(new_n938_), .A2(new_n753_), .A3(new_n869_), .A4(new_n925_), .ZN(new_n941_));
  INV_X1    g740(.A(G183gat), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n518_), .A2(new_n250_), .ZN(new_n943_));
  AOI22_X1  g742(.A1(new_n941_), .A2(new_n942_), .B1(new_n928_), .B2(new_n943_), .ZN(G1350gat));
  NAND4_X1  g743(.A1(new_n928_), .A2(new_n417_), .A3(new_n418_), .A4(new_n647_), .ZN(new_n945_));
  AND2_X1   g744(.A1(new_n928_), .A2(new_n704_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n945_), .B1(new_n946_), .B2(new_n414_), .ZN(G1351gat));
  NOR3_X1   g746(.A1(new_n488_), .A2(new_n373_), .A3(new_n456_), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n905_), .A2(new_n232_), .A3(new_n948_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n949_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g749(.A1(new_n905_), .A2(new_n607_), .A3(new_n948_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n951_), .B(G204gat), .ZN(G1353gat));
  NAND4_X1  g751(.A1(new_n868_), .A2(new_n290_), .A3(new_n867_), .A4(new_n948_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n954_));
  AND2_X1   g753(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n955_));
  NOR3_X1   g754(.A1(new_n953_), .A2(new_n954_), .A3(new_n955_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n956_), .B1(new_n953_), .B2(new_n954_), .ZN(G1354gat));
  NAND2_X1  g756(.A1(new_n905_), .A2(new_n948_), .ZN(new_n958_));
  OAI21_X1  g757(.A(G218gat), .B1(new_n958_), .B2(new_n694_), .ZN(new_n959_));
  OR2_X1    g758(.A1(new_n632_), .A2(G218gat), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n959_), .B1(new_n958_), .B2(new_n960_), .ZN(G1355gat));
endmodule


