//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 1 1 1 0 0 0 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n816_, new_n817_, new_n818_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n829_, new_n830_, new_n831_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n866_, new_n867_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_;
  OR2_X1    g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203_));
  NAND3_X1  g002(.A1(new_n202_), .A2(KEYINPUT24), .A3(new_n203_), .ZN(new_n204_));
  OAI21_X1  g003(.A(new_n204_), .B1(KEYINPUT24), .B2(new_n202_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n206_), .A2(G183gat), .A3(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT23), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n205_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT26), .B(G190gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT78), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT25), .B(G183gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT26), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n212_), .B1(new_n215_), .B2(G190gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n210_), .B1(new_n213_), .B2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT22), .B(G169gat), .ZN(new_n219_));
  INV_X1    g018(.A(G176gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(KEYINPUT79), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n209_), .B(KEYINPUT80), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n207_), .B(KEYINPUT81), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n223_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT82), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n222_), .B(new_n203_), .C1(new_n226_), .C2(new_n227_), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n226_), .A2(new_n227_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n218_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(G197gat), .A2(G204gat), .ZN(new_n231_));
  XOR2_X1   g030(.A(KEYINPUT85), .B(G197gat), .Z(new_n232_));
  AOI21_X1  g031(.A(new_n231_), .B1(new_n232_), .B2(G204gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G211gat), .B(G218gat), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n234_), .A2(KEYINPUT87), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT21), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n236_), .B1(new_n234_), .B2(KEYINPUT87), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n233_), .A2(new_n235_), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT88), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n233_), .A2(new_n235_), .A3(KEYINPUT88), .A4(new_n237_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n234_), .ZN(new_n243_));
  INV_X1    g042(.A(G204gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n232_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(G197gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n246_), .A2(KEYINPUT86), .A3(G204gat), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT86), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n248_), .B1(new_n244_), .B2(G197gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n245_), .A2(new_n247_), .A3(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n243_), .B1(new_n250_), .B2(KEYINPUT21), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n233_), .A2(KEYINPUT21), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n242_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n230_), .A2(new_n254_), .ZN(new_n255_));
  AND3_X1   g054(.A1(KEYINPUT19), .A2(G226gat), .A3(G233gat), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT19), .B1(G226gat), .B2(G233gat), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT20), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n240_), .A2(new_n241_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n205_), .B1(new_n211_), .B2(new_n214_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n224_), .A2(new_n225_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n209_), .A2(new_n207_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n264_), .B1(G183gat), .B2(G190gat), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n221_), .A2(new_n203_), .ZN(new_n266_));
  AOI22_X1  g065(.A1(new_n262_), .A2(new_n263_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n261_), .A2(new_n267_), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n268_), .A2(KEYINPUT90), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(KEYINPUT90), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n255_), .B(new_n260_), .C1(new_n269_), .C2(new_n270_), .ZN(new_n271_));
  XOR2_X1   g070(.A(new_n258_), .B(KEYINPUT89), .Z(new_n272_));
  NOR2_X1   g071(.A1(new_n230_), .A2(new_n254_), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT20), .B1(new_n261_), .B2(new_n267_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n272_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n271_), .A2(new_n275_), .ZN(new_n276_));
  XOR2_X1   g075(.A(G64gat), .B(G92gat), .Z(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT92), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G8gat), .B(G36gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n276_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n271_), .A2(new_n282_), .A3(new_n275_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  XOR2_X1   g085(.A(KEYINPUT98), .B(KEYINPUT27), .Z(new_n287_));
  AND2_X1   g086(.A1(new_n285_), .A2(KEYINPUT27), .ZN(new_n288_));
  OR3_X1    g087(.A1(new_n273_), .A2(new_n274_), .A3(new_n272_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n259_), .B1(new_n261_), .B2(new_n267_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(new_n255_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n291_), .A2(KEYINPUT96), .A3(new_n258_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(KEYINPUT96), .B1(new_n291_), .B2(new_n258_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n283_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  AOI22_X1  g094(.A1(new_n286_), .A2(new_n287_), .B1(new_n288_), .B2(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(G155gat), .B(G162gat), .Z(new_n297_));
  INV_X1    g096(.A(KEYINPUT1), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G141gat), .A2(G148gat), .ZN(new_n300_));
  INV_X1    g099(.A(G141gat), .ZN(new_n301_));
  INV_X1    g100(.A(G148gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n299_), .A2(new_n300_), .A3(new_n303_), .A4(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT84), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT3), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n306_), .A2(new_n307_), .A3(new_n301_), .A4(new_n302_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT2), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n300_), .A2(new_n309_), .ZN(new_n310_));
  OAI22_X1  g109(.A1(KEYINPUT84), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n308_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  OAI22_X1  g111(.A1(new_n300_), .A2(new_n309_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n297_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n305_), .A2(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n315_), .A2(KEYINPUT29), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n316_), .B(KEYINPUT28), .Z(new_n317_));
  AOI21_X1  g116(.A(new_n261_), .B1(KEYINPUT29), .B2(new_n315_), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n318_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G228gat), .A2(G233gat), .ZN(new_n321_));
  INV_X1    g120(.A(G78gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(G106gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G22gat), .B(G50gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n319_), .A2(new_n320_), .A3(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n327_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n296_), .A2(KEYINPUT99), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n288_), .A2(new_n295_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n285_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n282_), .B1(new_n271_), .B2(new_n275_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n287_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n332_), .A2(new_n330_), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT99), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n331_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT4), .ZN(new_n340_));
  INV_X1    g139(.A(new_n315_), .ZN(new_n341_));
  XOR2_X1   g140(.A(G127gat), .B(G134gat), .Z(new_n342_));
  XOR2_X1   g141(.A(G113gat), .B(G120gat), .Z(new_n343_));
  XOR2_X1   g142(.A(new_n342_), .B(new_n343_), .Z(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n340_), .B1(new_n341_), .B2(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(KEYINPUT93), .B1(new_n315_), .B2(new_n344_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n347_), .B1(new_n315_), .B2(new_n344_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n345_), .A2(KEYINPUT93), .A3(new_n305_), .A4(new_n314_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n346_), .B1(new_n350_), .B2(new_n340_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G225gat), .A2(G233gat), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n350_), .A2(new_n352_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(G1gat), .B(G29gat), .Z(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT94), .B(G85gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT0), .B(G57gat), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n359_), .B(new_n360_), .Z(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n356_), .A2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n354_), .A2(new_n361_), .A3(new_n355_), .ZN(new_n364_));
  AND3_X1   g163(.A1(new_n363_), .A2(KEYINPUT97), .A3(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(KEYINPUT97), .B1(new_n363_), .B2(new_n364_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n230_), .B(KEYINPUT30), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT83), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G71gat), .B(G99gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(G43gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G227gat), .A2(G233gat), .ZN(new_n373_));
  INV_X1    g172(.A(G15gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n372_), .B(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n370_), .A2(new_n377_), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n230_), .B(KEYINPUT30), .Z(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT83), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n376_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n344_), .B(KEYINPUT31), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n378_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n382_), .B1(new_n378_), .B2(new_n381_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n339_), .A2(new_n367_), .A3(new_n386_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n354_), .A2(KEYINPUT33), .A3(new_n361_), .A4(new_n355_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n351_), .A2(new_n352_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n361_), .B1(new_n350_), .B2(new_n353_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n284_), .A2(new_n388_), .A3(new_n391_), .A4(new_n285_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT33), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n364_), .A2(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n363_), .A2(new_n364_), .ZN(new_n396_));
  OAI211_X1 g195(.A(KEYINPUT32), .B(new_n282_), .C1(new_n293_), .C2(new_n294_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n282_), .A2(KEYINPUT32), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT95), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(new_n275_), .A3(new_n271_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n396_), .A2(new_n397_), .A3(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n330_), .B1(new_n395_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n330_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n296_), .A2(new_n367_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n385_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n387_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT70), .ZN(new_n409_));
  AND2_X1   g208(.A1(G230gat), .A2(G233gat), .ZN(new_n410_));
  OR2_X1    g209(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(new_n324_), .A3(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G99gat), .A2(G106gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT6), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT6), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n416_), .A2(G99gat), .A3(G106gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(G85gat), .ZN(new_n419_));
  INV_X1    g218(.A(G92gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G85gat), .A2(G92gat), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(KEYINPUT9), .A3(new_n422_), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n422_), .A2(KEYINPUT9), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n413_), .A2(new_n418_), .A3(new_n423_), .A4(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n421_), .A2(new_n422_), .ZN(new_n427_));
  INV_X1    g226(.A(G99gat), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT7), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n428_), .B(new_n324_), .C1(new_n429_), .C2(KEYINPUT64), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT64), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n431_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n429_), .A2(KEYINPUT64), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n430_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n415_), .A2(new_n417_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n427_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT8), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n418_), .A2(new_n432_), .A3(new_n430_), .A4(new_n433_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT8), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(new_n439_), .A3(new_n427_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n426_), .B1(new_n437_), .B2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G57gat), .B(G64gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G71gat), .B(G78gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n443_), .A3(KEYINPUT11), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(KEYINPUT11), .ZN(new_n445_));
  INV_X1    g244(.A(new_n443_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n442_), .A2(KEYINPUT11), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n444_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n410_), .B1(new_n441_), .B2(new_n449_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n438_), .A2(new_n439_), .A3(new_n427_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n439_), .B1(new_n438_), .B2(new_n427_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n425_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT12), .ZN(new_n454_));
  INV_X1    g253(.A(new_n449_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n453_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n454_), .B1(new_n453_), .B2(new_n455_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n450_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n425_), .B(new_n449_), .C1(new_n451_), .C2(new_n452_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT65), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n437_), .A2(new_n440_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT65), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n463_), .A2(new_n464_), .A3(new_n425_), .A4(new_n449_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n462_), .A2(KEYINPUT66), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n453_), .A2(new_n455_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(KEYINPUT66), .B1(new_n462_), .B2(new_n465_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n410_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT67), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  OAI211_X1 g271(.A(KEYINPUT67), .B(new_n410_), .C1(new_n468_), .C2(new_n469_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n460_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(G120gat), .B(G148gat), .Z(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT69), .ZN(new_n476_));
  XOR2_X1   g275(.A(G176gat), .B(G204gat), .Z(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n409_), .B1(new_n474_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n473_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT66), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n461_), .A2(KEYINPUT65), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n464_), .B1(new_n441_), .B2(new_n449_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n483_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n486_), .A2(new_n467_), .A3(new_n466_), .ZN(new_n487_));
  AOI21_X1  g286(.A(KEYINPUT67), .B1(new_n487_), .B2(new_n410_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n459_), .B1(new_n482_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n480_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(KEYINPUT70), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n481_), .A2(new_n491_), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n459_), .B(new_n480_), .C1(new_n482_), .C2(new_n488_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT71), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n474_), .A2(KEYINPUT71), .A3(new_n480_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n492_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT13), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n492_), .A2(new_n497_), .A3(KEYINPUT13), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G15gat), .B(G22gat), .ZN(new_n503_));
  INV_X1    g302(.A(G1gat), .ZN(new_n504_));
  INV_X1    g303(.A(G8gat), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT14), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n503_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G1gat), .B(G8gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(G29gat), .B(G36gat), .Z(new_n510_));
  XNOR2_X1  g309(.A(G43gat), .B(G50gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n509_), .B(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT76), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(G229gat), .A3(G233gat), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n512_), .B(KEYINPUT15), .Z(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n509_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G229gat), .A2(G233gat), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n509_), .A2(new_n512_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n515_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G113gat), .B(G141gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT77), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G169gat), .B(G197gat), .ZN(new_n524_));
  XOR2_X1   g323(.A(new_n523_), .B(new_n524_), .Z(new_n525_));
  OR2_X1    g324(.A1(new_n521_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n521_), .A2(new_n525_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n502_), .A2(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n408_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G232gat), .A2(G233gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT34), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n533_), .A2(KEYINPUT35), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n534_), .B1(new_n516_), .B2(new_n453_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n535_), .B1(new_n512_), .B2(new_n453_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n533_), .A2(KEYINPUT35), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT72), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n536_), .B(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G190gat), .B(G218gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G134gat), .B(G162gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n542_), .A2(KEYINPUT36), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(KEYINPUT36), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n539_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n539_), .A2(new_n543_), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT73), .B(KEYINPUT37), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n547_), .B(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G231gat), .A2(G233gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n509_), .B(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(new_n449_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT17), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT74), .ZN(new_n556_));
  NOR2_X1   g355(.A1(KEYINPUT75), .A2(KEYINPUT17), .ZN(new_n557_));
  AND2_X1   g356(.A1(KEYINPUT75), .A2(KEYINPUT17), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n555_), .B(new_n556_), .C1(new_n557_), .C2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G127gat), .B(G155gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT16), .ZN(new_n561_));
  XOR2_X1   g360(.A(G183gat), .B(G211gat), .Z(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT75), .ZN(new_n564_));
  OAI21_X1  g363(.A(KEYINPUT17), .B1(new_n556_), .B2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n563_), .B1(new_n554_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n559_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n555_), .A2(new_n563_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n551_), .A2(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n531_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n367_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n571_), .A2(new_n504_), .A3(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT38), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n408_), .A2(new_n547_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n569_), .B1(new_n575_), .B2(KEYINPUT100), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT100), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n408_), .A2(new_n577_), .A3(new_n547_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n576_), .A2(KEYINPUT101), .A3(new_n530_), .A4(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n385_), .B1(new_n331_), .B2(new_n338_), .ZN(new_n580_));
  AOI22_X1  g379(.A1(new_n580_), .A2(new_n367_), .B1(new_n406_), .B2(new_n385_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n547_), .ZN(new_n582_));
  OAI21_X1  g381(.A(KEYINPUT100), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n569_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n583_), .A2(new_n578_), .A3(new_n530_), .A4(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT101), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n367_), .B1(new_n579_), .B2(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n574_), .B1(new_n588_), .B2(new_n504_), .ZN(G1324gat));
  AOI21_X1  g388(.A(new_n505_), .B1(KEYINPUT102), .B2(KEYINPUT39), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n590_), .B1(new_n585_), .B2(new_n296_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(KEYINPUT102), .A2(KEYINPUT39), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  OAI221_X1 g392(.A(new_n590_), .B1(KEYINPUT102), .B2(KEYINPUT39), .C1(new_n585_), .C2(new_n296_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n296_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n571_), .A2(new_n505_), .A3(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n593_), .A2(new_n594_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT40), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(G1325gat));
  NAND3_X1  g398(.A1(new_n571_), .A2(new_n374_), .A3(new_n386_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n579_), .A2(new_n587_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(new_n386_), .ZN(new_n602_));
  AOI21_X1  g401(.A(KEYINPUT41), .B1(new_n602_), .B2(G15gat), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT41), .ZN(new_n604_));
  AOI211_X1 g403(.A(new_n604_), .B(new_n374_), .C1(new_n601_), .C2(new_n386_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n600_), .B1(new_n603_), .B2(new_n605_), .ZN(G1326gat));
  INV_X1    g405(.A(G22gat), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n571_), .A2(new_n607_), .A3(new_n404_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT42), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n601_), .A2(new_n404_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n609_), .B1(new_n610_), .B2(G22gat), .ZN(new_n611_));
  AOI211_X1 g410(.A(KEYINPUT42), .B(new_n607_), .C1(new_n601_), .C2(new_n404_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n608_), .B1(new_n611_), .B2(new_n612_), .ZN(G1327gat));
  NOR2_X1   g412(.A1(new_n547_), .A2(new_n584_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n531_), .A2(new_n614_), .ZN(new_n615_));
  OR3_X1    g414(.A1(new_n615_), .A2(G29gat), .A3(new_n367_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT43), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n617_), .B1(new_n581_), .B2(new_n550_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n408_), .A2(KEYINPUT43), .A3(new_n551_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n618_), .A2(new_n619_), .A3(new_n530_), .A4(new_n569_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT44), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  AOI211_X1 g421(.A(new_n572_), .B(new_n385_), .C1(new_n331_), .C2(new_n338_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n386_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n551_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n584_), .B1(new_n625_), .B2(new_n617_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n626_), .A2(KEYINPUT44), .A3(new_n530_), .A4(new_n619_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n622_), .A2(new_n627_), .A3(new_n572_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n628_), .A2(KEYINPUT103), .A3(G29gat), .ZN(new_n629_));
  AOI21_X1  g428(.A(KEYINPUT103), .B1(new_n628_), .B2(G29gat), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n616_), .B1(new_n629_), .B2(new_n630_), .ZN(G1328gat));
  NAND3_X1  g430(.A1(new_n622_), .A2(new_n627_), .A3(new_n595_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(G36gat), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n296_), .A2(G36gat), .ZN(new_n634_));
  OR3_X1    g433(.A1(new_n615_), .A2(KEYINPUT45), .A3(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(KEYINPUT45), .B1(new_n615_), .B2(new_n634_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n633_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT46), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n633_), .A2(KEYINPUT46), .A3(new_n637_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(G1329gat));
  NAND4_X1  g441(.A1(new_n622_), .A2(new_n627_), .A3(G43gat), .A4(new_n386_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n615_), .A2(new_n385_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n643_), .B1(G43gat), .B2(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g445(.A1(new_n622_), .A2(new_n627_), .A3(new_n404_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT104), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n647_), .A2(new_n648_), .A3(G50gat), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n647_), .B2(G50gat), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n330_), .A2(G50gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT105), .ZN(new_n652_));
  OAI22_X1  g451(.A1(new_n649_), .A2(new_n650_), .B1(new_n615_), .B2(new_n652_), .ZN(G1331gat));
  NAND2_X1  g452(.A1(new_n502_), .A2(new_n529_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n576_), .A2(new_n578_), .A3(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G57gat), .B1(new_n656_), .B2(new_n367_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n581_), .A2(new_n654_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n658_), .A2(new_n570_), .ZN(new_n659_));
  INV_X1    g458(.A(G57gat), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n659_), .A2(new_n660_), .A3(new_n572_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n657_), .A2(new_n661_), .ZN(G1332gat));
  INV_X1    g461(.A(G64gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n659_), .A2(new_n663_), .A3(new_n595_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n656_), .A2(new_n296_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT48), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n665_), .A2(new_n666_), .A3(G64gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n666_), .B1(new_n665_), .B2(G64gat), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n664_), .B1(new_n667_), .B2(new_n668_), .ZN(G1333gat));
  INV_X1    g468(.A(G71gat), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n659_), .A2(new_n670_), .A3(new_n386_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n576_), .A2(new_n386_), .A3(new_n578_), .A4(new_n655_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(G71gat), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT107), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT107), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n672_), .A2(new_n675_), .A3(G71gat), .ZN(new_n676_));
  XOR2_X1   g475(.A(KEYINPUT106), .B(KEYINPUT49), .Z(new_n677_));
  AND3_X1   g476(.A1(new_n674_), .A2(new_n676_), .A3(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n677_), .B1(new_n674_), .B2(new_n676_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n671_), .B1(new_n678_), .B2(new_n679_), .ZN(G1334gat));
  NAND3_X1  g479(.A1(new_n659_), .A2(new_n322_), .A3(new_n404_), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n656_), .A2(new_n330_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT50), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n682_), .A2(new_n683_), .A3(G78gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n682_), .B2(G78gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n681_), .B1(new_n684_), .B2(new_n685_), .ZN(G1335gat));
  NAND2_X1  g485(.A1(new_n658_), .A2(new_n614_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT108), .ZN(new_n688_));
  AOI21_X1  g487(.A(G85gat), .B1(new_n688_), .B2(new_n572_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n618_), .A2(new_n619_), .A3(new_n569_), .A4(new_n655_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT109), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n626_), .A2(KEYINPUT109), .A3(new_n619_), .A4(new_n655_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n367_), .A2(new_n419_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT110), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n690_), .A2(new_n698_), .A3(KEYINPUT111), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT111), .ZN(new_n700_));
  INV_X1    g499(.A(new_n698_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n700_), .B1(new_n701_), .B2(new_n689_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n699_), .A2(new_n702_), .ZN(G1336gat));
  NAND3_X1  g502(.A1(new_n688_), .A2(new_n420_), .A3(new_n595_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n296_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n704_), .B1(new_n420_), .B2(new_n705_), .ZN(G1337gat));
  AND2_X1   g505(.A1(new_n411_), .A2(new_n412_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n688_), .A2(new_n707_), .A3(new_n386_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n385_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n708_), .B1(new_n709_), .B2(new_n428_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT51), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT51), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n708_), .B(new_n712_), .C1(new_n709_), .C2(new_n428_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1338gat));
  NAND3_X1  g513(.A1(new_n688_), .A2(new_n324_), .A3(new_n404_), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n626_), .A2(new_n404_), .A3(new_n619_), .A4(new_n655_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT52), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n716_), .A2(new_n717_), .A3(G106gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n716_), .B2(G106gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n715_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n715_), .B(new_n721_), .C1(new_n718_), .C2(new_n719_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1339gat));
  AND2_X1   g524(.A1(new_n580_), .A2(new_n572_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n492_), .A2(new_n497_), .A3(KEYINPUT13), .ZN(new_n727_));
  AOI21_X1  g526(.A(KEYINPUT13), .B1(new_n492_), .B2(new_n497_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n569_), .A2(new_n528_), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT113), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n500_), .A2(KEYINPUT113), .A3(new_n501_), .A4(new_n730_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n550_), .ZN(new_n733_));
  OAI21_X1  g532(.A(KEYINPUT114), .B1(new_n731_), .B2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n500_), .A2(new_n501_), .A3(new_n730_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT113), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT114), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n737_), .A2(new_n738_), .A3(new_n550_), .A4(new_n732_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n734_), .A2(KEYINPUT54), .A3(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT54), .ZN(new_n741_));
  OAI211_X1 g540(.A(KEYINPUT114), .B(new_n741_), .C1(new_n731_), .C2(new_n733_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT117), .ZN(new_n744_));
  AOI22_X1  g543(.A1(new_n481_), .A2(new_n491_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n514_), .A2(new_n518_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n517_), .A2(new_n519_), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n746_), .B(new_n525_), .C1(new_n518_), .C2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n526_), .A2(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n744_), .B1(new_n745_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n749_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n498_), .A2(KEYINPUT117), .A3(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n497_), .A2(KEYINPUT115), .A3(new_n528_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n459_), .A2(KEYINPUT55), .ZN(new_n754_));
  INV_X1    g553(.A(new_n458_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n456_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT55), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(new_n757_), .A3(new_n450_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n754_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT116), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n457_), .A2(new_n458_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n462_), .A2(new_n465_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n410_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n759_), .A2(new_n760_), .A3(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n760_), .B1(new_n759_), .B2(new_n763_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n490_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT56), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n459_), .A2(KEYINPUT55), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n757_), .B1(new_n756_), .B2(new_n450_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n763_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT116), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n764_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(KEYINPUT56), .A3(new_n490_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n769_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n753_), .A2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT115), .B1(new_n497_), .B2(new_n528_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n750_), .B(new_n752_), .C1(new_n777_), .C2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n547_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT57), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT58), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT56), .B1(new_n774_), .B2(new_n490_), .ZN(new_n783_));
  AOI211_X1 g582(.A(new_n768_), .B(new_n480_), .C1(new_n773_), .C2(new_n764_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n751_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n497_), .ZN(new_n786_));
  OAI211_X1 g585(.A(KEYINPUT118), .B(new_n782_), .C1(new_n785_), .C2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(KEYINPUT118), .B1(new_n785_), .B2(new_n786_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n550_), .B1(new_n788_), .B2(KEYINPUT58), .ZN(new_n789_));
  AOI22_X1  g588(.A1(new_n780_), .A2(new_n781_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n779_), .A2(KEYINPUT57), .A3(new_n547_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n584_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n726_), .B1(new_n743_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(G113gat), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n794_), .A2(new_n795_), .A3(new_n528_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT59), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n793_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n780_), .A2(new_n781_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n789_), .A2(new_n787_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n799_), .A2(new_n791_), .A3(new_n800_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n742_), .B(new_n740_), .C1(new_n801_), .C2(new_n584_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n802_), .A2(KEYINPUT59), .A3(new_n726_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n529_), .B1(new_n798_), .B2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n796_), .B1(new_n804_), .B2(new_n795_), .ZN(G1340gat));
  AOI21_X1  g604(.A(new_n729_), .B1(new_n798_), .B2(new_n803_), .ZN(new_n806_));
  INV_X1    g605(.A(G120gat), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n807_), .B1(new_n729_), .B2(KEYINPUT60), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n808_), .B1(KEYINPUT60), .B2(new_n807_), .ZN(new_n809_));
  OAI22_X1  g608(.A1(new_n806_), .A2(new_n807_), .B1(new_n793_), .B2(new_n809_), .ZN(G1341gat));
  AOI21_X1  g609(.A(G127gat), .B1(new_n794_), .B2(new_n584_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n798_), .A2(new_n803_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n584_), .A2(G127gat), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT119), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n811_), .B1(new_n812_), .B2(new_n814_), .ZN(G1342gat));
  INV_X1    g614(.A(G134gat), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n794_), .A2(new_n816_), .A3(new_n582_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n550_), .B1(new_n798_), .B2(new_n803_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n817_), .B1(new_n818_), .B2(new_n816_), .ZN(G1343gat));
  NOR2_X1   g618(.A1(new_n743_), .A2(new_n792_), .ZN(new_n820_));
  NOR4_X1   g619(.A1(new_n386_), .A2(new_n595_), .A3(new_n367_), .A4(new_n330_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(KEYINPUT120), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n820_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n528_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(G141gat), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n824_), .A2(new_n301_), .A3(new_n528_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(G1344gat));
  XNOR2_X1  g627(.A(KEYINPUT121), .B(G148gat), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n824_), .A2(new_n502_), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n824_), .B2(new_n502_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(G1345gat));
  NAND2_X1  g631(.A1(new_n824_), .A2(new_n584_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(KEYINPUT61), .B(G155gat), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n834_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n824_), .A2(new_n584_), .A3(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n837_), .ZN(G1346gat));
  OAI211_X1 g637(.A(new_n551_), .B(new_n822_), .C1(new_n743_), .C2(new_n792_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(G162gat), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n547_), .A2(G162gat), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n802_), .A2(new_n822_), .A3(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(KEYINPUT122), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT122), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n840_), .A2(new_n845_), .A3(new_n842_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n844_), .A2(new_n846_), .ZN(G1347gat));
  NOR2_X1   g646(.A1(new_n820_), .A2(new_n404_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n572_), .A2(new_n385_), .A3(new_n296_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n848_), .A2(new_n528_), .A3(new_n219_), .A4(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n528_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(KEYINPUT123), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n802_), .A2(new_n330_), .A3(new_n852_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n854_));
  AND3_X1   g653(.A1(new_n853_), .A2(G169gat), .A3(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n853_), .B2(G169gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n850_), .B1(new_n855_), .B2(new_n856_), .ZN(G1348gat));
  NAND4_X1  g656(.A1(new_n802_), .A2(new_n502_), .A3(new_n330_), .A4(new_n849_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G176gat), .ZN(G1349gat));
  INV_X1    g658(.A(new_n214_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n848_), .A2(new_n860_), .A3(new_n584_), .A4(new_n849_), .ZN(new_n861_));
  INV_X1    g660(.A(G183gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n802_), .A2(new_n330_), .A3(new_n849_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n863_), .B2(new_n569_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n861_), .A2(new_n864_), .ZN(G1350gat));
  OAI21_X1  g664(.A(G190gat), .B1(new_n863_), .B2(new_n550_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n582_), .A2(new_n211_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n863_), .B2(new_n867_), .ZN(G1351gat));
  NAND3_X1  g667(.A1(new_n385_), .A2(new_n367_), .A3(new_n404_), .ZN(new_n869_));
  XOR2_X1   g668(.A(new_n869_), .B(KEYINPUT125), .Z(new_n870_));
  NOR2_X1   g669(.A1(new_n870_), .A2(new_n296_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n802_), .A2(G197gat), .A3(new_n528_), .A4(new_n871_), .ZN(new_n872_));
  AND2_X1   g671(.A1(new_n872_), .A2(KEYINPUT126), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n528_), .B(new_n871_), .C1(new_n743_), .C2(new_n792_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n246_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n875_), .B1(new_n872_), .B2(KEYINPUT126), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n873_), .A2(new_n876_), .ZN(G1352gat));
  AND2_X1   g676(.A1(new_n802_), .A2(new_n871_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n502_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(G204gat), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n878_), .A2(new_n244_), .A3(new_n502_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1353gat));
  NAND3_X1  g681(.A1(new_n802_), .A2(new_n584_), .A3(new_n871_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT63), .B(G211gat), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n885_), .B1(new_n883_), .B2(new_n886_), .ZN(G1354gat));
  NAND2_X1  g686(.A1(new_n878_), .A2(new_n582_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT127), .B(G218gat), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n550_), .A2(new_n889_), .ZN(new_n890_));
  AOI22_X1  g689(.A1(new_n888_), .A2(new_n889_), .B1(new_n878_), .B2(new_n890_), .ZN(G1355gat));
endmodule


