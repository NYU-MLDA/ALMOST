//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 0 0 1 0 1 0 1 0 1 1 1 1 1 1 1 1 1 1 1 1 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n611_,
    new_n612_, new_n613_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n854_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n863_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n892_, new_n894_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XOR2_X1   g002(.A(G1gat), .B(G8gat), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT71), .B(G15gat), .ZN(new_n206_));
  INV_X1    g005(.A(G22gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT72), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G1gat), .A2(G8gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT14), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n208_), .A2(new_n209_), .A3(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n209_), .B1(new_n208_), .B2(new_n211_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n205_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n214_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(new_n204_), .A3(new_n212_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G29gat), .B(G36gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT69), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G43gat), .B(G50gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n218_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n221_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n220_), .B(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n225_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n203_), .B1(new_n223_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n226_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT15), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n225_), .A2(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n222_), .A2(KEYINPUT15), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n217_), .B(new_n215_), .C1(new_n230_), .C2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n228_), .A2(new_n232_), .A3(new_n202_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G113gat), .B(G141gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G169gat), .B(G197gat), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n234_), .B(new_n235_), .Z(new_n236_));
  AND3_X1   g035(.A1(new_n227_), .A2(new_n233_), .A3(new_n236_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n236_), .B1(new_n227_), .B2(new_n233_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G183gat), .A2(G190gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT23), .ZN(new_n241_));
  NOR2_X1   g040(.A1(G169gat), .A2(G176gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT24), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT75), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT25), .B(G183gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT26), .B(G190gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n242_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G169gat), .A2(G176gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(KEYINPUT24), .A3(new_n251_), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n249_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT75), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n241_), .A2(new_n254_), .A3(new_n244_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n246_), .A2(new_n253_), .A3(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT76), .B(G176gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT22), .B(G169gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n259_), .A2(new_n251_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n241_), .B1(G183gat), .B2(G190gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n256_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT30), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT78), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n256_), .A2(KEYINPUT30), .A3(new_n262_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT31), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT31), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n265_), .A2(new_n266_), .A3(new_n270_), .A4(new_n267_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G71gat), .B(G99gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(G43gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT77), .B(G15gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G227gat), .A2(G233gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n266_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G127gat), .B(G134gat), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  XOR2_X1   g080(.A(G113gat), .B(G120gat), .Z(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G113gat), .B(G120gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n280_), .A2(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(KEYINPUT79), .B1(new_n283_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n283_), .A2(KEYINPUT79), .A3(new_n285_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NOR3_X1   g089(.A1(new_n278_), .A2(new_n279_), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n277_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n276_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n267_), .ZN(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT30), .B1(new_n256_), .B2(new_n262_), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT78), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n289_), .B1(new_n293_), .B2(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n272_), .B1(new_n291_), .B2(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n290_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n293_), .A2(new_n296_), .A3(new_n289_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n299_), .A2(new_n300_), .A3(new_n269_), .A4(new_n271_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G155gat), .A2(G162gat), .ZN(new_n304_));
  OR2_X1    g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305_));
  NOR3_X1   g104(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT81), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G141gat), .A2(G148gat), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT2), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT3), .ZN(new_n312_));
  NOR2_X1   g111(.A1(G141gat), .A2(G148gat), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n310_), .B(new_n311_), .C1(new_n312_), .C2(new_n313_), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n304_), .B(new_n305_), .C1(new_n307_), .C2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT29), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n304_), .A2(KEYINPUT1), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n304_), .A2(KEYINPUT1), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n317_), .A2(KEYINPUT80), .A3(new_n318_), .A4(new_n305_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n313_), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n320_), .A2(new_n308_), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n319_), .B(new_n321_), .C1(KEYINPUT80), .C2(new_n317_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n315_), .A2(new_n316_), .A3(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT28), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n315_), .A2(new_n322_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT29), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G211gat), .B(G218gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT83), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT21), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  XOR2_X1   g129(.A(G197gat), .B(G204gat), .Z(new_n331_));
  OAI211_X1 g130(.A(new_n330_), .B(new_n331_), .C1(KEYINPUT21), .C2(new_n328_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n331_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n333_), .B(KEYINPUT21), .C1(new_n329_), .C2(new_n328_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G78gat), .B(G106gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G228gat), .A2(G233gat), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n336_), .B(new_n337_), .Z(new_n338_));
  NAND3_X1  g137(.A1(new_n327_), .A2(new_n335_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT82), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n338_), .B1(new_n327_), .B2(new_n335_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n325_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G22gat), .B(G50gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n341_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n344_), .A2(new_n324_), .A3(KEYINPUT82), .A4(new_n339_), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n342_), .A2(new_n343_), .A3(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n343_), .B1(new_n342_), .B2(new_n345_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n303_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n289_), .A2(new_n326_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n283_), .A2(new_n285_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT86), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n283_), .A2(KEYINPUT86), .A3(new_n285_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n353_), .A2(new_n315_), .A3(new_n322_), .A4(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G225gat), .A2(G233gat), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n350_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  AND3_X1   g156(.A1(new_n350_), .A2(KEYINPUT4), .A3(new_n355_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT4), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n289_), .A2(new_n359_), .A3(new_n326_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n360_), .A2(G225gat), .A3(G233gat), .ZN(new_n361_));
  NOR3_X1   g160(.A1(new_n358_), .A2(new_n361_), .A3(KEYINPUT87), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT87), .ZN(new_n363_));
  INV_X1    g162(.A(new_n356_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n360_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n350_), .A2(KEYINPUT4), .A3(new_n355_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n363_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n357_), .B1(new_n362_), .B2(new_n367_), .ZN(new_n368_));
  XOR2_X1   g167(.A(G1gat), .B(G29gat), .Z(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT88), .B(KEYINPUT0), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G57gat), .B(G85gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n368_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n357_), .A2(new_n373_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT87), .B1(new_n358_), .B2(new_n361_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n365_), .A2(new_n366_), .A3(new_n363_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n376_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT92), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  AOI211_X1 g180(.A(KEYINPUT92), .B(new_n376_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n375_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G226gat), .A2(G233gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT19), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n249_), .A2(new_n252_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(KEYINPUT84), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n241_), .B(new_n244_), .C1(new_n386_), .C2(KEYINPUT84), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n262_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n335_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT20), .B1(new_n263_), .B2(new_n335_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n385_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n335_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n395_), .B(new_n262_), .C1(new_n388_), .C2(new_n389_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n385_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n263_), .A2(new_n335_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n396_), .A2(KEYINPUT20), .A3(new_n397_), .A4(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n394_), .A2(new_n399_), .ZN(new_n400_));
  XOR2_X1   g199(.A(G8gat), .B(G36gat), .Z(new_n401_));
  XNOR2_X1  g200(.A(G64gat), .B(G92gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT85), .B(KEYINPUT18), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT32), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n400_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT20), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n256_), .A2(new_n262_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n409_), .B1(new_n410_), .B2(new_n395_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(new_n397_), .A3(new_n391_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT91), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT91), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n411_), .A2(new_n414_), .A3(new_n397_), .A4(new_n391_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT90), .B(KEYINPUT20), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n396_), .A2(new_n398_), .A3(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n385_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n413_), .A2(new_n415_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n408_), .B1(new_n407_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n383_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n405_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n400_), .A2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n394_), .A2(new_n405_), .A3(new_n399_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n366_), .A2(new_n356_), .A3(new_n360_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n350_), .A2(new_n355_), .A3(new_n364_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n427_), .A2(new_n374_), .ZN(new_n428_));
  AOI22_X1  g227(.A1(new_n379_), .A2(KEYINPUT33), .B1(new_n426_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n376_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n430_), .B1(new_n362_), .B2(new_n367_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT33), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(KEYINPUT89), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT89), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n434_), .B1(new_n379_), .B2(KEYINPUT33), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n425_), .A2(new_n429_), .A3(new_n433_), .A4(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n349_), .B1(new_n421_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(KEYINPUT27), .B1(new_n423_), .B2(new_n424_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n424_), .A2(KEYINPUT27), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n405_), .B(KEYINPUT93), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  AOI22_X1  g241(.A1(new_n412_), .A2(KEYINPUT91), .B1(new_n417_), .B2(new_n385_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n442_), .B1(new_n443_), .B2(new_n415_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT94), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n440_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n419_), .A2(new_n441_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT94), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n439_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n342_), .A2(new_n345_), .A3(new_n343_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n347_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n302_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n301_), .B(new_n298_), .C1(new_n346_), .C2(new_n347_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n383_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n449_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n239_), .B1(new_n438_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT68), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G230gat), .A2(G233gat), .ZN(new_n459_));
  NOR2_X1   g258(.A1(G85gat), .A2(G92gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G85gat), .A2(G92gat), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT9), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n460_), .B1(new_n463_), .B2(KEYINPUT64), .ZN(new_n464_));
  NAND3_X1  g263(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT65), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT65), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n467_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT64), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n461_), .A2(new_n470_), .A3(new_n462_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n464_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n472_));
  AND2_X1   g271(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n473_));
  NOR2_X1   g272(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n474_));
  NOR3_X1   g273(.A1(new_n473_), .A2(new_n474_), .A3(G106gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G99gat), .A2(G106gat), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT6), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n475_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n472_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT7), .ZN(new_n483_));
  INV_X1    g282(.A(G99gat), .ZN(new_n484_));
  INV_X1    g283(.A(G106gat), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n483_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n486_), .A2(new_n478_), .A3(new_n479_), .A4(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT8), .ZN(new_n489_));
  XOR2_X1   g288(.A(G85gat), .B(G92gat), .Z(new_n490_));
  AND3_X1   g289(.A1(new_n488_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n489_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n482_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G57gat), .B(G64gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT11), .ZN(new_n495_));
  XOR2_X1   g294(.A(G71gat), .B(G78gat), .Z(new_n496_));
  NOR2_X1   g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n496_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n494_), .A2(KEYINPUT11), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n497_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT66), .B1(new_n493_), .B2(new_n502_), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n491_), .A2(new_n492_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n497_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n505_), .B1(new_n498_), .B2(new_n500_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n504_), .A2(new_n482_), .A3(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n459_), .B1(new_n503_), .B2(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n508_), .B1(new_n507_), .B2(new_n503_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT67), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT12), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n493_), .A2(new_n502_), .A3(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n510_), .A2(new_n511_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n493_), .A2(new_n502_), .A3(new_n514_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n516_), .A2(new_n459_), .A3(new_n507_), .A4(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G120gat), .B(G148gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT5), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G176gat), .B(G204gat), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n520_), .B(new_n521_), .Z(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n509_), .A2(new_n518_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n523_), .B1(new_n509_), .B2(new_n518_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n458_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n526_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n529_), .A2(KEYINPUT68), .A3(new_n524_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT13), .ZN(new_n532_));
  NOR3_X1   g331(.A1(new_n528_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(KEYINPUT13), .B1(new_n527_), .B2(new_n530_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n225_), .B(new_n229_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(new_n493_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n222_), .A2(new_n504_), .A3(new_n482_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G232gat), .A2(G233gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT34), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT70), .B1(new_n540_), .B2(KEYINPUT35), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n537_), .A2(new_n538_), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n540_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT35), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G190gat), .B(G218gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G134gat), .B(G162gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n550_), .A2(KEYINPUT36), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n541_), .B1(new_n536_), .B2(new_n493_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n546_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n552_), .A2(new_n553_), .A3(new_n538_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n547_), .A2(new_n551_), .A3(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n550_), .B(KEYINPUT36), .Z(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n557_), .B1(new_n547_), .B2(new_n554_), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT37), .B1(new_n555_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n554_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n553_), .B1(new_n552_), .B2(new_n538_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n556_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n547_), .A2(new_n551_), .A3(new_n554_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT37), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n562_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n559_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G231gat), .A2(G233gat), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n568_), .B(KEYINPUT73), .Z(new_n569_));
  NOR2_X1   g368(.A1(new_n218_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n569_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n571_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(new_n506_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n502_), .B1(new_n570_), .B2(new_n572_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(G127gat), .B(G155gat), .Z(new_n577_));
  XNOR2_X1  g376(.A(G183gat), .B(G211gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n581_), .A2(KEYINPUT17), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n576_), .A2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n581_), .A2(KEYINPUT17), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n574_), .A2(new_n575_), .A3(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n586_), .ZN(new_n587_));
  NOR3_X1   g386(.A1(new_n535_), .A2(new_n567_), .A3(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n457_), .A2(new_n588_), .ZN(new_n589_));
  NOR3_X1   g388(.A1(new_n589_), .A2(G1gat), .A3(new_n455_), .ZN(new_n590_));
  XOR2_X1   g389(.A(KEYINPUT95), .B(KEYINPUT38), .Z(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n555_), .A2(new_n558_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n593_), .B1(new_n438_), .B2(new_n456_), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n535_), .A2(new_n587_), .A3(new_n239_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(G1gat), .B1(new_n596_), .B2(new_n455_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n592_), .A2(new_n597_), .ZN(G1324gat));
  NOR3_X1   g397(.A1(new_n589_), .A2(G8gat), .A3(new_n449_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT96), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n600_), .B1(new_n596_), .B2(new_n449_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n449_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n594_), .A2(new_n595_), .A3(KEYINPUT96), .A4(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n601_), .A2(G8gat), .A3(new_n603_), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n604_), .A2(KEYINPUT39), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(KEYINPUT39), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n599_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(KEYINPUT97), .B(KEYINPUT40), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n607_), .B(new_n609_), .ZN(G1325gat));
  OAI21_X1  g409(.A(G15gat), .B1(new_n596_), .B2(new_n303_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT41), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n589_), .A2(G15gat), .A3(new_n303_), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n612_), .A2(new_n613_), .ZN(G1326gat));
  OAI21_X1  g413(.A(G22gat), .B1(new_n596_), .B2(new_n348_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT42), .ZN(new_n616_));
  INV_X1    g415(.A(new_n348_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(new_n207_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT98), .Z(new_n619_));
  OAI21_X1  g418(.A(new_n616_), .B1(new_n589_), .B2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT99), .ZN(G1327gat));
  AND2_X1   g420(.A1(new_n425_), .A2(new_n429_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n433_), .A2(new_n435_), .ZN(new_n623_));
  AOI22_X1  g422(.A1(new_n622_), .A2(new_n623_), .B1(new_n383_), .B2(new_n420_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n456_), .B1(new_n624_), .B2(new_n349_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n535_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n239_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n593_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n587_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n625_), .A2(new_n626_), .A3(new_n627_), .A4(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(KEYINPUT102), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT102), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n457_), .A2(new_n633_), .A3(new_n626_), .A4(new_n630_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(G29gat), .B1(new_n636_), .B2(new_n383_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT43), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n449_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n567_), .B(new_n638_), .C1(new_n639_), .C2(new_n437_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(KEYINPUT100), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n567_), .B1(new_n639_), .B2(new_n437_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT43), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n625_), .A2(new_n644_), .A3(new_n638_), .A4(new_n567_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n641_), .A2(new_n643_), .A3(new_n645_), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n535_), .A2(new_n629_), .A3(new_n239_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n646_), .A2(KEYINPUT44), .A3(new_n647_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n648_), .A2(G29gat), .A3(new_n383_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n647_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(KEYINPUT101), .B(KEYINPUT44), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n637_), .B1(new_n649_), .B2(new_n653_), .ZN(G1328gat));
  NOR2_X1   g453(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT106), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n449_), .A2(G36gat), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n632_), .A2(new_n634_), .A3(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n659_), .B(KEYINPUT104), .Z(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n658_), .A2(new_n661_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n632_), .A2(new_n634_), .A3(new_n657_), .A4(new_n660_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n646_), .A2(KEYINPUT44), .A3(new_n647_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n651_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n666_), .A2(new_n667_), .A3(new_n449_), .ZN(new_n668_));
  INV_X1    g467(.A(G36gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n665_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n656_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n653_), .A2(new_n602_), .A3(new_n648_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n664_), .B1(new_n673_), .B2(G36gat), .ZN(new_n674_));
  INV_X1    g473(.A(new_n671_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n656_), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n674_), .A2(new_n675_), .A3(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n672_), .A2(new_n677_), .ZN(G1329gat));
  INV_X1    g477(.A(KEYINPUT47), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n666_), .A2(new_n667_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(new_n302_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(G43gat), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n635_), .A2(G43gat), .A3(new_n303_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n679_), .B1(new_n682_), .B2(new_n684_), .ZN(new_n685_));
  AOI211_X1 g484(.A(KEYINPUT47), .B(new_n683_), .C1(new_n681_), .C2(G43gat), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1330gat));
  AOI21_X1  g486(.A(G50gat), .B1(new_n636_), .B2(new_n617_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n617_), .A2(G50gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n680_), .B2(new_n689_), .ZN(G1331gat));
  INV_X1    g489(.A(G57gat), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n535_), .A2(new_n239_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n438_), .B2(new_n456_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n587_), .B1(new_n559_), .B2(new_n565_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n691_), .B1(new_n695_), .B2(new_n455_), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT107), .Z(new_n697_));
  NOR2_X1   g496(.A1(new_n692_), .A2(new_n587_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(new_n594_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n699_), .A2(new_n691_), .A3(new_n455_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n697_), .A2(new_n700_), .ZN(G1332gat));
  OAI21_X1  g500(.A(G64gat), .B1(new_n699_), .B2(new_n449_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT48), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n449_), .A2(G64gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(new_n695_), .B2(new_n704_), .ZN(G1333gat));
  OR3_X1    g504(.A1(new_n695_), .A2(G71gat), .A3(new_n303_), .ZN(new_n706_));
  OAI21_X1  g505(.A(G71gat), .B1(new_n699_), .B2(new_n303_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n707_), .A2(KEYINPUT49), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(KEYINPUT49), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n706_), .B1(new_n708_), .B2(new_n709_), .ZN(G1334gat));
  NAND3_X1  g509(.A1(new_n698_), .A2(new_n617_), .A3(new_n594_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT50), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n711_), .A2(new_n712_), .A3(G78gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n711_), .B2(G78gat), .ZN(new_n714_));
  OR2_X1    g513(.A1(new_n348_), .A2(G78gat), .ZN(new_n715_));
  OAI22_X1  g514(.A1(new_n713_), .A2(new_n714_), .B1(new_n695_), .B2(new_n715_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT108), .Z(G1335gat));
  NOR2_X1   g516(.A1(new_n692_), .A2(new_n629_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n646_), .A2(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n719_), .A2(KEYINPUT109), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT110), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT109), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n722_), .B1(new_n646_), .B2(new_n718_), .ZN(new_n723_));
  OR3_X1    g522(.A1(new_n720_), .A2(new_n721_), .A3(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n721_), .B1(new_n720_), .B2(new_n723_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n724_), .A2(new_n383_), .A3(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(G85gat), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n693_), .A2(new_n630_), .ZN(new_n728_));
  OR3_X1    g527(.A1(new_n728_), .A2(G85gat), .A3(new_n455_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1336gat));
  INV_X1    g529(.A(new_n728_), .ZN(new_n731_));
  AOI21_X1  g530(.A(G92gat), .B1(new_n731_), .B2(new_n602_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n724_), .A2(new_n725_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n602_), .A2(G92gat), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT111), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n732_), .B1(new_n733_), .B2(new_n735_), .ZN(G1337gat));
  NOR3_X1   g535(.A1(new_n303_), .A2(new_n474_), .A3(new_n473_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(KEYINPUT112), .B1(new_n728_), .B2(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n302_), .B1(new_n720_), .B2(new_n723_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n740_), .B2(G99gat), .ZN(new_n741_));
  XNOR2_X1  g540(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n741_), .B(new_n743_), .ZN(G1338gat));
  NAND3_X1  g543(.A1(new_n731_), .A2(new_n485_), .A3(new_n617_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT114), .ZN(new_n746_));
  OAI21_X1  g545(.A(G106gat), .B1(new_n719_), .B2(new_n348_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n748_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n746_), .A2(new_n749_), .A3(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT53), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT53), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n746_), .A2(new_n749_), .A3(new_n753_), .A4(new_n750_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(G1339gat));
  INV_X1    g554(.A(KEYINPUT120), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n694_), .B(new_n239_), .C1(new_n533_), .C2(new_n534_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT54), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n757_), .B(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n227_), .A2(new_n233_), .A3(new_n236_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n202_), .B1(new_n223_), .B2(new_n226_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n228_), .A2(new_n232_), .A3(new_n203_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n236_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n761_), .A2(new_n762_), .A3(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n760_), .A2(new_n764_), .A3(new_n524_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n518_), .A2(KEYINPUT115), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT55), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n518_), .A2(KEYINPUT115), .A3(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n459_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n513_), .A2(new_n515_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n507_), .A2(new_n517_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n771_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT116), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n776_), .B(new_n771_), .C1(new_n772_), .C2(new_n773_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n768_), .A2(new_n770_), .A3(new_n775_), .A4(new_n777_), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n778_), .A2(KEYINPUT56), .A3(new_n522_), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT56), .B1(new_n778_), .B2(new_n522_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n766_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT118), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n566_), .B1(new_n782_), .B2(KEYINPUT58), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT58), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n781_), .A2(KEYINPUT118), .A3(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n524_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n778_), .A2(new_n522_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT56), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n778_), .A2(KEYINPUT56), .A3(new_n522_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n786_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n760_), .A2(new_n764_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n792_), .A2(new_n527_), .A3(new_n530_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  OAI211_X1 g593(.A(KEYINPUT57), .B(new_n628_), .C1(new_n791_), .C2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT119), .ZN(new_n796_));
  AOI22_X1  g595(.A1(new_n783_), .A2(new_n785_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n628_), .B1(new_n791_), .B2(new_n794_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT117), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT117), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n801_), .B(new_n628_), .C1(new_n791_), .C2(new_n794_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n799_), .A2(new_n800_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n238_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n525_), .B1(new_n804_), .B2(new_n760_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n805_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n593_), .B1(new_n806_), .B2(new_n793_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n807_), .A2(KEYINPUT119), .A3(KEYINPUT57), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n797_), .A2(new_n803_), .A3(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n759_), .B1(new_n809_), .B2(new_n587_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n602_), .A2(new_n455_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n452_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n756_), .B1(new_n810_), .B2(new_n813_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n799_), .A2(new_n800_), .A3(new_n802_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n765_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT118), .ZN(new_n817_));
  OAI21_X1  g616(.A(KEYINPUT58), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n818_), .A2(new_n567_), .A3(new_n785_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n795_), .A2(new_n796_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n820_), .A3(new_n808_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n587_), .B1(new_n815_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n759_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n813_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n824_), .A2(KEYINPUT120), .A3(new_n825_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n814_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(G113gat), .B1(new_n827_), .B2(new_n627_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT59), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n810_), .B2(new_n813_), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n819_), .A2(new_n820_), .A3(new_n808_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n629_), .B1(new_n831_), .B2(new_n803_), .ZN(new_n832_));
  OAI211_X1 g631(.A(KEYINPUT59), .B(new_n825_), .C1(new_n832_), .C2(new_n759_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n830_), .A2(new_n833_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n239_), .A2(KEYINPUT121), .ZN(new_n835_));
  MUX2_X1   g634(.A(KEYINPUT121), .B(new_n835_), .S(G113gat), .Z(new_n836_));
  AOI21_X1  g635(.A(new_n828_), .B1(new_n834_), .B2(new_n836_), .ZN(G1340gat));
  NAND2_X1  g636(.A1(new_n834_), .A2(new_n535_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(G120gat), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n626_), .A2(KEYINPUT60), .ZN(new_n840_));
  MUX2_X1   g639(.A(new_n840_), .B(KEYINPUT60), .S(G120gat), .Z(new_n841_));
  NAND2_X1  g640(.A1(new_n827_), .A2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n839_), .A2(new_n842_), .ZN(G1341gat));
  INV_X1    g642(.A(G127gat), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n814_), .A2(new_n826_), .A3(new_n844_), .A4(new_n629_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n587_), .B1(new_n830_), .B2(new_n833_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(new_n844_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT122), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT122), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n845_), .B(new_n849_), .C1(new_n846_), .C2(new_n844_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n850_), .ZN(G1342gat));
  INV_X1    g650(.A(G134gat), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n827_), .A2(new_n852_), .A3(new_n593_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n566_), .B1(new_n830_), .B2(new_n833_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n852_), .B2(new_n854_), .ZN(G1343gat));
  INV_X1    g654(.A(new_n453_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n811_), .A2(new_n856_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(KEYINPUT123), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n824_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n627_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n535_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G148gat), .ZN(G1345gat));
  OR3_X1    g663(.A1(new_n859_), .A2(KEYINPUT124), .A3(new_n587_), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT124), .B1(new_n859_), .B2(new_n587_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(KEYINPUT61), .B(G155gat), .ZN(new_n867_));
  AND3_X1   g666(.A1(new_n865_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n868_), .A2(new_n869_), .ZN(G1346gat));
  OR3_X1    g669(.A1(new_n859_), .A2(G162gat), .A3(new_n628_), .ZN(new_n871_));
  OAI21_X1  g670(.A(G162gat), .B1(new_n859_), .B2(new_n566_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(G1347gat));
  NOR3_X1   g672(.A1(new_n449_), .A2(new_n383_), .A3(new_n452_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n824_), .A2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n627_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(G169gat), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT62), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n876_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n880_));
  INV_X1    g679(.A(new_n258_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n879_), .B(new_n880_), .C1(new_n881_), .C2(new_n876_), .ZN(G1348gat));
  NAND3_X1  g681(.A1(new_n824_), .A2(new_n535_), .A3(new_n874_), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n883_), .A2(G176gat), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT125), .ZN(new_n885_));
  INV_X1    g684(.A(new_n257_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n883_), .A2(new_n886_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n884_), .A2(new_n885_), .A3(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n885_), .B1(new_n884_), .B2(new_n887_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1349gat));
  NAND2_X1  g690(.A1(new_n875_), .A2(new_n629_), .ZN(new_n892_));
  MUX2_X1   g691(.A(new_n247_), .B(G183gat), .S(new_n892_), .Z(G1350gat));
  NAND3_X1  g692(.A1(new_n875_), .A2(new_n248_), .A3(new_n593_), .ZN(new_n894_));
  AND2_X1   g693(.A1(new_n875_), .A2(new_n567_), .ZN(new_n895_));
  INV_X1    g694(.A(G190gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n894_), .B1(new_n895_), .B2(new_n896_), .ZN(G1351gat));
  NOR2_X1   g696(.A1(new_n449_), .A2(new_n383_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n856_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(KEYINPUT126), .B1(new_n824_), .B2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT126), .ZN(new_n902_));
  AOI211_X1 g701(.A(new_n902_), .B(new_n899_), .C1(new_n822_), .C2(new_n823_), .ZN(new_n903_));
  OAI211_X1 g702(.A(G197gat), .B(new_n627_), .C1(new_n901_), .C2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(KEYINPUT127), .ZN(new_n905_));
  INV_X1    g704(.A(G197gat), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n901_), .A2(new_n903_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n907_), .B2(new_n239_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n902_), .B1(new_n810_), .B2(new_n899_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n824_), .A2(KEYINPUT126), .A3(new_n900_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT127), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n911_), .A2(new_n912_), .A3(G197gat), .A4(new_n627_), .ZN(new_n913_));
  AND3_X1   g712(.A1(new_n905_), .A2(new_n908_), .A3(new_n913_), .ZN(G1352gat));
  NAND2_X1  g713(.A1(new_n911_), .A2(new_n535_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(G204gat), .ZN(G1353gat));
  OR2_X1    g715(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n917_));
  NAND2_X1  g716(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n918_));
  AND4_X1   g717(.A1(new_n629_), .A2(new_n911_), .A3(new_n917_), .A4(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n917_), .B1(new_n911_), .B2(new_n629_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n919_), .A2(new_n920_), .ZN(G1354gat));
  OR3_X1    g720(.A1(new_n907_), .A2(G218gat), .A3(new_n628_), .ZN(new_n922_));
  OAI21_X1  g721(.A(G218gat), .B1(new_n907_), .B2(new_n566_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(G1355gat));
endmodule


