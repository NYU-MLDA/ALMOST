//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 1 0 0 1 1 1 1 1 0 0 0 0 1 0 1 1 0 0 0 1 1 0 0 1 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n921_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n955_, new_n956_, new_n957_, new_n959_,
    new_n960_, new_n961_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n968_, new_n969_, new_n970_, new_n971_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n978_, new_n980_,
    new_n981_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n990_, new_n991_, new_n992_;
  INV_X1    g000(.A(KEYINPUT38), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT7), .ZN(new_n203_));
  INV_X1    g002(.A(G99gat), .ZN(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT6), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n206_), .A2(new_n209_), .A3(new_n210_), .A4(new_n211_), .ZN(new_n212_));
  OR2_X1    g011(.A1(G85gat), .A2(G92gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G85gat), .A2(G92gat), .ZN(new_n214_));
  AND2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT8), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n204_), .A2(KEYINPUT10), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n204_), .A2(KEYINPUT10), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n205_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n209_), .A2(new_n210_), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n214_), .A2(KEYINPUT9), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n213_), .A2(KEYINPUT9), .A3(new_n214_), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .A4(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n212_), .A2(KEYINPUT8), .A3(new_n215_), .ZN(new_n226_));
  AND3_X1   g025(.A1(new_n218_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n228_));
  INV_X1    g027(.A(G57gat), .ZN(new_n229_));
  INV_X1    g028(.A(G64gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G57gat), .A2(G64gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT11), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G71gat), .B(G78gat), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT11), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n231_), .A2(new_n237_), .A3(new_n232_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n234_), .A2(new_n236_), .A3(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n233_), .A2(new_n235_), .A3(KEYINPUT11), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n227_), .A2(new_n228_), .A3(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n218_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n241_), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT64), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n242_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n243_), .A2(new_n244_), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n247_), .A2(KEYINPUT65), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(KEYINPUT65), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n246_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G230gat), .A2(G233gat), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n247_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT12), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT12), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n247_), .A2(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n252_), .B1(new_n227_), .B2(new_n241_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n255_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(G120gat), .B(G148gat), .Z(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT66), .B(KEYINPUT5), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G176gat), .B(G204gat), .ZN(new_n263_));
  XOR2_X1   g062(.A(new_n262_), .B(new_n263_), .Z(new_n264_));
  NAND3_X1  g063(.A1(new_n253_), .A2(new_n259_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n264_), .B1(new_n253_), .B2(new_n259_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT67), .ZN(new_n268_));
  OAI22_X1  g067(.A1(new_n266_), .A2(new_n267_), .B1(new_n268_), .B2(KEYINPUT13), .ZN(new_n269_));
  INV_X1    g068(.A(new_n267_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT67), .B(KEYINPUT13), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n270_), .A2(new_n265_), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n269_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT37), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G190gat), .B(G218gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(G134gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(G162gat), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n279_), .A2(KEYINPUT36), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G232gat), .A2(G233gat), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT68), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT34), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT35), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(G50gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G29gat), .A2(G36gat), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(G29gat), .A2(G36gat), .ZN(new_n291_));
  NOR3_X1   g090(.A1(new_n290_), .A2(new_n291_), .A3(G43gat), .ZN(new_n292_));
  INV_X1    g091(.A(G43gat), .ZN(new_n293_));
  INV_X1    g092(.A(G29gat), .ZN(new_n294_));
  INV_X1    g093(.A(G36gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n293_), .B1(new_n296_), .B2(new_n289_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n288_), .B1(new_n292_), .B2(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(G43gat), .B1(new_n290_), .B2(new_n291_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n296_), .A2(new_n293_), .A3(new_n289_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n299_), .A2(new_n300_), .A3(G50gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n287_), .B1(new_n243_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT69), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n285_), .A2(new_n286_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n298_), .A2(KEYINPUT15), .A3(new_n301_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(KEYINPUT15), .B1(new_n298_), .B2(new_n301_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n243_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n304_), .A2(new_n305_), .A3(new_n306_), .A4(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n306_), .A2(new_n305_), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT69), .B1(new_n285_), .B2(new_n286_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n226_), .ZN(new_n314_));
  AOI21_X1  g113(.A(KEYINPUT8), .B1(new_n212_), .B2(new_n215_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT15), .ZN(new_n317_));
  AND3_X1   g116(.A1(new_n299_), .A2(new_n300_), .A3(G50gat), .ZN(new_n318_));
  AOI21_X1  g117(.A(G50gat), .B1(new_n299_), .B2(new_n300_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n317_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  AOI22_X1  g119(.A1(new_n316_), .A2(new_n225_), .B1(new_n320_), .B2(new_n307_), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n312_), .B(new_n313_), .C1(new_n321_), .C2(new_n303_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n311_), .A2(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n281_), .B1(new_n323_), .B2(KEYINPUT70), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT70), .ZN(new_n325_));
  AOI211_X1 g124(.A(new_n325_), .B(new_n280_), .C1(new_n311_), .C2(new_n322_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n279_), .A2(KEYINPUT36), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n311_), .A2(new_n322_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n276_), .B1(new_n327_), .B2(new_n330_), .ZN(new_n331_));
  NOR4_X1   g130(.A1(new_n324_), .A2(new_n326_), .A3(KEYINPUT71), .A4(new_n329_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n275_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n323_), .A2(KEYINPUT70), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n280_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n323_), .A2(KEYINPUT70), .A3(new_n281_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(new_n336_), .A3(new_n330_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT71), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n327_), .A2(new_n276_), .A3(new_n330_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n338_), .A2(new_n339_), .A3(KEYINPUT37), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n333_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT16), .B(G183gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(G211gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G127gat), .B(G155gat), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n344_), .B(new_n345_), .Z(new_n346_));
  INV_X1    g145(.A(KEYINPUT17), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT72), .B(G22gat), .ZN(new_n349_));
  INV_X1    g148(.A(G15gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(G1gat), .ZN(new_n352_));
  INV_X1    g151(.A(G8gat), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT14), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n351_), .A2(new_n354_), .ZN(new_n355_));
  XOR2_X1   g154(.A(G1gat), .B(G8gat), .Z(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n351_), .A2(new_n356_), .A3(new_n354_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(new_n244_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G231gat), .A2(G233gat), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n358_), .A2(new_n359_), .A3(new_n241_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n361_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n362_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n348_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n366_), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n346_), .A2(new_n347_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(new_n364_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT73), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n367_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n371_), .B1(new_n367_), .B2(new_n370_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n342_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT27), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G226gat), .A2(G233gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT19), .ZN(new_n379_));
  XOR2_X1   g178(.A(G211gat), .B(G218gat), .Z(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(G204gat), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n382_), .A2(G197gat), .ZN(new_n383_));
  INV_X1    g182(.A(G197gat), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT85), .B1(new_n384_), .B2(G204gat), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT85), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(new_n382_), .A3(G197gat), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n383_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT21), .ZN(new_n389_));
  NOR3_X1   g188(.A1(new_n381_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n382_), .A2(G197gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n384_), .A2(G204gat), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(new_n392_), .A3(KEYINPUT84), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n393_), .B(KEYINPUT21), .C1(KEYINPUT84), .C2(new_n391_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT86), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n385_), .A2(new_n387_), .ZN(new_n396_));
  AND4_X1   g195(.A1(new_n395_), .A2(new_n396_), .A3(new_n389_), .A4(new_n392_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n395_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n394_), .B(new_n381_), .C1(new_n397_), .C2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT87), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n386_), .B1(G197gat), .B2(new_n382_), .ZN(new_n401_));
  NOR3_X1   g200(.A1(new_n384_), .A2(KEYINPUT85), .A3(G204gat), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n389_), .B(new_n392_), .C1(new_n401_), .C2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT86), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n388_), .A2(new_n395_), .A3(new_n389_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT87), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n406_), .A2(new_n407_), .A3(new_n394_), .A4(new_n381_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n390_), .B1(new_n400_), .B2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT25), .B(G183gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT26), .B(G190gat), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT92), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n413_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n411_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G169gat), .A2(G176gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NOR3_X1   g219(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G183gat), .A2(G190gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT75), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT75), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n426_), .A2(G183gat), .A3(G190gat), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n425_), .A2(new_n427_), .A3(KEYINPUT23), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT23), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n424_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(new_n430_), .ZN(new_n431_));
  NOR3_X1   g230(.A1(new_n416_), .A2(new_n423_), .A3(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n425_), .A2(new_n427_), .A3(new_n429_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n424_), .A2(KEYINPUT23), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(G183gat), .ZN(new_n436_));
  INV_X1    g235(.A(G190gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT76), .B(G176gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT22), .B(G169gat), .ZN(new_n440_));
  AOI22_X1  g239(.A1(new_n435_), .A2(new_n438_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(new_n417_), .B(KEYINPUT93), .Z(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT94), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n441_), .A2(KEYINPUT94), .A3(new_n442_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n432_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT20), .B1(new_n409_), .B2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n428_), .A2(new_n438_), .A3(new_n430_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n439_), .A2(new_n440_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(new_n417_), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n410_), .A2(new_n412_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n435_), .A2(new_n422_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  AOI211_X1 g253(.A(new_n454_), .B(new_n390_), .C1(new_n400_), .C2(new_n408_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n379_), .B1(new_n448_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n457_));
  INV_X1    g256(.A(new_n390_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n408_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n380_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n407_), .B1(new_n460_), .B2(new_n394_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n458_), .B1(new_n459_), .B2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n457_), .B1(new_n462_), .B2(new_n454_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n379_), .B1(new_n409_), .B2(new_n447_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(G8gat), .B(G36gat), .Z(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G64gat), .B(G92gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  AND3_X1   g269(.A1(new_n456_), .A2(new_n465_), .A3(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n470_), .B1(new_n456_), .B2(new_n465_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n377_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n470_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n379_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n432_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n409_), .A2(new_n476_), .A3(new_n443_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n475_), .B1(new_n463_), .B2(new_n477_), .ZN(new_n478_));
  NOR3_X1   g277(.A1(new_n448_), .A2(new_n379_), .A3(new_n455_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n474_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n456_), .A2(new_n465_), .A3(new_n470_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n480_), .A2(KEYINPUT27), .A3(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT0), .B(G57gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(G85gat), .ZN(new_n484_));
  XOR2_X1   g283(.A(G1gat), .B(G29gat), .Z(new_n485_));
  XOR2_X1   g284(.A(new_n484_), .B(new_n485_), .Z(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT4), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT78), .ZN(new_n489_));
  OR2_X1    g288(.A1(G127gat), .A2(G134gat), .ZN(new_n490_));
  INV_X1    g289(.A(G113gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G127gat), .A2(G134gat), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  AND2_X1   g292(.A1(G127gat), .A2(G134gat), .ZN(new_n494_));
  NOR2_X1   g293(.A1(G127gat), .A2(G134gat), .ZN(new_n495_));
  OAI21_X1  g294(.A(G113gat), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n493_), .A2(new_n496_), .A3(G120gat), .ZN(new_n497_));
  AOI21_X1  g296(.A(G120gat), .B1(new_n493_), .B2(new_n496_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n489_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n493_), .A2(new_n496_), .ZN(new_n500_));
  INV_X1    g299(.A(G120gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n493_), .A2(new_n496_), .A3(G120gat), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(KEYINPUT78), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n499_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G155gat), .A2(G162gat), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT81), .B1(new_n506_), .B2(KEYINPUT1), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT81), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT1), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n508_), .A2(new_n509_), .A3(G155gat), .A4(G162gat), .ZN(new_n510_));
  OR2_X1    g309(.A1(G155gat), .A2(G162gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n506_), .A2(KEYINPUT1), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n507_), .A2(new_n510_), .A3(new_n511_), .A4(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(G141gat), .ZN(new_n514_));
  INV_X1    g313(.A(G148gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G141gat), .A2(G148gat), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n513_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT3), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n519_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT2), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n517_), .A2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n523_));
  NAND3_X1  g322(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n520_), .A2(new_n522_), .A3(new_n523_), .A4(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT82), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n511_), .B(new_n506_), .C1(new_n525_), .C2(new_n526_), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n525_), .A2(new_n526_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n518_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n505_), .A2(new_n529_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n525_), .A2(new_n526_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n525_), .A2(new_n526_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n531_), .A2(new_n532_), .A3(new_n511_), .A4(new_n506_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT96), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n534_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n502_), .A2(KEYINPUT96), .A3(new_n503_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n533_), .A2(new_n535_), .A3(new_n536_), .A4(new_n518_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n488_), .B1(new_n530_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G225gat), .A2(G233gat), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT4), .B1(new_n505_), .B2(new_n529_), .ZN(new_n540_));
  NOR3_X1   g339(.A1(new_n538_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n530_), .A2(new_n537_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(new_n539_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n487_), .B1(new_n541_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(KEYINPUT4), .ZN(new_n546_));
  INV_X1    g345(.A(new_n539_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n540_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n546_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n549_), .A2(new_n543_), .A3(new_n486_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n545_), .A2(new_n550_), .A3(KEYINPUT98), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT98), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n552_), .B(new_n487_), .C1(new_n541_), .C2(new_n544_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n473_), .A2(new_n482_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT80), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G15gat), .B(G43gat), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G227gat), .A2(G233gat), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n557_), .B(new_n558_), .Z(new_n559_));
  INV_X1    g358(.A(KEYINPUT30), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n451_), .A2(new_n453_), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n560_), .B1(new_n451_), .B2(new_n453_), .ZN(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT79), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n454_), .A2(KEYINPUT30), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT79), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n565_), .A2(new_n566_), .A3(new_n561_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n505_), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n564_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n568_), .B1(new_n564_), .B2(new_n567_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n559_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G71gat), .B(G99gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT77), .B(KEYINPUT31), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n562_), .A2(new_n563_), .A3(KEYINPUT79), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n566_), .B1(new_n565_), .B2(new_n561_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n505_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n564_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n559_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n577_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n571_), .A2(new_n574_), .A3(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n574_), .B1(new_n571_), .B2(new_n580_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n556_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n574_), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n569_), .A2(new_n570_), .A3(new_n559_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n579_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n584_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n571_), .A2(new_n580_), .A3(new_n574_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(KEYINPUT80), .A3(new_n588_), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n529_), .A2(KEYINPUT29), .ZN(new_n590_));
  XOR2_X1   g389(.A(KEYINPUT83), .B(KEYINPUT28), .Z(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G22gat), .B(G50gat), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n592_), .B(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(G228gat), .ZN(new_n596_));
  INV_X1    g395(.A(G233gat), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT88), .B(KEYINPUT29), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n529_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT89), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n529_), .A2(KEYINPUT89), .A3(new_n599_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n598_), .B1(new_n604_), .B2(new_n409_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n598_), .B1(new_n529_), .B2(KEYINPUT29), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n462_), .A2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G78gat), .B(G106gat), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT90), .Z(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n605_), .A2(new_n607_), .A3(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n605_), .A2(new_n607_), .A3(KEYINPUT91), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(new_n608_), .ZN(new_n613_));
  AOI21_X1  g412(.A(KEYINPUT91), .B1(new_n605_), .B2(new_n607_), .ZN(new_n614_));
  OAI211_X1 g413(.A(new_n595_), .B(new_n611_), .C1(new_n613_), .C2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n592_), .B(new_n593_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n611_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n610_), .B1(new_n605_), .B2(new_n607_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n616_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  AOI22_X1  g418(.A1(new_n583_), .A2(new_n589_), .B1(new_n615_), .B2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n587_), .A2(new_n588_), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n615_), .A2(new_n621_), .A3(new_n619_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n555_), .B1(new_n620_), .B2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n456_), .A2(new_n465_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(new_n474_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT97), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n542_), .A2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n530_), .A2(new_n537_), .A3(KEYINPUT97), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(new_n547_), .A3(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n539_), .B1(new_n538_), .B2(new_n540_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(new_n486_), .A3(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n625_), .A2(new_n481_), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT33), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n545_), .B(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n470_), .A2(KEYINPUT32), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n456_), .A2(new_n465_), .A3(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n551_), .A2(new_n553_), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n478_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n479_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n635_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  OAI22_X1  g439(.A1(new_n632_), .A2(new_n634_), .B1(new_n637_), .B2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n583_), .A2(new_n589_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n615_), .A2(new_n619_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n641_), .A2(new_n642_), .A3(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n623_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n302_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n358_), .A2(new_n359_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n647_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n650_));
  OAI211_X1 g449(.A(G229gat), .B(G233gat), .C1(new_n649_), .C2(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n360_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(G229gat), .A2(G233gat), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(new_n653_), .A3(new_n648_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n651_), .A2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(G169gat), .B(G197gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(G141gat), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT74), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(new_n491_), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n655_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n655_), .A2(new_n659_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT99), .B1(new_n646_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT99), .ZN(new_n664_));
  INV_X1    g463(.A(new_n662_), .ZN(new_n665_));
  AOI211_X1 g464(.A(new_n664_), .B(new_n665_), .C1(new_n623_), .C2(new_n645_), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n274_), .B(new_n376_), .C1(new_n663_), .C2(new_n666_), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n667_), .A2(KEYINPUT100), .ZN(new_n668_));
  INV_X1    g467(.A(new_n554_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(KEYINPUT100), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n668_), .A2(new_n352_), .A3(new_n669_), .A4(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT101), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n671_), .A2(KEYINPUT101), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n202_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n671_), .A2(KEYINPUT101), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n676_), .A2(KEYINPUT38), .A3(new_n672_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n646_), .A2(new_n662_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n274_), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n680_), .A2(new_n375_), .A3(new_n337_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(G1gat), .B1(new_n682_), .B2(new_n554_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n675_), .A2(new_n677_), .A3(new_n683_), .ZN(G1324gat));
  NAND2_X1  g483(.A1(new_n473_), .A2(new_n482_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n679_), .A2(new_n685_), .A3(new_n681_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n686_), .A2(new_n687_), .A3(G8gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n686_), .B2(G8gat), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT39), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n688_), .A2(new_n689_), .A3(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n686_), .A2(G8gat), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT102), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n686_), .A2(new_n687_), .A3(G8gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(KEYINPUT39), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n691_), .A2(new_n695_), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n668_), .A2(new_n353_), .A3(new_n685_), .A4(new_n670_), .ZN(new_n697_));
  XOR2_X1   g496(.A(KEYINPUT103), .B(KEYINPUT104), .Z(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT40), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n696_), .A2(new_n697_), .A3(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1325gat));
  OAI21_X1  g501(.A(G15gat), .B1(new_n682_), .B2(new_n642_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT41), .Z(new_n704_));
  NAND2_X1  g503(.A1(new_n668_), .A2(new_n670_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n642_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(new_n350_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n704_), .B1(new_n705_), .B2(new_n707_), .ZN(G1326gat));
  OAI21_X1  g507(.A(G22gat), .B1(new_n682_), .B2(new_n644_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT105), .Z(new_n710_));
  AND2_X1   g509(.A1(new_n710_), .A2(KEYINPUT42), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(KEYINPUT42), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n644_), .A2(G22gat), .ZN(new_n713_));
  OAI22_X1  g512(.A1(new_n711_), .A2(new_n712_), .B1(new_n705_), .B2(new_n713_), .ZN(G1327gat));
  NOR3_X1   g513(.A1(new_n680_), .A2(new_n665_), .A3(new_n374_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n646_), .B2(new_n342_), .ZN(new_n717_));
  AOI211_X1 g516(.A(KEYINPUT43), .B(new_n341_), .C1(new_n623_), .C2(new_n645_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n715_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  OAI211_X1 g520(.A(KEYINPUT44), .B(new_n715_), .C1(new_n717_), .C2(new_n718_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n723_), .A2(G29gat), .A3(new_n669_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n337_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n374_), .A2(new_n725_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n274_), .B(new_n726_), .C1(new_n663_), .C2(new_n666_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n294_), .B1(new_n727_), .B2(new_n554_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n724_), .A2(new_n728_), .ZN(G1328gat));
  NOR2_X1   g528(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT45), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT107), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n727_), .A2(G36gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(new_n685_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n685_), .ZN(new_n735_));
  NOR4_X1   g534(.A1(new_n727_), .A2(KEYINPUT107), .A3(G36gat), .A4(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n731_), .B1(new_n734_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n663_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n646_), .A2(KEYINPUT99), .A3(new_n662_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n680_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n740_), .A2(new_n295_), .A3(new_n685_), .A4(new_n726_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT107), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n733_), .A2(new_n732_), .A3(new_n685_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n742_), .A2(new_n743_), .A3(KEYINPUT45), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n737_), .A2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n721_), .A2(new_n685_), .A3(new_n722_), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n746_), .A2(KEYINPUT106), .A3(G36gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(KEYINPUT106), .B1(new_n746_), .B2(G36gat), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n730_), .B1(new_n745_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n746_), .A2(G36gat), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT106), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n746_), .A2(KEYINPUT106), .A3(G36gat), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n730_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n755_), .A2(new_n756_), .A3(new_n744_), .A4(new_n737_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n750_), .A2(new_n757_), .ZN(G1329gat));
  INV_X1    g557(.A(KEYINPUT47), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n721_), .A2(new_n621_), .A3(new_n722_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(G43gat), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n762_));
  INV_X1    g561(.A(new_n727_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n763_), .A2(new_n293_), .A3(new_n706_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n761_), .A2(new_n762_), .A3(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n762_), .B1(new_n761_), .B2(new_n764_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n759_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n767_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n769_), .A2(KEYINPUT47), .A3(new_n765_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(G1330gat));
  AOI21_X1  g570(.A(G50gat), .B1(new_n763_), .B2(new_n643_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n644_), .A2(new_n288_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n723_), .B2(new_n773_), .ZN(G1331gat));
  AND2_X1   g573(.A1(new_n623_), .A2(new_n645_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n274_), .A2(new_n662_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n775_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n376_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(G57gat), .B1(new_n780_), .B2(new_n669_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n375_), .A2(new_n337_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n778_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n229_), .B1(new_n669_), .B2(KEYINPUT110), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n229_), .A2(KEYINPUT110), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n781_), .B1(new_n786_), .B2(new_n787_), .ZN(G1332gat));
  AOI21_X1  g587(.A(new_n230_), .B1(new_n783_), .B2(new_n685_), .ZN(new_n789_));
  XOR2_X1   g588(.A(new_n789_), .B(KEYINPUT48), .Z(new_n790_));
  NAND3_X1  g589(.A1(new_n780_), .A2(new_n230_), .A3(new_n685_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(G1333gat));
  INV_X1    g591(.A(G71gat), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n793_), .B1(new_n783_), .B2(new_n706_), .ZN(new_n794_));
  XOR2_X1   g593(.A(new_n794_), .B(KEYINPUT49), .Z(new_n795_));
  NAND3_X1  g594(.A1(new_n780_), .A2(new_n793_), .A3(new_n706_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(G1334gat));
  INV_X1    g596(.A(G78gat), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n798_), .B1(new_n783_), .B2(new_n643_), .ZN(new_n799_));
  XOR2_X1   g598(.A(new_n799_), .B(KEYINPUT50), .Z(new_n800_));
  NAND3_X1  g599(.A1(new_n780_), .A2(new_n798_), .A3(new_n643_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(G1335gat));
  OAI211_X1 g601(.A(new_n375_), .B(new_n776_), .C1(new_n717_), .C2(new_n718_), .ZN(new_n803_));
  INV_X1    g602(.A(G85gat), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n803_), .A2(new_n804_), .A3(new_n554_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n778_), .A2(new_n726_), .ZN(new_n806_));
  AOI21_X1  g605(.A(G85gat), .B1(new_n806_), .B2(new_n669_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n805_), .A2(new_n807_), .ZN(G1336gat));
  AOI21_X1  g607(.A(G92gat), .B1(new_n806_), .B2(new_n685_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n803_), .A2(new_n735_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(G92gat), .ZN(G1337gat));
  OAI211_X1 g610(.A(new_n806_), .B(new_n621_), .C1(new_n219_), .C2(new_n220_), .ZN(new_n812_));
  OAI21_X1  g611(.A(G99gat), .B1(new_n803_), .B2(new_n642_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n815_), .A2(KEYINPUT111), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n814_), .B(new_n816_), .ZN(G1338gat));
  NOR2_X1   g616(.A1(new_n644_), .A2(G106gat), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n806_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n820_));
  INV_X1    g619(.A(new_n717_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n718_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n823_), .A2(new_n643_), .A3(new_n375_), .A4(new_n776_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n820_), .B1(new_n824_), .B2(G106gat), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n820_), .B(G106gat), .C1(new_n803_), .C2(new_n644_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n819_), .B1(new_n825_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT112), .ZN(new_n829_));
  OAI21_X1  g628(.A(G106gat), .B1(new_n803_), .B2(new_n644_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT52), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n826_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT112), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(new_n833_), .A3(new_n819_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n829_), .A2(KEYINPUT53), .A3(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT53), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n833_), .B1(new_n832_), .B2(new_n819_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n819_), .ZN(new_n838_));
  AOI211_X1 g637(.A(KEYINPUT112), .B(new_n838_), .C1(new_n831_), .C2(new_n826_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n836_), .B1(new_n837_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n835_), .A2(new_n840_), .ZN(G1339gat));
  NOR2_X1   g640(.A1(new_n685_), .A2(new_n554_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n653_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n652_), .A2(new_n648_), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n843_), .B(new_n659_), .C1(new_n844_), .C2(new_n653_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n660_), .A2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n846_), .B1(new_n267_), .B2(new_n266_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT55), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n259_), .A2(new_n848_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n247_), .B(KEYINPUT12), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n850_), .A2(KEYINPUT55), .A3(new_n258_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n850_), .A2(new_n246_), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n849_), .B(new_n851_), .C1(new_n852_), .C2(new_n251_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT56), .ZN(new_n854_));
  INV_X1    g653(.A(new_n264_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n853_), .A2(KEYINPUT115), .A3(new_n854_), .A4(new_n855_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n853_), .A2(new_n855_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n265_), .B(new_n856_), .C1(new_n857_), .C2(new_n854_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n662_), .B1(new_n857_), .B2(KEYINPUT115), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n847_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n860_), .A2(KEYINPUT57), .A3(new_n725_), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT57), .B1(new_n860_), .B2(new_n725_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n857_), .A2(new_n854_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n853_), .A2(new_n855_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n266_), .B1(new_n865_), .B2(KEYINPUT56), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n864_), .A2(new_n866_), .A3(new_n846_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT58), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n864_), .A2(new_n866_), .A3(KEYINPUT58), .A4(new_n846_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n342_), .A2(new_n869_), .A3(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n374_), .B1(new_n863_), .B2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n662_), .B1(new_n269_), .B2(new_n273_), .ZN(new_n873_));
  AND3_X1   g672(.A1(new_n873_), .A2(KEYINPUT113), .A3(new_n374_), .ZN(new_n874_));
  AOI21_X1  g673(.A(KEYINPUT113), .B1(new_n873_), .B2(new_n374_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT114), .ZN(new_n878_));
  OR2_X1    g677(.A1(new_n877_), .A2(KEYINPUT114), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n876_), .A2(new_n341_), .A3(new_n878_), .A4(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n274_), .A2(new_n665_), .A3(new_n374_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT113), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n873_), .A2(KEYINPUT113), .A3(new_n374_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n883_), .A2(new_n341_), .A3(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n885_), .A2(KEYINPUT114), .A3(new_n877_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n880_), .A2(new_n886_), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n622_), .B(new_n842_), .C1(new_n872_), .C2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(G113gat), .B1(new_n889_), .B2(new_n662_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT116), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n888_), .A2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n888_), .A2(new_n892_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n891_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n889_), .A2(KEYINPUT59), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n897_), .A2(KEYINPUT116), .A3(new_n893_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n665_), .B1(new_n896_), .B2(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n890_), .B1(new_n899_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g699(.A(new_n501_), .B1(new_n274_), .B2(KEYINPUT60), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n889_), .B(new_n901_), .C1(KEYINPUT60), .C2(new_n501_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n274_), .B1(new_n897_), .B2(new_n893_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n903_), .B2(new_n501_), .ZN(G1341gat));
  AOI21_X1  g703(.A(G127gat), .B1(new_n889_), .B2(new_n374_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n375_), .B1(new_n896_), .B2(new_n898_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n905_), .B1(new_n906_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g706(.A(G134gat), .B1(new_n889_), .B2(new_n337_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n341_), .B1(new_n896_), .B2(new_n898_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n908_), .B1(new_n909_), .B2(G134gat), .ZN(G1343gat));
  AND2_X1   g709(.A1(new_n880_), .A2(new_n886_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n862_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n860_), .A2(KEYINPUT57), .A3(new_n725_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n912_), .A2(new_n913_), .A3(new_n871_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(new_n375_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n911_), .A2(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n842_), .A2(new_n620_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(KEYINPUT117), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n916_), .A2(new_n662_), .A3(new_n918_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g719(.A1(new_n916_), .A2(new_n680_), .A3(new_n918_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g721(.A1(new_n916_), .A2(new_n374_), .A3(new_n918_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(KEYINPUT61), .B(G155gat), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n923_), .B(new_n924_), .ZN(G1346gat));
  NAND4_X1  g724(.A1(new_n916_), .A2(G162gat), .A3(new_n342_), .A4(new_n918_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n916_), .A2(new_n337_), .A3(new_n918_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  OR3_X1    g728(.A1(new_n929_), .A2(KEYINPUT118), .A3(G162gat), .ZN(new_n930_));
  OAI21_X1  g729(.A(KEYINPUT118), .B1(new_n929_), .B2(G162gat), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n927_), .B1(new_n930_), .B2(new_n931_), .ZN(G1347gat));
  INV_X1    g731(.A(KEYINPUT119), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n735_), .A2(new_n669_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n642_), .A2(new_n643_), .ZN(new_n935_));
  OAI211_X1 g734(.A(new_n934_), .B(new_n935_), .C1(new_n872_), .C2(new_n887_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n933_), .B1(new_n936_), .B2(new_n665_), .ZN(new_n937_));
  INV_X1    g736(.A(new_n934_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n938_), .B1(new_n911_), .B2(new_n915_), .ZN(new_n939_));
  NAND4_X1  g738(.A1(new_n939_), .A2(KEYINPUT119), .A3(new_n662_), .A4(new_n935_), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n937_), .A2(new_n940_), .A3(G169gat), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(KEYINPUT121), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT121), .ZN(new_n943_));
  NAND4_X1  g742(.A1(new_n937_), .A2(new_n940_), .A3(new_n943_), .A4(G169gat), .ZN(new_n944_));
  XOR2_X1   g743(.A(KEYINPUT120), .B(KEYINPUT62), .Z(new_n945_));
  NAND3_X1  g744(.A1(new_n942_), .A2(new_n944_), .A3(new_n945_), .ZN(new_n946_));
  INV_X1    g745(.A(KEYINPUT122), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n939_), .A2(new_n947_), .A3(new_n935_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n936_), .A2(KEYINPUT122), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n948_), .A2(new_n949_), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n950_), .A2(new_n662_), .A3(new_n440_), .ZN(new_n951_));
  INV_X1    g750(.A(new_n945_), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n941_), .A2(KEYINPUT121), .A3(new_n952_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n946_), .A2(new_n951_), .A3(new_n953_), .ZN(G1348gat));
  NAND4_X1  g753(.A1(new_n939_), .A2(G176gat), .A3(new_n680_), .A4(new_n935_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n955_), .B(KEYINPUT123), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n950_), .A2(new_n680_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n956_), .B1(new_n439_), .B2(new_n957_), .ZN(G1349gat));
  INV_X1    g757(.A(KEYINPUT124), .ZN(new_n959_));
  AOI211_X1 g758(.A(new_n410_), .B(new_n375_), .C1(new_n948_), .C2(new_n949_), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n939_), .A2(new_n374_), .A3(new_n935_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n961_), .A2(new_n436_), .ZN(new_n962_));
  INV_X1    g761(.A(new_n962_), .ZN(new_n963_));
  OAI21_X1  g762(.A(new_n959_), .B1(new_n960_), .B2(new_n963_), .ZN(new_n964_));
  NAND3_X1  g763(.A1(new_n950_), .A2(new_n411_), .A3(new_n374_), .ZN(new_n965_));
  NAND3_X1  g764(.A1(new_n965_), .A2(KEYINPUT124), .A3(new_n962_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n964_), .A2(new_n966_), .ZN(G1350gat));
  AND2_X1   g766(.A1(new_n414_), .A2(new_n415_), .ZN(new_n968_));
  INV_X1    g767(.A(new_n968_), .ZN(new_n969_));
  NAND3_X1  g768(.A1(new_n950_), .A2(new_n969_), .A3(new_n337_), .ZN(new_n970_));
  AOI21_X1  g769(.A(new_n341_), .B1(new_n948_), .B2(new_n949_), .ZN(new_n971_));
  OAI21_X1  g770(.A(new_n970_), .B1(new_n971_), .B2(new_n437_), .ZN(G1351gat));
  NAND2_X1  g771(.A1(new_n939_), .A2(new_n620_), .ZN(new_n973_));
  INV_X1    g772(.A(new_n973_), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n974_), .A2(new_n662_), .ZN(new_n975_));
  OR2_X1    g774(.A1(new_n384_), .A2(KEYINPUT125), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n384_), .A2(KEYINPUT125), .ZN(new_n977_));
  NAND3_X1  g776(.A1(new_n975_), .A2(new_n976_), .A3(new_n977_), .ZN(new_n978_));
  OAI21_X1  g777(.A(new_n978_), .B1(new_n975_), .B2(new_n977_), .ZN(G1352gat));
  NOR2_X1   g778(.A1(new_n973_), .A2(new_n274_), .ZN(new_n980_));
  XNOR2_X1  g779(.A(KEYINPUT126), .B(G204gat), .ZN(new_n981_));
  XNOR2_X1  g780(.A(new_n980_), .B(new_n981_), .ZN(G1353gat));
  AOI21_X1  g781(.A(new_n375_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n983_));
  NAND2_X1  g782(.A1(new_n983_), .A2(KEYINPUT127), .ZN(new_n984_));
  INV_X1    g783(.A(new_n984_), .ZN(new_n985_));
  NOR2_X1   g784(.A1(new_n983_), .A2(KEYINPUT127), .ZN(new_n986_));
  NOR3_X1   g785(.A1(new_n973_), .A2(new_n985_), .A3(new_n986_), .ZN(new_n987_));
  NOR2_X1   g786(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n988_));
  XNOR2_X1  g787(.A(new_n987_), .B(new_n988_), .ZN(G1354gat));
  INV_X1    g788(.A(G218gat), .ZN(new_n990_));
  NOR3_X1   g789(.A1(new_n973_), .A2(new_n990_), .A3(new_n341_), .ZN(new_n991_));
  NAND2_X1  g790(.A1(new_n974_), .A2(new_n337_), .ZN(new_n992_));
  AOI21_X1  g791(.A(new_n991_), .B1(new_n990_), .B2(new_n992_), .ZN(G1355gat));
endmodule


