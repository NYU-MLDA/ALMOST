//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 0 1 1 0 1 1 1 0 0 0 0 0 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n855_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n920_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT70), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT11), .ZN(new_n205_));
  XOR2_X1   g004(.A(G71gat), .B(G78gat), .Z(new_n206_));
  OR2_X1    g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n202_), .B(KEYINPUT70), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT11), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n205_), .A2(new_n210_), .A3(new_n206_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n207_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT6), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G99gat), .A3(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G99gat), .ZN(new_n219_));
  INV_X1    g018(.A(G106gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT7), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n218_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n224_));
  AOI21_X1  g023(.A(KEYINPUT7), .B1(new_n221_), .B2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n219_), .A2(new_n220_), .A3(KEYINPUT66), .ZN(new_n226_));
  AOI21_X1  g025(.A(KEYINPUT67), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n224_), .B1(G99gat), .B2(G106gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT7), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n226_), .A2(new_n228_), .A3(KEYINPUT67), .A4(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n223_), .B1(new_n227_), .B2(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(G85gat), .B(G92gat), .Z(new_n233_));
  INV_X1    g032(.A(KEYINPUT8), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n232_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n233_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n215_), .A2(new_n217_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(new_n222_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n239_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n226_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(new_n230_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n238_), .B1(new_n243_), .B2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n237_), .B1(new_n248_), .B2(new_n234_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n233_), .A2(KEYINPUT9), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT9), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n251_), .A2(G85gat), .A3(G92gat), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n250_), .A2(new_n252_), .A3(new_n218_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  OR2_X1    g053(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT64), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT64), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n255_), .A2(new_n259_), .A3(new_n256_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  AND3_X1   g060(.A1(new_n261_), .A2(KEYINPUT65), .A3(new_n220_), .ZN(new_n262_));
  AOI21_X1  g061(.A(KEYINPUT65), .B1(new_n261_), .B2(new_n220_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n254_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n249_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n213_), .A2(new_n265_), .A3(KEYINPUT12), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n235_), .B1(new_n247_), .B2(new_n223_), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n246_), .A2(new_n230_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n242_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n269_), .A2(new_n240_), .A3(new_n222_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n233_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n267_), .B1(new_n271_), .B2(KEYINPUT8), .ZN(new_n272_));
  INV_X1    g071(.A(new_n263_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n261_), .A2(KEYINPUT65), .A3(new_n220_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n253_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT69), .B1(new_n272_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n249_), .A2(new_n277_), .A3(new_n264_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n276_), .A2(new_n278_), .A3(new_n212_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G230gat), .A2(G233gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n212_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n284_));
  NOR3_X1   g083(.A1(new_n283_), .A2(new_n284_), .A3(KEYINPUT12), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n249_), .A2(new_n277_), .A3(new_n264_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n277_), .B1(new_n249_), .B2(new_n264_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n213_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT12), .ZN(new_n289_));
  AOI21_X1  g088(.A(KEYINPUT72), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  OAI211_X1 g089(.A(new_n266_), .B(new_n282_), .C1(new_n285_), .C2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT73), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n284_), .B1(new_n283_), .B2(KEYINPUT12), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n288_), .A2(KEYINPUT72), .A3(new_n289_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n296_), .A2(KEYINPUT73), .A3(new_n266_), .A4(new_n282_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n288_), .A2(new_n279_), .A3(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n280_), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n299_), .B(new_n300_), .C1(new_n298_), .C2(new_n288_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n293_), .A2(new_n297_), .A3(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G120gat), .B(G148gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT5), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G176gat), .B(G204gat), .ZN(new_n305_));
  XOR2_X1   g104(.A(new_n304_), .B(new_n305_), .Z(new_n306_));
  NAND2_X1  g105(.A1(new_n302_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n306_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n293_), .A2(new_n297_), .A3(new_n301_), .A4(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(KEYINPUT74), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT74), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n302_), .A2(new_n311_), .A3(new_n306_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT13), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT75), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n313_), .A2(new_n314_), .ZN(new_n318_));
  AOI21_X1  g117(.A(KEYINPUT13), .B1(new_n310_), .B2(new_n312_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT75), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n317_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  XOR2_X1   g122(.A(G29gat), .B(G36gat), .Z(new_n324_));
  XOR2_X1   g123(.A(G43gat), .B(G50gat), .Z(new_n325_));
  XOR2_X1   g124(.A(new_n324_), .B(new_n325_), .Z(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT15), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n327_), .B1(new_n264_), .B2(new_n249_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT35), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G232gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT34), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n328_), .B1(new_n329_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n326_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n276_), .A2(new_n278_), .A3(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n332_), .A2(new_n329_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n333_), .B(new_n335_), .C1(new_n329_), .C2(new_n332_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G190gat), .B(G218gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G134gat), .B(G162gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n342_), .A2(KEYINPUT36), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n338_), .A2(new_n339_), .A3(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT76), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n338_), .A2(new_n339_), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n342_), .B(KEYINPUT36), .Z(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n345_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT77), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n349_), .A2(KEYINPUT37), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(KEYINPUT37), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n353_), .A2(new_n345_), .A3(new_n348_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G231gat), .A2(G233gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n212_), .B(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G1gat), .B(G8gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT78), .ZN(new_n359_));
  INV_X1    g158(.A(G15gat), .ZN(new_n360_));
  INV_X1    g159(.A(G22gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G15gat), .A2(G22gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G1gat), .A2(G8gat), .ZN(new_n364_));
  AOI22_X1  g163(.A1(new_n362_), .A2(new_n363_), .B1(KEYINPUT14), .B2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n359_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n357_), .B(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(G127gat), .B(G155gat), .Z(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT16), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G183gat), .B(G211gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT17), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n371_), .A2(new_n372_), .ZN(new_n374_));
  NOR3_X1   g173(.A1(new_n367_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n367_), .A2(new_n373_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT79), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n355_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G141gat), .A2(G148gat), .ZN(new_n381_));
  AND2_X1   g180(.A1(KEYINPUT88), .A2(KEYINPUT2), .ZN(new_n382_));
  NOR2_X1   g181(.A1(KEYINPUT88), .A2(KEYINPUT2), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n381_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT89), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(G141gat), .A2(G148gat), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT2), .ZN(new_n389_));
  OAI22_X1  g188(.A1(new_n387_), .A2(new_n388_), .B1(new_n381_), .B2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n390_), .B1(new_n388_), .B2(new_n387_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n386_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT86), .ZN(new_n393_));
  INV_X1    g192(.A(G155gat), .ZN(new_n394_));
  INV_X1    g193(.A(G162gat), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n393_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT86), .B1(G155gat), .B2(G162gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n394_), .A2(new_n395_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n392_), .A2(new_n398_), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT1), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n398_), .B1(new_n402_), .B2(new_n399_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT87), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  OAI22_X1  g204(.A1(new_n403_), .A2(KEYINPUT87), .B1(KEYINPUT1), .B2(new_n400_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n387_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n381_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n401_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  XOR2_X1   g209(.A(G127gat), .B(G134gat), .Z(new_n411_));
  XNOR2_X1  g210(.A(G113gat), .B(G120gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n410_), .B(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G225gat), .A2(G233gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT96), .B(KEYINPUT4), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n410_), .A2(new_n413_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n416_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT4), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n419_), .B(new_n420_), .C1(new_n414_), .C2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n417_), .A2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G1gat), .B(G29gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(G85gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT0), .B(G57gat), .ZN(new_n426_));
  XOR2_X1   g225(.A(new_n425_), .B(new_n426_), .Z(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n423_), .A2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n417_), .A2(new_n422_), .A3(new_n427_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT27), .ZN(new_n433_));
  INV_X1    g232(.A(G169gat), .ZN(new_n434_));
  INV_X1    g233(.A(G176gat), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n434_), .A2(new_n435_), .A3(KEYINPUT84), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT84), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n437_), .B1(G169gat), .B2(G176gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT24), .B1(new_n434_), .B2(new_n435_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT85), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G183gat), .A2(G190gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT23), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT25), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(G183gat), .ZN(new_n446_));
  XOR2_X1   g245(.A(new_n446_), .B(KEYINPUT83), .Z(new_n447_));
  XNOR2_X1  g246(.A(KEYINPUT26), .B(G190gat), .ZN(new_n448_));
  INV_X1    g247(.A(G183gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT25), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT82), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n448_), .A2(new_n451_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n447_), .B(new_n452_), .C1(KEYINPUT82), .C2(new_n450_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT24), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n439_), .A2(new_n454_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n442_), .A2(new_n444_), .A3(new_n453_), .A4(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G197gat), .B(G204gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT91), .ZN(new_n458_));
  INV_X1    g257(.A(G197gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(G204gat), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n458_), .B(KEYINPUT21), .C1(KEYINPUT91), .C2(new_n460_), .ZN(new_n461_));
  XOR2_X1   g260(.A(G211gat), .B(G218gat), .Z(new_n462_));
  INV_X1    g261(.A(KEYINPUT21), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n462_), .B1(new_n463_), .B2(new_n457_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n461_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n457_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(new_n462_), .A3(KEYINPUT21), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n444_), .B1(G183gat), .B2(G190gat), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT22), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n471_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n472_));
  OAI21_X1  g271(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n470_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n456_), .A2(new_n469_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT20), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n474_), .A2(KEYINPUT94), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n470_), .A2(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n474_), .A2(KEYINPUT94), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n446_), .A2(new_n450_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n448_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n454_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(new_n444_), .A3(new_n484_), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n440_), .A2(KEYINPUT93), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n440_), .A2(KEYINPUT93), .ZN(new_n487_));
  NOR3_X1   g286(.A1(new_n486_), .A2(new_n487_), .A3(new_n439_), .ZN(new_n488_));
  OAI22_X1  g287(.A1(new_n480_), .A2(new_n481_), .B1(new_n485_), .B2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n478_), .B1(new_n489_), .B2(new_n468_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n477_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G226gat), .A2(G233gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT19), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT20), .B1(new_n489_), .B2(new_n468_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n495_), .A2(new_n493_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n456_), .A2(new_n476_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(new_n468_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G8gat), .B(G36gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT18), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G64gat), .B(G92gat), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n501_), .B(new_n502_), .Z(new_n503_));
  NAND3_X1  g302(.A1(new_n494_), .A2(new_n499_), .A3(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT101), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n495_), .A2(KEYINPUT100), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n498_), .A2(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n495_), .A2(KEYINPUT100), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n493_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n491_), .A2(new_n493_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n503_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n433_), .B1(new_n505_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n504_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n503_), .B1(new_n494_), .B2(new_n499_), .ZN(new_n516_));
  NOR3_X1   g315(.A1(new_n515_), .A2(KEYINPUT27), .A3(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n432_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n520_));
  INV_X1    g319(.A(G228gat), .ZN(new_n521_));
  INV_X1    g320(.A(G233gat), .ZN(new_n522_));
  NOR3_X1   g321(.A1(new_n521_), .A2(new_n522_), .A3(KEYINPUT92), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n520_), .B(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n381_), .B(new_n408_), .C1(new_n405_), .C2(new_n406_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n526_), .A2(new_n401_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT29), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n468_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(G78gat), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n521_), .A2(new_n522_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT92), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n529_), .A2(new_n530_), .A3(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n469_), .B1(new_n410_), .B2(KEYINPUT29), .ZN(new_n536_));
  OAI21_X1  g335(.A(G78gat), .B1(new_n536_), .B2(new_n533_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n535_), .A2(new_n537_), .A3(G106gat), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(G106gat), .B1(new_n535_), .B2(new_n537_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n527_), .A2(new_n528_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G22gat), .B(G50gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  NOR3_X1   g342(.A1(new_n539_), .A2(new_n540_), .A3(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n543_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n535_), .A2(new_n537_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n220_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n545_), .B1(new_n547_), .B2(new_n538_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n525_), .B1(new_n544_), .B2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G71gat), .B(G99gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(G43gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n497_), .B(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(new_n413_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G227gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(new_n360_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT30), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT31), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n553_), .A2(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n553_), .A2(new_n557_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n543_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n547_), .A2(new_n538_), .A3(new_n545_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n561_), .A2(new_n562_), .A3(new_n524_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n549_), .A2(new_n560_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n560_), .B1(new_n549_), .B2(new_n563_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n519_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n558_), .A2(new_n559_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n568_), .A2(new_n549_), .A3(new_n563_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n494_), .A2(new_n499_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT99), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n503_), .A2(KEYINPUT32), .ZN(new_n573_));
  NOR3_X1   g372(.A1(new_n571_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n509_), .B(new_n510_), .C1(new_n571_), .C2(KEYINPUT99), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n574_), .B1(new_n575_), .B2(new_n573_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n431_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n430_), .A2(KEYINPUT97), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT97), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n417_), .A2(new_n422_), .A3(new_n579_), .A4(new_n427_), .ZN(new_n580_));
  XOR2_X1   g379(.A(KEYINPUT98), .B(KEYINPUT33), .Z(new_n581_));
  NAND3_X1  g380(.A1(new_n578_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n427_), .B1(new_n415_), .B2(new_n420_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n419_), .B1(new_n414_), .B2(new_n421_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n584_), .B1(new_n585_), .B2(new_n420_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n417_), .A2(new_n422_), .A3(KEYINPUT33), .A4(new_n427_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n516_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n588_), .A2(new_n504_), .A3(KEYINPUT95), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT95), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n590_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n586_), .A2(new_n587_), .A3(new_n589_), .A4(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n577_), .B1(new_n583_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n570_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n567_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n366_), .B(new_n334_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G229gat), .A2(G233gat), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT80), .Z(new_n600_));
  OR2_X1    g399(.A1(new_n327_), .A2(new_n366_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n366_), .A2(new_n334_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n601_), .A2(new_n602_), .A3(new_n597_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n600_), .A2(new_n603_), .ZN(new_n604_));
  XOR2_X1   g403(.A(G113gat), .B(G141gat), .Z(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT81), .ZN(new_n606_));
  XOR2_X1   g405(.A(G169gat), .B(G197gat), .Z(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n604_), .B(new_n608_), .Z(new_n609_));
  NAND2_X1  g408(.A1(new_n595_), .A2(new_n609_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n323_), .A2(new_n380_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(G1gat), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n431_), .B(KEYINPUT102), .Z(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n611_), .A2(new_n612_), .A3(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT103), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT38), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n615_), .A2(KEYINPUT103), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n615_), .A2(KEYINPUT103), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(KEYINPUT38), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n609_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n320_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n595_), .A2(new_n349_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n377_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n623_), .A2(new_n626_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n627_), .A2(KEYINPUT104), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(KEYINPUT104), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(new_n431_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(G1gat), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n618_), .A2(new_n621_), .A3(new_n632_), .ZN(G1324gat));
  NOR2_X1   g432(.A1(new_n514_), .A2(new_n517_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(G8gat), .B1(new_n627_), .B2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT39), .ZN(new_n637_));
  INV_X1    g436(.A(G8gat), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n611_), .A2(new_n638_), .A3(new_n634_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g440(.A(KEYINPUT41), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n568_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n643_));
  OAI21_X1  g442(.A(KEYINPUT105), .B1(new_n643_), .B2(new_n360_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n643_), .A2(KEYINPUT105), .A3(new_n360_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n642_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n646_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n648_), .A2(KEYINPUT41), .A3(new_n644_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n611_), .A2(new_n360_), .A3(new_n560_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n647_), .A2(new_n649_), .A3(new_n650_), .ZN(G1326gat));
  INV_X1    g450(.A(new_n563_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n524_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n654_), .A2(KEYINPUT106), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(KEYINPUT106), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n361_), .B1(new_n630_), .B2(new_n657_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT42), .Z(new_n659_));
  NAND3_X1  g458(.A1(new_n611_), .A2(new_n361_), .A3(new_n657_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1327gat));
  INV_X1    g460(.A(new_n349_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(new_n378_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT111), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n664_), .A2(new_n320_), .A3(new_n610_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  OR3_X1    g465(.A1(new_n666_), .A2(G29gat), .A3(new_n432_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n568_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n518_), .B1(new_n669_), .B2(new_n564_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n592_), .ZN(new_n671_));
  AOI22_X1  g470(.A1(new_n671_), .A2(new_n582_), .B1(new_n576_), .B2(new_n431_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n672_), .A2(new_n569_), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n354_), .B(new_n352_), .C1(new_n670_), .C2(new_n673_), .ZN(new_n674_));
  XOR2_X1   g473(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT108), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT108), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n674_), .A2(new_n678_), .A3(new_n675_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT109), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n680_), .B1(new_n674_), .B2(KEYINPUT43), .ZN(new_n681_));
  INV_X1    g480(.A(new_n355_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n682_), .A2(KEYINPUT109), .A3(new_n595_), .A4(new_n683_), .ZN(new_n684_));
  AOI22_X1  g483(.A1(new_n677_), .A2(new_n679_), .B1(new_n681_), .B2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n315_), .A2(new_n378_), .A3(new_n609_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n668_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n669_), .A2(new_n564_), .ZN(new_n688_));
  AOI22_X1  g487(.A1(new_n688_), .A2(new_n519_), .B1(new_n570_), .B2(new_n593_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n689_), .A2(new_n355_), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT109), .B1(new_n690_), .B2(new_n683_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n674_), .A2(new_n680_), .A3(KEYINPUT43), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n674_), .A2(new_n678_), .A3(new_n675_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n678_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n694_));
  OAI22_X1  g493(.A1(new_n691_), .A2(new_n692_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n686_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n695_), .A2(KEYINPUT44), .A3(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n687_), .A2(new_n697_), .A3(new_n614_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n698_), .A2(KEYINPUT110), .ZN(new_n699_));
  OAI21_X1  g498(.A(G29gat), .B1(new_n698_), .B2(KEYINPUT110), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n667_), .B1(new_n699_), .B2(new_n700_), .ZN(G1328gat));
  NOR2_X1   g500(.A1(new_n635_), .A2(G36gat), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(KEYINPUT113), .B1(new_n666_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT113), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n665_), .A2(new_n705_), .A3(new_n702_), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n704_), .A2(KEYINPUT45), .A3(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(KEYINPUT45), .B1(new_n704_), .B2(new_n706_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n687_), .A2(new_n697_), .A3(new_n634_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT112), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n687_), .A2(new_n697_), .A3(KEYINPUT112), .A4(new_n634_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(G36gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n709_), .B1(new_n712_), .B2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(KEYINPUT114), .B(KEYINPUT46), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n709_), .B(new_n716_), .C1(new_n712_), .C2(new_n714_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1329gat));
  NAND4_X1  g519(.A1(new_n687_), .A2(new_n697_), .A3(G43gat), .A4(new_n560_), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n721_), .A2(KEYINPUT115), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n665_), .A2(new_n560_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n721_), .B(KEYINPUT115), .C1(G43gat), .C2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n722_), .A2(new_n725_), .A3(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n722_), .B2(new_n725_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1330gat));
  INV_X1    g528(.A(new_n654_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n687_), .A2(new_n697_), .A3(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(G50gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(G50gat), .B1(new_n655_), .B2(new_n656_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT116), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n732_), .B1(new_n666_), .B2(new_n734_), .ZN(G1331gat));
  NAND2_X1  g534(.A1(new_n595_), .A2(new_n622_), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n315_), .A2(new_n736_), .A3(new_n380_), .ZN(new_n737_));
  INV_X1    g536(.A(G57gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n737_), .A2(new_n738_), .A3(new_n614_), .ZN(new_n739_));
  NOR4_X1   g538(.A1(new_n322_), .A2(new_n378_), .A3(new_n609_), .A4(new_n624_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n740_), .A2(new_n431_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n739_), .B1(new_n741_), .B2(new_n738_), .ZN(G1332gat));
  INV_X1    g541(.A(G64gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n740_), .B2(new_n634_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(KEYINPUT117), .B(KEYINPUT48), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n744_), .B(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n737_), .A2(new_n743_), .A3(new_n634_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1333gat));
  INV_X1    g547(.A(G71gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n740_), .B2(new_n560_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT49), .Z(new_n751_));
  NAND3_X1  g550(.A1(new_n737_), .A2(new_n749_), .A3(new_n560_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1334gat));
  AOI21_X1  g552(.A(new_n530_), .B1(new_n740_), .B2(new_n657_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT50), .Z(new_n755_));
  NAND3_X1  g554(.A1(new_n737_), .A2(new_n530_), .A3(new_n657_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1335gat));
  NOR3_X1   g556(.A1(new_n322_), .A2(new_n664_), .A3(new_n736_), .ZN(new_n758_));
  INV_X1    g557(.A(G85gat), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n758_), .A2(new_n759_), .A3(new_n614_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n320_), .A2(new_n378_), .A3(new_n622_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n685_), .A2(new_n432_), .A3(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n760_), .B1(new_n762_), .B2(new_n759_), .ZN(G1336gat));
  AOI21_X1  g562(.A(G92gat), .B1(new_n758_), .B2(new_n634_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT118), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n685_), .A2(new_n761_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n634_), .A2(G92gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n765_), .B1(new_n766_), .B2(new_n767_), .ZN(G1337gat));
  NAND3_X1  g567(.A1(new_n758_), .A2(new_n261_), .A3(new_n560_), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n685_), .A2(new_n568_), .A3(new_n761_), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n769_), .B(KEYINPUT119), .C1(new_n770_), .C2(new_n219_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g571(.A1(new_n758_), .A2(new_n220_), .A3(new_n730_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n220_), .B1(new_n766_), .B2(new_n730_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT52), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n774_), .A2(new_n775_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT53), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n780_), .B(new_n773_), .C1(new_n776_), .C2(new_n777_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1339gat));
  NAND3_X1  g581(.A1(new_n600_), .A2(new_n603_), .A3(new_n608_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n608_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n784_));
  OR2_X1    g583(.A1(new_n784_), .A2(KEYINPUT121), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(KEYINPUT121), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n601_), .A2(new_n602_), .A3(new_n598_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n785_), .A2(new_n786_), .A3(new_n787_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n783_), .A2(new_n788_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n309_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT55), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n293_), .A2(new_n791_), .A3(new_n297_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n266_), .ZN(new_n793_));
  AOI211_X1 g592(.A(new_n793_), .B(new_n281_), .C1(new_n294_), .C2(new_n295_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n266_), .B(new_n279_), .C1(new_n285_), .C2(new_n290_), .ZN(new_n795_));
  AOI22_X1  g594(.A1(new_n794_), .A2(KEYINPUT55), .B1(new_n795_), .B2(new_n300_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n792_), .A2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT56), .B1(new_n797_), .B2(new_n306_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT56), .ZN(new_n799_));
  AOI211_X1 g598(.A(new_n799_), .B(new_n308_), .C1(new_n792_), .C2(new_n796_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n790_), .B1(new_n798_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT58), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  OAI211_X1 g602(.A(KEYINPUT58), .B(new_n790_), .C1(new_n798_), .C2(new_n800_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n803_), .A2(new_n682_), .A3(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT57), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n609_), .A2(new_n309_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n807_), .B1(new_n798_), .B2(new_n800_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n310_), .A2(new_n312_), .A3(new_n789_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n806_), .B1(new_n810_), .B2(new_n349_), .ZN(new_n811_));
  AOI211_X1 g610(.A(KEYINPUT57), .B(new_n662_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n805_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n625_), .ZN(new_n814_));
  AOI211_X1 g613(.A(new_n378_), .B(new_n609_), .C1(new_n352_), .C2(new_n354_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n315_), .A2(new_n815_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(KEYINPUT120), .B(KEYINPUT54), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n315_), .A2(new_n815_), .A3(new_n817_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n814_), .A2(new_n821_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n613_), .A2(new_n634_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n565_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n822_), .A2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(G113gat), .B1(new_n825_), .B2(new_n609_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n813_), .A2(new_n378_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n821_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n824_), .A2(KEYINPUT59), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT59), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n825_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(G113gat), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n834_), .B1(new_n609_), .B2(KEYINPUT122), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n835_), .B1(KEYINPUT122), .B2(new_n834_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n826_), .B1(new_n833_), .B2(new_n836_), .ZN(G1340gat));
  OAI21_X1  g636(.A(G120gat), .B1(new_n832_), .B2(new_n322_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n825_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT60), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(G120gat), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n315_), .A2(KEYINPUT60), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n842_), .B2(G120gat), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n838_), .B1(new_n839_), .B2(new_n843_), .ZN(G1341gat));
  OAI21_X1  g643(.A(G127gat), .B1(new_n832_), .B2(new_n625_), .ZN(new_n845_));
  OR2_X1    g644(.A1(new_n378_), .A2(G127gat), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n845_), .B1(new_n839_), .B2(new_n846_), .ZN(G1342gat));
  AOI21_X1  g646(.A(G134gat), .B1(new_n825_), .B2(new_n662_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n682_), .A2(G134gat), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(KEYINPUT123), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n848_), .B1(new_n833_), .B2(new_n850_), .ZN(G1343gat));
  NOR2_X1   g650(.A1(new_n822_), .A2(new_n669_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n852_), .A2(new_n609_), .A3(new_n823_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g653(.A1(new_n852_), .A2(new_n323_), .A3(new_n823_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g655(.A1(new_n852_), .A2(new_n379_), .A3(new_n823_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(KEYINPUT61), .B(G155gat), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(G1346gat));
  NAND4_X1  g658(.A1(new_n852_), .A2(new_n395_), .A3(new_n662_), .A4(new_n823_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n852_), .A2(new_n682_), .A3(new_n823_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n861_), .B2(new_n395_), .ZN(G1347gat));
  INV_X1    g661(.A(KEYINPUT62), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n614_), .A2(new_n568_), .A3(new_n635_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n864_), .A2(new_n656_), .A3(new_n655_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n865_), .B1(new_n827_), .B2(new_n821_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n866_), .A2(new_n609_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n863_), .B1(new_n867_), .B2(new_n471_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(G169gat), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n434_), .B1(new_n867_), .B2(new_n863_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n868_), .B2(new_n870_), .ZN(G1348gat));
  AOI21_X1  g670(.A(G176gat), .B1(new_n866_), .B2(new_n320_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n822_), .A2(new_n730_), .ZN(new_n873_));
  AND3_X1   g672(.A1(new_n323_), .A2(G176gat), .A3(new_n864_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n872_), .B1(new_n873_), .B2(new_n874_), .ZN(G1349gat));
  NOR2_X1   g674(.A1(new_n625_), .A2(new_n482_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n866_), .A2(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(KEYINPUT124), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n877_), .A2(KEYINPUT124), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n873_), .A2(new_n379_), .A3(new_n864_), .ZN(new_n880_));
  AOI211_X1 g679(.A(new_n878_), .B(new_n879_), .C1(new_n449_), .C2(new_n880_), .ZN(G1350gat));
  NAND3_X1  g680(.A1(new_n866_), .A2(new_n662_), .A3(new_n448_), .ZN(new_n882_));
  INV_X1    g681(.A(G190gat), .ZN(new_n883_));
  AOI211_X1 g682(.A(KEYINPUT125), .B(new_n883_), .C1(new_n866_), .C2(new_n682_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT125), .ZN(new_n885_));
  INV_X1    g684(.A(new_n865_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n609_), .A2(new_n309_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n797_), .A2(new_n306_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n799_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n797_), .A2(KEYINPUT56), .A3(new_n306_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n887_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n809_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n349_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(KEYINPUT57), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n810_), .A2(new_n806_), .A3(new_n349_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n379_), .B1(new_n896_), .B2(new_n805_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n820_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n817_), .B1(new_n315_), .B2(new_n815_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n682_), .B(new_n886_), .C1(new_n897_), .C2(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n885_), .B1(new_n901_), .B2(G190gat), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n882_), .B1(new_n884_), .B2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT126), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  OAI211_X1 g704(.A(KEYINPUT126), .B(new_n882_), .C1(new_n884_), .C2(new_n902_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1351gat));
  NOR2_X1   g706(.A1(new_n635_), .A2(new_n431_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n852_), .A2(new_n609_), .A3(new_n908_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g709(.A1(new_n852_), .A2(new_n323_), .A3(new_n908_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G204gat), .ZN(G1353gat));
  XNOR2_X1  g711(.A(KEYINPUT63), .B(G211gat), .ZN(new_n913_));
  OR2_X1    g712(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n852_), .A2(new_n377_), .A3(new_n908_), .ZN(new_n915_));
  MUX2_X1   g714(.A(new_n913_), .B(new_n914_), .S(new_n915_), .Z(G1354gat));
  AND2_X1   g715(.A1(new_n852_), .A2(new_n908_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n662_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(KEYINPUT127), .B(G218gat), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n355_), .A2(new_n919_), .ZN(new_n920_));
  AOI22_X1  g719(.A1(new_n918_), .A2(new_n919_), .B1(new_n917_), .B2(new_n920_), .ZN(G1355gat));
endmodule


