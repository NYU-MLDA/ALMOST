//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1 1 1 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 0 0 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n833_, new_n834_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_;
  INV_X1    g000(.A(KEYINPUT97), .ZN(new_n202_));
  OR2_X1    g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(KEYINPUT24), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205_));
  AND3_X1   g004(.A1(new_n203_), .A2(KEYINPUT24), .A3(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT25), .B(G183gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT26), .B(G190gat), .ZN(new_n208_));
  AOI211_X1 g007(.A(new_n204_), .B(new_n206_), .C1(new_n207_), .C2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT23), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(KEYINPUT80), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n211_), .B1(new_n212_), .B2(KEYINPUT23), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n209_), .A2(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT80), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n210_), .B(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n215_), .B1(new_n217_), .B2(KEYINPUT23), .ZN(new_n218_));
  INV_X1    g017(.A(G183gat), .ZN(new_n219_));
  INV_X1    g018(.A(G190gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n218_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(G176gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT22), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT81), .B1(new_n224_), .B2(G169gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT22), .B(G169gat), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n223_), .B(new_n225_), .C1(new_n226_), .C2(KEYINPUT81), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n222_), .A2(new_n205_), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n214_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G71gat), .B(G99gat), .ZN(new_n230_));
  INV_X1    g029(.A(G43gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n229_), .B(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G127gat), .B(G134gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT82), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G113gat), .B(G120gat), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n235_), .A2(new_n237_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n234_), .A2(KEYINPUT82), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n234_), .A2(KEYINPUT82), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n240_), .A3(new_n236_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n233_), .B(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G227gat), .A2(G233gat), .ZN(new_n244_));
  INV_X1    g043(.A(G15gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT30), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT31), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n243_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n243_), .A2(new_n248_), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G155gat), .A2(G162gat), .ZN(new_n252_));
  NOR2_X1   g051(.A1(G155gat), .A2(G162gat), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(G141gat), .A2(G148gat), .ZN(new_n255_));
  XOR2_X1   g054(.A(new_n255_), .B(KEYINPUT3), .Z(new_n256_));
  NAND2_X1  g055(.A1(G141gat), .A2(G148gat), .ZN(new_n257_));
  XOR2_X1   g056(.A(new_n257_), .B(KEYINPUT2), .Z(new_n258_));
  OAI211_X1 g057(.A(new_n252_), .B(new_n254_), .C1(new_n256_), .C2(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n253_), .B1(KEYINPUT1), .B2(new_n252_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n260_), .B1(KEYINPUT1), .B2(new_n252_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n255_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n261_), .A2(new_n262_), .A3(new_n257_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n259_), .A2(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n264_), .A2(KEYINPUT29), .ZN(new_n265_));
  XOR2_X1   g064(.A(KEYINPUT83), .B(KEYINPUT28), .Z(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G228gat), .A2(G233gat), .ZN(new_n268_));
  INV_X1    g067(.A(G78gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(G106gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n267_), .B(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G211gat), .B(G218gat), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(G197gat), .B(G204gat), .Z(new_n275_));
  NAND3_X1  g074(.A1(new_n274_), .A2(KEYINPUT21), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(G197gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n277_), .A2(KEYINPUT84), .A3(G204gat), .ZN(new_n278_));
  OAI211_X1 g077(.A(KEYINPUT21), .B(new_n278_), .C1(new_n275_), .C2(KEYINPUT84), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n273_), .B1(new_n275_), .B2(KEYINPUT21), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n276_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n283_), .B1(new_n264_), .B2(KEYINPUT29), .ZN(new_n284_));
  XOR2_X1   g083(.A(G22gat), .B(G50gat), .Z(new_n285_));
  XOR2_X1   g084(.A(new_n284_), .B(new_n285_), .Z(new_n286_));
  OR2_X1    g085(.A1(new_n272_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n272_), .A2(new_n286_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT20), .B1(new_n229_), .B2(new_n282_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n209_), .A2(new_n218_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n226_), .A2(new_n223_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n205_), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n294_), .A2(KEYINPUT85), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT86), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n213_), .A2(new_n296_), .A3(new_n221_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n294_), .A2(KEYINPUT85), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n295_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n296_), .B1(new_n213_), .B2(new_n221_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n292_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n282_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT87), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT87), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n301_), .A2(new_n304_), .A3(new_n282_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n291_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G226gat), .A2(G233gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT19), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT88), .B1(new_n306_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n229_), .A2(new_n282_), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n311_), .B(KEYINPUT20), .C1(new_n301_), .C2(new_n282_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n312_), .A2(new_n308_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n291_), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n301_), .A2(new_n304_), .A3(new_n282_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n304_), .B1(new_n301_), .B2(new_n282_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n314_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT88), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n317_), .A2(new_n318_), .A3(new_n308_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G8gat), .B(G36gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT18), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G64gat), .B(G92gat), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n321_), .B(new_n322_), .Z(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT32), .ZN(new_n324_));
  AND4_X1   g123(.A1(new_n310_), .A2(new_n313_), .A3(new_n319_), .A4(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n242_), .A2(new_n264_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n238_), .A2(new_n259_), .A3(new_n241_), .A4(new_n263_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n326_), .A2(KEYINPUT4), .A3(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G225gat), .A2(G233gat), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT4), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n242_), .A2(new_n264_), .A3(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n328_), .A2(new_n330_), .A3(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n326_), .A2(new_n329_), .A3(new_n327_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT90), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n326_), .A2(KEYINPUT90), .A3(new_n329_), .A4(new_n327_), .ZN(new_n337_));
  AND3_X1   g136(.A1(new_n333_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G1gat), .B(G29gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT89), .B(KEYINPUT0), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G57gat), .B(G85gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n338_), .A2(KEYINPUT94), .A3(new_n343_), .ZN(new_n344_));
  NAND4_X1  g143(.A1(new_n333_), .A2(new_n336_), .A3(new_n343_), .A4(new_n337_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT94), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n333_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n343_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n344_), .A2(new_n347_), .A3(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n312_), .A2(new_n308_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n352_), .B1(new_n317_), .B2(new_n308_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n324_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n351_), .A2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n325_), .A2(new_n356_), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n326_), .A2(new_n327_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n343_), .B1(new_n358_), .B2(new_n330_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n328_), .A2(new_n329_), .A3(new_n332_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT92), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n360_), .A2(new_n361_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n359_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT33), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n338_), .A2(KEYINPUT91), .A3(KEYINPUT33), .A4(new_n343_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT91), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT33), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n367_), .B1(new_n345_), .B2(new_n368_), .ZN(new_n369_));
  AOI22_X1  g168(.A1(new_n365_), .A2(new_n345_), .B1(new_n366_), .B2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n310_), .A2(new_n313_), .A3(new_n319_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n323_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n310_), .A2(new_n323_), .A3(new_n313_), .A4(new_n319_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n370_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n357_), .B1(new_n375_), .B2(KEYINPUT93), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT93), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n370_), .A2(new_n373_), .A3(new_n377_), .A4(new_n374_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n290_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n379_));
  XOR2_X1   g178(.A(KEYINPUT95), .B(KEYINPUT27), .Z(new_n380_));
  AOI21_X1  g179(.A(new_n380_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n353_), .A2(new_n372_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n374_), .A2(KEYINPUT27), .A3(new_n382_), .ZN(new_n383_));
  NOR4_X1   g182(.A1(new_n381_), .A2(new_n383_), .A3(new_n289_), .A4(new_n351_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n251_), .B1(new_n379_), .B2(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n251_), .A2(new_n351_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n381_), .A2(new_n383_), .ZN(new_n387_));
  AOI21_X1  g186(.A(KEYINPUT96), .B1(new_n387_), .B2(new_n289_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT96), .ZN(new_n389_));
  NOR4_X1   g188(.A1(new_n381_), .A2(new_n383_), .A3(new_n290_), .A4(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n386_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n385_), .A2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G29gat), .B(G36gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G43gat), .B(G50gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT79), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G15gat), .B(G22gat), .ZN(new_n398_));
  INV_X1    g197(.A(G1gat), .ZN(new_n399_));
  INV_X1    g198(.A(G8gat), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT14), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n398_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G1gat), .B(G8gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n397_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G229gat), .A2(G233gat), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n395_), .B(KEYINPUT15), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n404_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n397_), .B(new_n404_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n406_), .ZN(new_n411_));
  AOI22_X1  g210(.A1(new_n407_), .A2(new_n409_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  XOR2_X1   g211(.A(G113gat), .B(G141gat), .Z(new_n413_));
  XNOR2_X1  g212(.A(G169gat), .B(G197gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  OR2_X1    g214(.A1(new_n412_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n412_), .A2(new_n415_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n202_), .B1(new_n392_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n418_), .ZN(new_n420_));
  AOI211_X1 g219(.A(KEYINPUT97), .B(new_n420_), .C1(new_n385_), .C2(new_n391_), .ZN(new_n421_));
  OR2_X1    g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  XOR2_X1   g221(.A(KEYINPUT10), .B(G99gat), .Z(new_n423_));
  INV_X1    g222(.A(G106gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(G85gat), .B(G92gat), .Z(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT9), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G99gat), .A2(G106gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT6), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT6), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(G99gat), .A3(G106gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(G85gat), .ZN(new_n433_));
  INV_X1    g232(.A(G92gat), .ZN(new_n434_));
  OR3_X1    g233(.A1(new_n433_), .A2(new_n434_), .A3(KEYINPUT9), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n425_), .A2(new_n427_), .A3(new_n432_), .A4(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT7), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT64), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT64), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT7), .ZN(new_n441_));
  NOR2_X1   g240(.A1(G99gat), .A2(G106gat), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n439_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT65), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n439_), .A2(new_n441_), .A3(KEYINPUT65), .A4(new_n442_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT67), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT66), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT66), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT67), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n432_), .A2(new_n453_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n429_), .A2(new_n431_), .A3(new_n450_), .A4(new_n452_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n426_), .B1(new_n448_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT8), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .A4(new_n432_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n426_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n460_), .A2(KEYINPUT8), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n437_), .B1(new_n458_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n395_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT73), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n457_), .A2(KEYINPUT8), .B1(new_n459_), .B2(new_n461_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n408_), .B1(new_n466_), .B2(new_n437_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G232gat), .A2(G233gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT34), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT35), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n464_), .A2(new_n465_), .A3(new_n467_), .A4(new_n472_), .ZN(new_n473_));
  AOI211_X1 g272(.A(new_n471_), .B(new_n470_), .C1(new_n467_), .C2(KEYINPUT73), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n470_), .A2(new_n471_), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n464_), .A2(new_n467_), .A3(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n473_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(G190gat), .B(G218gat), .Z(new_n478_));
  XNOR2_X1  g277(.A(G134gat), .B(G162gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT36), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(new_n482_), .B(KEYINPUT74), .Z(new_n483_));
  NAND2_X1  g282(.A1(new_n477_), .A2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n480_), .B(KEYINPUT36), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n473_), .B(new_n485_), .C1(new_n474_), .C2(new_n476_), .ZN(new_n486_));
  AND3_X1   g285(.A1(new_n484_), .A2(KEYINPUT37), .A3(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n477_), .A2(KEYINPUT75), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT75), .ZN(new_n489_));
  OAI211_X1 g288(.A(new_n489_), .B(new_n473_), .C1(new_n474_), .C2(new_n476_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n491_), .A2(KEYINPUT76), .A3(new_n485_), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT76), .B1(new_n491_), .B2(new_n485_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n484_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT37), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n487_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  XOR2_X1   g295(.A(G127gat), .B(G155gat), .Z(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT16), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G183gat), .B(G211gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT17), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G231gat), .A2(G233gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT77), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n404_), .B(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(G64gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(G57gat), .ZN(new_n507_));
  INV_X1    g306(.A(G57gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(G64gat), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT68), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n507_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n510_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT11), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n508_), .A2(G64gat), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n506_), .A2(G57gat), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT68), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT11), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n507_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n516_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G71gat), .B(G78gat), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n513_), .A2(new_n519_), .A3(new_n521_), .ZN(new_n522_));
  OAI211_X1 g321(.A(KEYINPUT11), .B(new_n520_), .C1(new_n511_), .C2(new_n512_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n502_), .B1(new_n505_), .B2(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n525_), .B1(new_n524_), .B2(new_n505_), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n526_), .B(KEYINPUT78), .Z(new_n527_));
  AND2_X1   g326(.A1(new_n500_), .A2(new_n501_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT69), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n522_), .A2(new_n529_), .A3(new_n523_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n529_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  AOI211_X1 g332(.A(new_n502_), .B(new_n528_), .C1(new_n533_), .C2(new_n505_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n534_), .B1(new_n533_), .B2(new_n505_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n527_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n496_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G230gat), .A2(G233gat), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT70), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n532_), .A2(new_n463_), .A3(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n541_), .B1(new_n532_), .B2(new_n463_), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n458_), .A2(new_n462_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n524_), .A2(KEYINPUT69), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n522_), .A2(new_n529_), .A3(new_n523_), .ZN(new_n547_));
  AOI22_X1  g346(.A1(new_n545_), .A2(new_n436_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n540_), .B1(new_n544_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT12), .ZN(new_n550_));
  OR3_X1    g349(.A1(new_n463_), .A2(new_n550_), .A3(new_n524_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n540_), .B1(new_n532_), .B2(new_n463_), .ZN(new_n552_));
  OAI22_X1  g351(.A1(new_n466_), .A2(new_n437_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT71), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n553_), .A2(new_n554_), .A3(new_n550_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n554_), .B1(new_n553_), .B2(new_n550_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n551_), .B(new_n552_), .C1(new_n555_), .C2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n549_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G120gat), .B(G148gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT5), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G176gat), .B(G204gat), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n560_), .B(new_n561_), .Z(new_n562_));
  NAND2_X1  g361(.A1(new_n558_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n562_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n549_), .A2(new_n557_), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT13), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n563_), .B(new_n565_), .C1(KEYINPUT72), .C2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT72), .B(KEYINPUT13), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n565_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n564_), .B1(new_n549_), .B2(new_n557_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n569_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n567_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n538_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n422_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n351_), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n576_), .A2(G1gat), .A3(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n579_));
  OR2_X1    g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n579_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n573_), .A2(new_n418_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n582_), .A2(new_n536_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n392_), .A2(new_n494_), .A3(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(G1gat), .B1(new_n584_), .B2(new_n577_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n580_), .A2(new_n581_), .A3(new_n585_), .ZN(G1324gat));
  XNOR2_X1  g385(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n584_), .A2(new_n387_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(G8gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT39), .ZN(new_n590_));
  INV_X1    g389(.A(new_n387_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n422_), .A2(new_n400_), .A3(new_n591_), .A4(new_n575_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n587_), .B1(new_n590_), .B2(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n589_), .A2(KEYINPUT39), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT39), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n595_), .B1(new_n588_), .B2(G8gat), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n592_), .B(new_n587_), .C1(new_n594_), .C2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n593_), .A2(new_n598_), .ZN(G1325gat));
  OAI21_X1  g398(.A(G15gat), .B1(new_n584_), .B2(new_n251_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT41), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n600_), .A2(new_n601_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n251_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(new_n245_), .ZN(new_n605_));
  OAI22_X1  g404(.A1(new_n602_), .A2(new_n603_), .B1(new_n576_), .B2(new_n605_), .ZN(G1326gat));
  OAI21_X1  g405(.A(G22gat), .B1(new_n584_), .B2(new_n289_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n607_), .A2(KEYINPUT42), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(KEYINPUT42), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n289_), .A2(G22gat), .ZN(new_n610_));
  OAI22_X1  g409(.A1(new_n608_), .A2(new_n609_), .B1(new_n576_), .B2(new_n610_), .ZN(G1327gat));
  NOR2_X1   g410(.A1(new_n582_), .A2(new_n537_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT43), .ZN(new_n613_));
  INV_X1    g412(.A(new_n496_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n613_), .B1(new_n392_), .B2(new_n614_), .ZN(new_n615_));
  AOI211_X1 g414(.A(KEYINPUT43), .B(new_n496_), .C1(new_n385_), .C2(new_n391_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n612_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT44), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  OAI211_X1 g418(.A(KEYINPUT44), .B(new_n612_), .C1(new_n615_), .C2(new_n616_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(new_n351_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(G29gat), .ZN(new_n622_));
  NOR3_X1   g421(.A1(new_n574_), .A2(new_n537_), .A3(new_n494_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n422_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(G29gat), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n624_), .A2(new_n625_), .A3(new_n351_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n622_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT100), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT100), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n622_), .A2(new_n626_), .A3(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(G1328gat));
  NAND3_X1  g430(.A1(new_n619_), .A2(new_n591_), .A3(new_n620_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(G36gat), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n387_), .A2(G36gat), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n623_), .B(new_n634_), .C1(new_n419_), .C2(new_n421_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT45), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n633_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT46), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n633_), .A2(new_n636_), .A3(KEYINPUT46), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1329gat));
  NAND4_X1  g440(.A1(new_n619_), .A2(G43gat), .A3(new_n604_), .A4(new_n620_), .ZN(new_n642_));
  OAI211_X1 g441(.A(new_n604_), .B(new_n623_), .C1(new_n419_), .C2(new_n421_), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n643_), .A2(KEYINPUT101), .A3(new_n231_), .ZN(new_n644_));
  AOI21_X1  g443(.A(KEYINPUT101), .B1(new_n643_), .B2(new_n231_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n642_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g446(.A1(new_n619_), .A2(new_n290_), .A3(new_n620_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(G50gat), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n289_), .A2(G50gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT102), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n624_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n649_), .A2(new_n652_), .ZN(G1331gat));
  NAND3_X1  g452(.A1(new_n420_), .A2(new_n527_), .A3(new_n535_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n392_), .A2(new_n574_), .A3(new_n494_), .A4(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(KEYINPUT103), .B(G57gat), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n351_), .A2(new_n657_), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n659_), .A2(KEYINPUT104), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(KEYINPUT104), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n418_), .B1(new_n385_), .B2(new_n391_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n538_), .A2(new_n573_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(G57gat), .B1(new_n665_), .B2(new_n351_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n660_), .A2(new_n661_), .A3(new_n666_), .ZN(G1332gat));
  NAND3_X1  g466(.A1(new_n665_), .A2(new_n506_), .A3(new_n591_), .ZN(new_n668_));
  OAI21_X1  g467(.A(G64gat), .B1(new_n656_), .B2(new_n387_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n669_), .A2(KEYINPUT48), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(KEYINPUT48), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n668_), .B1(new_n670_), .B2(new_n671_), .ZN(G1333gat));
  OR3_X1    g471(.A1(new_n664_), .A2(G71gat), .A3(new_n251_), .ZN(new_n673_));
  OAI21_X1  g472(.A(G71gat), .B1(new_n656_), .B2(new_n251_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n674_), .A2(KEYINPUT49), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n674_), .A2(KEYINPUT49), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n673_), .B1(new_n675_), .B2(new_n676_), .ZN(G1334gat));
  NAND3_X1  g476(.A1(new_n665_), .A2(new_n269_), .A3(new_n290_), .ZN(new_n678_));
  OAI21_X1  g477(.A(G78gat), .B1(new_n656_), .B2(new_n289_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n679_), .A2(KEYINPUT50), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n679_), .A2(KEYINPUT50), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n678_), .B1(new_n680_), .B2(new_n681_), .ZN(G1335gat));
  INV_X1    g481(.A(new_n494_), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n662_), .A2(new_n574_), .A3(new_n536_), .A4(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n433_), .B1(new_n684_), .B2(new_n577_), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n685_), .A2(KEYINPUT105), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(KEYINPUT105), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n615_), .A2(new_n616_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n573_), .A2(new_n418_), .A3(new_n537_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n577_), .A2(new_n433_), .ZN(new_n691_));
  AOI22_X1  g490(.A1(new_n686_), .A2(new_n687_), .B1(new_n690_), .B2(new_n691_), .ZN(G1336gat));
  OAI21_X1  g491(.A(new_n434_), .B1(new_n684_), .B2(new_n387_), .ZN(new_n693_));
  OR2_X1    g492(.A1(new_n693_), .A2(KEYINPUT106), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(KEYINPUT106), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n387_), .A2(new_n434_), .ZN(new_n696_));
  AOI22_X1  g495(.A1(new_n694_), .A2(new_n695_), .B1(new_n690_), .B2(new_n696_), .ZN(G1337gat));
  NAND2_X1  g496(.A1(new_n604_), .A2(new_n423_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n684_), .A2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n688_), .A2(new_n604_), .A3(new_n689_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n700_), .B2(G99gat), .ZN(new_n701_));
  XOR2_X1   g500(.A(KEYINPUT107), .B(KEYINPUT51), .Z(new_n702_));
  XNOR2_X1  g501(.A(new_n701_), .B(new_n702_), .ZN(G1338gat));
  OAI211_X1 g502(.A(new_n290_), .B(new_n689_), .C1(new_n615_), .C2(new_n616_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT52), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n704_), .A2(new_n705_), .A3(G106gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n704_), .B2(G106gat), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n290_), .A2(new_n424_), .ZN(new_n708_));
  OAI22_X1  g507(.A1(new_n706_), .A2(new_n707_), .B1(new_n684_), .B2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g509(.A(KEYINPUT54), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n573_), .A2(new_n655_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT108), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n573_), .A2(new_n714_), .A3(new_n655_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n711_), .B1(new_n716_), .B2(new_n496_), .ZN(new_n717_));
  AOI211_X1 g516(.A(KEYINPUT108), .B(new_n654_), .C1(new_n567_), .C2(new_n572_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n714_), .B1(new_n573_), .B2(new_n655_), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n711_), .B(new_n496_), .C1(new_n718_), .C2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n717_), .A2(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n405_), .A2(new_n409_), .A3(new_n411_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n415_), .B1(new_n410_), .B2(new_n406_), .ZN(new_n724_));
  AOI22_X1  g523(.A1(new_n412_), .A2(new_n415_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n565_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n562_), .A2(KEYINPUT56), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT55), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n557_), .A2(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT71), .B1(new_n548_), .B2(KEYINPUT12), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n553_), .A2(new_n554_), .A3(new_n550_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n732_), .A2(KEYINPUT55), .A3(new_n551_), .A4(new_n552_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n729_), .A2(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n551_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n735_));
  OAI21_X1  g534(.A(KEYINPUT109), .B1(new_n735_), .B2(new_n544_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT109), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n542_), .A2(new_n543_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n732_), .A2(new_n737_), .A3(new_n738_), .A4(new_n551_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n736_), .A2(new_n540_), .A3(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n727_), .B1(new_n734_), .B2(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n564_), .B1(new_n734_), .B2(new_n740_), .ZN(new_n742_));
  OAI22_X1  g541(.A1(KEYINPUT111), .A2(new_n741_), .B1(new_n742_), .B2(KEYINPUT56), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n741_), .A2(KEYINPUT111), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n726_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT58), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  OAI211_X1 g546(.A(KEYINPUT58), .B(new_n726_), .C1(new_n743_), .C2(new_n744_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n747_), .A2(new_n614_), .A3(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT57), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n683_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n563_), .A2(new_n565_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(new_n725_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n418_), .A2(new_n565_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT56), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n729_), .A2(new_n733_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n732_), .A2(new_n738_), .A3(new_n551_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n539_), .B1(new_n757_), .B2(KEYINPUT109), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n756_), .B1(new_n739_), .B2(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n755_), .B1(new_n759_), .B2(new_n564_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n741_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n754_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n753_), .B1(new_n762_), .B2(KEYINPUT110), .ZN(new_n763_));
  INV_X1    g562(.A(new_n754_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n734_), .A2(new_n740_), .ZN(new_n765_));
  AOI21_X1  g564(.A(KEYINPUT56), .B1(new_n765_), .B2(new_n562_), .ZN(new_n766_));
  OAI211_X1 g565(.A(KEYINPUT110), .B(new_n764_), .C1(new_n766_), .C2(new_n741_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n751_), .B1(new_n763_), .B2(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n764_), .B1(new_n766_), .B2(new_n741_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT110), .ZN(new_n771_));
  AOI22_X1  g570(.A1(new_n770_), .A2(new_n771_), .B1(new_n752_), .B2(new_n725_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n683_), .B1(new_n772_), .B2(new_n767_), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n749_), .B(new_n769_), .C1(new_n773_), .C2(KEYINPUT57), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n722_), .B1(new_n774_), .B2(new_n536_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n604_), .B(new_n351_), .C1(new_n388_), .C2(new_n390_), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT112), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT112), .ZN(new_n778_));
  INV_X1    g577(.A(new_n776_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n496_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n736_), .A2(new_n540_), .A3(new_n739_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n562_), .B1(new_n781_), .B2(new_n756_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n741_), .B1(new_n782_), .B2(new_n755_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n771_), .B1(new_n783_), .B2(new_n754_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n784_), .A2(new_n767_), .A3(new_n753_), .ZN(new_n785_));
  AOI22_X1  g584(.A1(new_n780_), .A2(new_n748_), .B1(new_n785_), .B2(new_n751_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n494_), .B1(new_n763_), .B2(new_n768_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n750_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n537_), .B1(new_n786_), .B2(new_n788_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n778_), .B(new_n779_), .C1(new_n789_), .C2(new_n722_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n777_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(G113gat), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n792_), .A3(new_n418_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n749_), .A2(new_n769_), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT57), .B1(new_n785_), .B2(new_n494_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n536_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n722_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT59), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n798_), .B(new_n779_), .C1(KEYINPUT113), .C2(new_n799_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n799_), .A2(KEYINPUT113), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n799_), .A2(KEYINPUT113), .ZN(new_n802_));
  OAI22_X1  g601(.A1(new_n775_), .A2(new_n776_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n800_), .A2(new_n418_), .A3(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n793_), .B1(new_n792_), .B2(new_n804_), .ZN(G1340gat));
  NAND3_X1  g604(.A1(new_n800_), .A2(new_n574_), .A3(new_n803_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(G120gat), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n573_), .A2(KEYINPUT60), .ZN(new_n808_));
  MUX2_X1   g607(.A(new_n808_), .B(KEYINPUT60), .S(G120gat), .Z(new_n809_));
  NAND2_X1  g608(.A1(new_n791_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n807_), .A2(new_n810_), .ZN(G1341gat));
  AND4_X1   g610(.A1(G127gat), .A2(new_n800_), .A3(new_n537_), .A4(new_n803_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n777_), .A2(new_n537_), .A3(new_n790_), .ZN(new_n813_));
  INV_X1    g612(.A(G127gat), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n813_), .A2(KEYINPUT114), .A3(new_n814_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n812_), .B1(new_n817_), .B2(new_n818_), .ZN(G1342gat));
  AND4_X1   g618(.A1(G134gat), .A2(new_n800_), .A3(new_n614_), .A4(new_n803_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n777_), .A2(new_n683_), .A3(new_n790_), .ZN(new_n821_));
  INV_X1    g620(.A(G134gat), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n821_), .A2(KEYINPUT115), .A3(new_n822_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n820_), .B1(new_n825_), .B2(new_n826_), .ZN(G1343gat));
  NOR3_X1   g626(.A1(new_n775_), .A2(new_n604_), .A3(new_n289_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n591_), .A2(new_n577_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n418_), .A3(new_n829_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(KEYINPUT116), .B(G141gat), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n830_), .B(new_n831_), .ZN(G1344gat));
  NAND3_X1  g631(.A1(new_n828_), .A2(new_n574_), .A3(new_n829_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(KEYINPUT117), .B(G148gat), .ZN(new_n834_));
  XOR2_X1   g633(.A(new_n833_), .B(new_n834_), .Z(G1345gat));
  NAND3_X1  g634(.A1(new_n828_), .A2(new_n537_), .A3(new_n829_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(KEYINPUT61), .B(G155gat), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n836_), .B(new_n837_), .ZN(G1346gat));
  NOR2_X1   g637(.A1(new_n494_), .A2(G162gat), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n828_), .A2(new_n829_), .A3(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n604_), .A2(new_n289_), .ZN(new_n841_));
  AND4_X1   g640(.A1(new_n614_), .A2(new_n798_), .A3(new_n841_), .A4(new_n829_), .ZN(new_n842_));
  INV_X1    g641(.A(G162gat), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n840_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n840_), .B(KEYINPUT118), .C1(new_n843_), .C2(new_n842_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(G1347gat));
  XNOR2_X1  g647(.A(KEYINPUT120), .B(KEYINPUT62), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n387_), .A2(new_n351_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n604_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n852_), .A2(new_n420_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n798_), .A2(new_n850_), .A3(new_n289_), .A4(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(G169gat), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n290_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n850_), .B1(new_n856_), .B2(new_n853_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n849_), .B1(new_n855_), .B2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n798_), .A2(new_n289_), .A3(new_n853_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(KEYINPUT119), .ZN(new_n860_));
  INV_X1    g659(.A(new_n849_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n860_), .A2(new_n854_), .A3(G169gat), .A4(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n858_), .A2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n418_), .A2(new_n226_), .ZN(new_n864_));
  XOR2_X1   g663(.A(new_n864_), .B(KEYINPUT122), .Z(new_n865_));
  INV_X1    g664(.A(new_n852_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n289_), .B(new_n866_), .C1(new_n789_), .C2(new_n722_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(KEYINPUT121), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT121), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n798_), .A2(new_n870_), .A3(new_n289_), .A4(new_n866_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n865_), .B1(new_n869_), .B2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n863_), .A2(new_n873_), .ZN(G1348gat));
  OAI211_X1 g673(.A(new_n223_), .B(new_n574_), .C1(new_n869_), .C2(new_n872_), .ZN(new_n875_));
  OAI21_X1  g674(.A(G176gat), .B1(new_n867_), .B2(new_n573_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(G1349gat));
  OAI21_X1  g676(.A(new_n219_), .B1(new_n867_), .B2(new_n536_), .ZN(new_n878_));
  OR2_X1    g677(.A1(new_n536_), .A2(new_n207_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n879_), .B1(new_n868_), .B2(new_n871_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n878_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  AOI211_X1 g681(.A(KEYINPUT123), .B(new_n879_), .C1(new_n868_), .C2(new_n871_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1350gat));
  OAI211_X1 g683(.A(new_n208_), .B(new_n683_), .C1(new_n869_), .C2(new_n872_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n496_), .B1(new_n868_), .B2(new_n871_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n220_), .B2(new_n886_), .ZN(G1351gat));
  AND3_X1   g686(.A1(new_n798_), .A2(new_n841_), .A3(new_n851_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n888_), .A2(G197gat), .A3(new_n418_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT124), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n888_), .A2(new_n418_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n277_), .ZN(new_n893_));
  NAND4_X1  g692(.A1(new_n888_), .A2(KEYINPUT124), .A3(G197gat), .A4(new_n418_), .ZN(new_n894_));
  AND3_X1   g693(.A1(new_n891_), .A2(new_n893_), .A3(new_n894_), .ZN(G1352gat));
  NAND2_X1  g694(.A1(new_n888_), .A2(new_n574_), .ZN(new_n896_));
  INV_X1    g695(.A(G204gat), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(KEYINPUT125), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n897_), .A2(KEYINPUT125), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n896_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n900_), .B1(new_n896_), .B2(new_n898_), .ZN(G1353gat));
  AOI21_X1  g700(.A(new_n536_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n902_));
  XOR2_X1   g701(.A(new_n902_), .B(KEYINPUT126), .Z(new_n903_));
  NAND2_X1  g702(.A1(new_n888_), .A2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT127), .ZN(new_n905_));
  NOR2_X1   g704(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n904_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n906_), .B(KEYINPUT127), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n908_), .B1(new_n888_), .B2(new_n903_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n907_), .A2(new_n909_), .ZN(G1354gat));
  INV_X1    g709(.A(G218gat), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n888_), .A2(new_n911_), .A3(new_n683_), .ZN(new_n912_));
  AND2_X1   g711(.A1(new_n888_), .A2(new_n614_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n911_), .ZN(G1355gat));
endmodule


