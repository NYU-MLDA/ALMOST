//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1 1 1 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n740_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n841_, new_n842_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  OR3_X1    g003(.A1(new_n203_), .A2(new_n204_), .A3(KEYINPUT1), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT91), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT91), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n208_), .A2(G141gat), .A3(G148gat), .ZN(new_n209_));
  AND2_X1   g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n211_), .B1(new_n203_), .B2(KEYINPUT1), .ZN(new_n212_));
  AND3_X1   g011(.A1(new_n205_), .A2(new_n210_), .A3(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n203_), .A2(new_n204_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n207_), .A2(new_n209_), .A3(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT93), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT93), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n207_), .A2(new_n209_), .A3(new_n218_), .A4(new_n215_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n211_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT92), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n222_), .A2(KEYINPUT3), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(KEYINPUT3), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n221_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n222_), .A2(KEYINPUT3), .ZN(new_n226_));
  OAI22_X1  g025(.A1(new_n226_), .A2(new_n211_), .B1(new_n215_), .B2(new_n206_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n220_), .A2(KEYINPUT94), .A3(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(KEYINPUT94), .B1(new_n220_), .B2(new_n228_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n214_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT95), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n213_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  OAI211_X1 g032(.A(KEYINPUT95), .B(new_n214_), .C1(new_n229_), .C2(new_n230_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT29), .ZN(new_n236_));
  XOR2_X1   g035(.A(G197gat), .B(G204gat), .Z(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT21), .ZN(new_n238_));
  XOR2_X1   g037(.A(G211gat), .B(G218gat), .Z(new_n239_));
  AND2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G197gat), .B(G204gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT21), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n239_), .B1(new_n238_), .B2(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n240_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n236_), .A2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(G106gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n231_), .A2(new_n232_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT29), .ZN(new_n249_));
  INV_X1    g048(.A(new_n213_), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n248_), .A2(new_n249_), .A3(new_n234_), .A4(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(G22gat), .B(G50gat), .Z(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT96), .B(KEYINPUT28), .ZN(new_n254_));
  INV_X1    g053(.A(new_n252_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n233_), .A2(new_n249_), .A3(new_n234_), .A4(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n253_), .A2(new_n254_), .A3(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n254_), .B1(new_n253_), .B2(new_n256_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G228gat), .A2(G233gat), .ZN(new_n260_));
  INV_X1    g059(.A(G78gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  NOR3_X1   g061(.A1(new_n258_), .A2(new_n259_), .A3(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n262_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n253_), .A2(new_n256_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n254_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n264_), .B1(new_n267_), .B2(new_n257_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n247_), .B1(new_n263_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(G106gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n246_), .B(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n262_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n267_), .A2(new_n257_), .A3(new_n264_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n271_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G226gat), .A2(G233gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT19), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT20), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G183gat), .A2(G190gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT23), .ZN(new_n280_));
  OR2_X1    g079(.A1(G183gat), .A2(G190gat), .ZN(new_n281_));
  AOI22_X1  g080(.A1(new_n280_), .A2(new_n281_), .B1(G169gat), .B2(G176gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT22), .B(G169gat), .ZN(new_n283_));
  INV_X1    g082(.A(G176gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT25), .B(G183gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT26), .B(G190gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(G169gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(new_n284_), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n291_), .A2(KEYINPUT24), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n291_), .A2(KEYINPUT24), .A3(new_n293_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n289_), .A2(new_n280_), .A3(new_n292_), .A4(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n286_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n240_), .A2(new_n244_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n278_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n289_), .A2(new_n280_), .A3(new_n292_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT86), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n294_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT22), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n290_), .B1(new_n303_), .B2(KEYINPUT87), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT87), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n305_), .A2(KEYINPUT88), .A3(KEYINPUT22), .A4(G169gat), .ZN(new_n306_));
  OAI211_X1 g105(.A(new_n304_), .B(new_n306_), .C1(KEYINPUT88), .C2(KEYINPUT22), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n284_), .ZN(new_n308_));
  AOI22_X1  g107(.A1(new_n300_), .A2(new_n302_), .B1(new_n282_), .B2(new_n308_), .ZN(new_n309_));
  NOR3_X1   g108(.A1(new_n298_), .A2(new_n309_), .A3(KEYINPUT98), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT98), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n282_), .A2(new_n308_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n289_), .A2(new_n280_), .A3(new_n292_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n294_), .B(KEYINPUT86), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n312_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n311_), .B1(new_n315_), .B2(new_n245_), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n277_), .B(new_n299_), .C1(new_n310_), .C2(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(G64gat), .B(G92gat), .Z(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT100), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G8gat), .B(G36gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT20), .B1(new_n315_), .B2(new_n245_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT97), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n325_), .B1(new_n296_), .B2(new_n245_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n296_), .A2(new_n245_), .A3(new_n325_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n324_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n317_), .B(new_n323_), .C1(new_n329_), .C2(new_n277_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT104), .ZN(new_n331_));
  INV_X1    g130(.A(new_n328_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n332_), .A2(new_n326_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n276_), .B1(new_n333_), .B2(new_n324_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT104), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n334_), .A2(new_n335_), .A3(new_n323_), .A4(new_n317_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n278_), .B1(new_n298_), .B2(new_n309_), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n277_), .B(new_n337_), .C1(new_n332_), .C2(new_n326_), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT20), .B1(new_n296_), .B2(new_n245_), .ZN(new_n339_));
  OAI21_X1  g138(.A(KEYINPUT98), .B1(new_n298_), .B2(new_n309_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n315_), .A2(new_n311_), .A3(new_n245_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n339_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n338_), .B1(new_n342_), .B2(new_n277_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n323_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n331_), .A2(new_n336_), .A3(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT27), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n327_), .A2(new_n328_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n277_), .B1(new_n348_), .B2(new_n337_), .ZN(new_n349_));
  AOI211_X1 g148(.A(new_n276_), .B(new_n339_), .C1(new_n340_), .C2(new_n341_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n344_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT27), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(new_n352_), .A3(new_n330_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n347_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n269_), .A2(new_n274_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT105), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G15gat), .B(G43gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT89), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT30), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT31), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G227gat), .A2(G233gat), .ZN(new_n362_));
  INV_X1    g161(.A(G71gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(G99gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n309_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n361_), .B(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n367_), .B(KEYINPUT90), .Z(new_n368_));
  XNOR2_X1  g167(.A(G127gat), .B(G134gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G113gat), .B(G120gat), .ZN(new_n370_));
  XOR2_X1   g169(.A(new_n369_), .B(new_n370_), .Z(new_n371_));
  XNOR2_X1  g170(.A(new_n368_), .B(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n235_), .A2(new_n371_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n371_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n233_), .A2(new_n374_), .A3(new_n234_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n373_), .A2(KEYINPUT4), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT4), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n235_), .A2(new_n377_), .A3(new_n371_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G225gat), .A2(G233gat), .ZN(new_n379_));
  XOR2_X1   g178(.A(new_n379_), .B(KEYINPUT101), .Z(new_n380_));
  NAND3_X1  g179(.A1(new_n376_), .A2(new_n378_), .A3(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G1gat), .B(G29gat), .ZN(new_n382_));
  INV_X1    g181(.A(G85gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT0), .B(G57gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n373_), .A2(new_n375_), .A3(new_n379_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n381_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n386_), .B1(new_n381_), .B2(new_n387_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n269_), .A2(new_n354_), .A3(new_n274_), .A4(KEYINPUT105), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n357_), .A2(new_n372_), .A3(new_n391_), .A4(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT102), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n394_), .A2(KEYINPUT33), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n388_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n351_), .A2(new_n330_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n373_), .A2(new_n375_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n386_), .B1(new_n398_), .B2(new_n380_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n376_), .A2(new_n379_), .A3(new_n378_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n397_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n395_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n381_), .A2(new_n386_), .A3(new_n387_), .A4(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n396_), .A2(new_n401_), .A3(new_n403_), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n323_), .A2(KEYINPUT32), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT103), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n405_), .A2(new_n343_), .A3(new_n406_), .ZN(new_n407_));
  NOR3_X1   g206(.A1(new_n405_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n406_), .B1(new_n405_), .B2(new_n343_), .ZN(new_n409_));
  NOR3_X1   g208(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n410_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n404_), .A2(new_n411_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n269_), .A2(new_n274_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n351_), .A2(new_n352_), .A3(new_n330_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n414_), .B1(KEYINPUT27), .B2(new_n346_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n415_), .B1(new_n269_), .B2(new_n274_), .ZN(new_n416_));
  AOI22_X1  g215(.A1(new_n412_), .A2(new_n413_), .B1(new_n416_), .B2(new_n391_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n393_), .B1(new_n417_), .B2(new_n372_), .ZN(new_n418_));
  INV_X1    g217(.A(G36gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(G29gat), .ZN(new_n420_));
  INV_X1    g219(.A(G29gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(G36gat), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n420_), .A2(new_n422_), .A3(KEYINPUT75), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT75), .B1(new_n420_), .B2(new_n422_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT76), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT75), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n421_), .A2(G36gat), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n419_), .A2(G29gat), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n426_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT76), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n420_), .A2(new_n422_), .A3(KEYINPUT75), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n429_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n425_), .A2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G43gat), .B(G50gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n425_), .A2(new_n432_), .A3(new_n434_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G15gat), .B(G22gat), .ZN(new_n439_));
  INV_X1    g238(.A(G1gat), .ZN(new_n440_));
  INV_X1    g239(.A(G8gat), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT14), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n439_), .A2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G1gat), .B(G8gat), .ZN(new_n444_));
  XOR2_X1   g243(.A(new_n443_), .B(new_n444_), .Z(new_n445_));
  XNOR2_X1  g244(.A(new_n438_), .B(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n446_), .A2(G229gat), .A3(G233gat), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT15), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n425_), .A2(new_n434_), .A3(new_n432_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n434_), .B1(new_n425_), .B2(new_n432_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n448_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n436_), .A2(KEYINPUT15), .A3(new_n437_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n445_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n451_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G229gat), .A2(G233gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n438_), .A2(new_n445_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n454_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n447_), .B1(new_n457_), .B2(KEYINPUT85), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n458_), .B1(KEYINPUT85), .B2(new_n457_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G113gat), .B(G141gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G169gat), .B(G197gat), .ZN(new_n461_));
  XOR2_X1   g260(.A(new_n460_), .B(new_n461_), .Z(new_n462_));
  XNOR2_X1  g261(.A(new_n459_), .B(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT8), .ZN(new_n464_));
  NOR2_X1   g263(.A1(G85gat), .A2(G92gat), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT69), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G85gat), .A2(G92gat), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  AND2_X1   g268(.A1(G85gat), .A2(G92gat), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT69), .B1(new_n470_), .B2(new_n465_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n473_));
  NOR2_X1   g272(.A1(G99gat), .A2(G106gat), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT7), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT6), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n477_), .B1(G99gat), .B2(G106gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G99gat), .A2(G106gat), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n479_), .A2(KEYINPUT6), .ZN(new_n480_));
  OAI211_X1 g279(.A(new_n473_), .B(new_n476_), .C1(new_n478_), .C2(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n464_), .B1(new_n472_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT68), .B(KEYINPUT8), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n469_), .A2(new_n471_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n476_), .A2(new_n473_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT65), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n488_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n479_), .A2(KEYINPUT6), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n477_), .A2(G99gat), .A3(G106gat), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(KEYINPUT65), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n487_), .B1(new_n489_), .B2(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n486_), .B1(new_n493_), .B2(KEYINPUT67), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n476_), .A2(new_n473_), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n490_), .A2(new_n491_), .A3(KEYINPUT65), .ZN(new_n496_));
  AOI21_X1  g295(.A(KEYINPUT65), .B1(new_n490_), .B2(new_n491_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n495_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT67), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n483_), .B1(new_n494_), .B2(new_n500_), .ZN(new_n501_));
  OR2_X1    g300(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(new_n270_), .A3(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n504_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n465_), .B1(new_n470_), .B2(KEYINPUT9), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT64), .B1(new_n470_), .B2(KEYINPUT9), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT64), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT9), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n468_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n506_), .A2(new_n507_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT66), .ZN(new_n512_));
  NOR3_X1   g311(.A1(new_n505_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n502_), .A2(new_n270_), .A3(new_n503_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n514_), .B1(new_n489_), .B2(new_n492_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n506_), .A2(new_n507_), .A3(new_n510_), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT66), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n513_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n501_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G57gat), .B(G64gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT11), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT71), .ZN(new_n522_));
  XOR2_X1   g321(.A(G71gat), .B(G78gat), .Z(new_n523_));
  OAI21_X1  g322(.A(new_n523_), .B1(KEYINPUT11), .B2(new_n520_), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n522_), .A2(new_n524_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n519_), .A2(KEYINPUT12), .A3(new_n525_), .A4(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n526_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT70), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n485_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n493_), .A2(KEYINPUT67), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n482_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n512_), .B1(new_n505_), .B2(new_n511_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n515_), .A2(KEYINPUT66), .A3(new_n516_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n529_), .B1(new_n532_), .B2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n501_), .A2(new_n518_), .A3(KEYINPUT70), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n528_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT74), .B(KEYINPUT12), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n527_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n536_), .A2(new_n537_), .A3(new_n528_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G230gat), .A2(G233gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT72), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n541_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n541_), .A2(new_n545_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n538_), .B1(new_n548_), .B2(KEYINPUT73), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT73), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n546_), .A2(new_n550_), .A3(new_n547_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n542_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n544_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G120gat), .B(G148gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT5), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G176gat), .B(G204gat), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n556_), .B(new_n557_), .Z(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n554_), .A2(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n542_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n558_), .B1(new_n561_), .B2(new_n544_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n560_), .A2(KEYINPUT13), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(KEYINPUT13), .B1(new_n560_), .B2(new_n562_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n418_), .A2(new_n463_), .A3(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n536_), .A2(new_n537_), .A3(new_n438_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT79), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n536_), .A2(new_n537_), .A3(KEYINPUT79), .A4(new_n438_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G232gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT34), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT35), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n570_), .A2(new_n571_), .A3(new_n576_), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n451_), .B(new_n452_), .C1(new_n532_), .C2(new_n535_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT77), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT77), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n519_), .A2(new_n580_), .A3(new_n452_), .A4(new_n451_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n582_), .B1(new_n575_), .B2(new_n574_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n577_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT80), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n568_), .A2(new_n569_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n571_), .A2(new_n576_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n585_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n579_), .A2(new_n581_), .A3(KEYINPUT78), .ZN(new_n589_));
  AOI21_X1  g388(.A(KEYINPUT78), .B1(new_n579_), .B2(new_n581_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n570_), .A2(KEYINPUT80), .A3(new_n571_), .A4(new_n576_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n588_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n574_), .A2(new_n575_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n584_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G190gat), .B(G218gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G134gat), .B(G162gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT36), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n595_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT82), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n593_), .A2(new_n594_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n584_), .ZN(new_n603_));
  XOR2_X1   g402(.A(KEYINPUT81), .B(KEYINPUT36), .Z(new_n604_));
  NOR2_X1   g403(.A1(new_n598_), .A2(new_n604_), .ZN(new_n605_));
  AND4_X1   g404(.A1(new_n601_), .A2(new_n602_), .A3(new_n603_), .A4(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n601_), .B1(new_n595_), .B2(new_n605_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n600_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT83), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT37), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n608_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n602_), .A2(new_n603_), .A3(new_n605_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT82), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n595_), .A2(new_n601_), .A3(new_n605_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(KEYINPUT83), .A2(KEYINPUT37), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n609_), .A2(new_n610_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n615_), .A2(new_n600_), .A3(new_n616_), .A4(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n611_), .A2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G127gat), .B(G155gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT16), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G183gat), .B(G211gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(G231gat), .A2(G233gat), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n445_), .B(new_n624_), .Z(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(new_n528_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n623_), .B1(new_n626_), .B2(KEYINPUT84), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT17), .B1(new_n626_), .B2(new_n623_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  OAI211_X1 g428(.A(KEYINPUT17), .B(new_n623_), .C1(new_n626_), .C2(KEYINPUT84), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n619_), .A2(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n567_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n391_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n634_), .A2(new_n440_), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT38), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n637_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n608_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n640_), .A2(new_n632_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n567_), .A2(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G1gat), .B1(new_n642_), .B2(new_n391_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n638_), .A2(new_n639_), .A3(new_n643_), .ZN(G1324gat));
  NAND3_X1  g443(.A1(new_n634_), .A2(new_n441_), .A3(new_n415_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n646_));
  INV_X1    g445(.A(new_n642_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(new_n415_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n646_), .B1(new_n648_), .B2(G8gat), .ZN(new_n649_));
  AOI211_X1 g448(.A(KEYINPUT39), .B(new_n441_), .C1(new_n647_), .C2(new_n415_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n645_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g451(.A(new_n372_), .ZN(new_n653_));
  OAI21_X1  g452(.A(G15gat), .B1(new_n642_), .B2(new_n653_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT41), .Z(new_n655_));
  INV_X1    g454(.A(G15gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n634_), .A2(new_n656_), .A3(new_n372_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(G1326gat));
  XOR2_X1   g457(.A(new_n413_), .B(KEYINPUT106), .Z(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(G22gat), .B1(new_n642_), .B2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT42), .ZN(new_n662_));
  INV_X1    g461(.A(G22gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n634_), .A2(new_n663_), .A3(new_n659_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(G1327gat));
  OR2_X1    g464(.A1(new_n564_), .A2(new_n565_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n463_), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n666_), .A2(new_n667_), .A3(new_n631_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT43), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n619_), .A2(new_n418_), .A3(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n669_), .B1(new_n619_), .B2(new_n418_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n668_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  OAI211_X1 g473(.A(new_n668_), .B(KEYINPUT44), .C1(new_n670_), .C2(new_n671_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n391_), .A2(new_n421_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n608_), .A2(new_n631_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n567_), .A2(new_n635_), .A3(new_n678_), .ZN(new_n679_));
  AOI22_X1  g478(.A1(new_n676_), .A2(new_n677_), .B1(new_n421_), .B2(new_n679_), .ZN(G1328gat));
  XNOR2_X1  g479(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n674_), .A2(new_n415_), .A3(new_n675_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(G36gat), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT107), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n682_), .A2(KEYINPUT107), .A3(G36gat), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n567_), .A2(new_n419_), .A3(new_n415_), .A4(new_n678_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT45), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n681_), .B1(new_n687_), .B2(new_n689_), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n682_), .A2(KEYINPUT107), .A3(G36gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(KEYINPUT107), .B1(new_n682_), .B2(G36gat), .ZN(new_n692_));
  OAI211_X1 g491(.A(new_n689_), .B(new_n681_), .C1(new_n691_), .C2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n690_), .A2(new_n694_), .ZN(G1329gat));
  NAND3_X1  g494(.A1(new_n676_), .A2(G43gat), .A3(new_n372_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n567_), .A2(new_n678_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n697_), .A2(new_n653_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n696_), .B1(G43gat), .B2(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g499(.A(new_n413_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n676_), .A2(G50gat), .A3(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(G50gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n703_), .B1(new_n697_), .B2(new_n660_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n702_), .A2(new_n704_), .ZN(G1331gat));
  AND3_X1   g504(.A1(new_n418_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n706_), .A2(new_n633_), .ZN(new_n707_));
  INV_X1    g506(.A(G57gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n707_), .A2(new_n708_), .A3(new_n635_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n706_), .A2(new_n641_), .ZN(new_n710_));
  OAI21_X1  g509(.A(G57gat), .B1(new_n710_), .B2(new_n391_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n711_), .ZN(G1332gat));
  INV_X1    g511(.A(G64gat), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n707_), .A2(new_n713_), .A3(new_n415_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n710_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(new_n415_), .ZN(new_n716_));
  XOR2_X1   g515(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n717_));
  AND3_X1   g516(.A1(new_n716_), .A2(G64gat), .A3(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n716_), .B2(G64gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n714_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT110), .Z(G1333gat));
  NAND3_X1  g520(.A1(new_n707_), .A2(new_n363_), .A3(new_n372_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n715_), .A2(new_n372_), .ZN(new_n723_));
  XOR2_X1   g522(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n724_));
  AND3_X1   g523(.A1(new_n723_), .A2(G71gat), .A3(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n723_), .B2(G71gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n722_), .B1(new_n725_), .B2(new_n726_), .ZN(G1334gat));
  OAI21_X1  g526(.A(G78gat), .B1(new_n710_), .B2(new_n660_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT50), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n707_), .A2(new_n261_), .A3(new_n659_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1335gat));
  AND2_X1   g530(.A1(new_n706_), .A2(new_n678_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n732_), .A2(new_n383_), .A3(new_n635_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n566_), .A2(new_n463_), .A3(new_n631_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n734_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n735_));
  OAI21_X1  g534(.A(G85gat), .B1(new_n735_), .B2(new_n391_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n733_), .A2(new_n736_), .ZN(G1336gat));
  INV_X1    g536(.A(G92gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n732_), .A2(new_n738_), .A3(new_n415_), .ZN(new_n739_));
  OAI21_X1  g538(.A(G92gat), .B1(new_n735_), .B2(new_n354_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1337gat));
  NAND4_X1  g540(.A1(new_n732_), .A2(new_n502_), .A3(new_n503_), .A4(new_n372_), .ZN(new_n742_));
  OAI21_X1  g541(.A(G99gat), .B1(new_n735_), .B2(new_n653_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT51), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n745_), .A2(KEYINPUT112), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n744_), .B(new_n746_), .ZN(G1338gat));
  OAI211_X1 g546(.A(new_n701_), .B(new_n734_), .C1(new_n670_), .C2(new_n671_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT113), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(G106gat), .B1(new_n748_), .B2(KEYINPUT113), .ZN(new_n751_));
  OAI21_X1  g550(.A(KEYINPUT52), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n748_), .A2(KEYINPUT113), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n753_), .A2(new_n754_), .A3(G106gat), .A4(new_n749_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n752_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n732_), .A2(new_n270_), .A3(new_n701_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n756_), .A2(new_n757_), .A3(new_n759_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(G1339gat));
  NAND2_X1  g562(.A1(new_n454_), .A2(new_n456_), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n764_), .A2(new_n455_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n462_), .B1(new_n446_), .B2(new_n455_), .ZN(new_n766_));
  AOI22_X1  g565(.A1(new_n459_), .A2(new_n462_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n562_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n561_), .A2(new_n544_), .A3(new_n558_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n767_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n553_), .B1(new_n548_), .B2(new_n540_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n544_), .A2(KEYINPUT55), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n773_), .B1(new_n540_), .B2(new_n543_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n771_), .A2(new_n772_), .A3(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n558_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT115), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n777_), .B2(KEYINPUT56), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT56), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n775_), .A2(KEYINPUT115), .A3(new_n779_), .A4(new_n558_), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n778_), .A2(new_n560_), .A3(new_n463_), .A4(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n770_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT57), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n782_), .A2(new_n608_), .A3(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n786_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n776_), .A2(KEYINPUT56), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n775_), .A2(new_n779_), .A3(new_n558_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n560_), .A2(new_n788_), .A3(new_n767_), .A4(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT58), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n791_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n619_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n782_), .A2(KEYINPUT116), .A3(KEYINPUT57), .A4(new_n608_), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n787_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n611_), .A2(new_n618_), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n564_), .A2(new_n565_), .A3(new_n463_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(new_n631_), .A3(new_n798_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n799_), .A2(KEYINPUT54), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(KEYINPUT54), .ZN(new_n801_));
  OAI22_X1  g600(.A1(new_n796_), .A2(new_n631_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n357_), .A2(new_n372_), .A3(new_n392_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n802_), .A2(new_n635_), .A3(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n806_), .A2(KEYINPUT59), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n806_), .A2(KEYINPUT59), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n805_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n806_), .A2(KEYINPUT59), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n802_), .A2(new_n635_), .A3(new_n804_), .A4(new_n810_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n463_), .A2(G113gat), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT119), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n805_), .A2(KEYINPUT117), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT117), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n802_), .A2(new_n816_), .A3(new_n635_), .A4(new_n804_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n815_), .A2(new_n463_), .A3(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(G113gat), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n812_), .A2(new_n814_), .B1(new_n818_), .B2(new_n819_), .ZN(G1340gat));
  NAND3_X1  g619(.A1(new_n809_), .A2(new_n666_), .A3(new_n811_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(G120gat), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n566_), .A2(KEYINPUT60), .ZN(new_n823_));
  MUX2_X1   g622(.A(new_n823_), .B(KEYINPUT60), .S(G120gat), .Z(new_n824_));
  NAND3_X1  g623(.A1(new_n815_), .A2(new_n817_), .A3(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n822_), .A2(new_n825_), .ZN(G1341gat));
  NAND3_X1  g625(.A1(new_n809_), .A2(new_n631_), .A3(new_n811_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(G127gat), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n632_), .A2(G127gat), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n815_), .A2(new_n817_), .A3(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(G1342gat));
  NAND2_X1  g630(.A1(new_n619_), .A2(G134gat), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(KEYINPUT120), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n815_), .A2(new_n640_), .A3(new_n817_), .ZN(new_n834_));
  INV_X1    g633(.A(G134gat), .ZN(new_n835_));
  AOI22_X1  g634(.A1(new_n812_), .A2(new_n833_), .B1(new_n834_), .B2(new_n835_), .ZN(G1343gat));
  NOR3_X1   g635(.A1(new_n413_), .A2(new_n372_), .A3(new_n415_), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n802_), .A2(new_n635_), .A3(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n463_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n666_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(KEYINPUT121), .B(G148gat), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n841_), .B(new_n842_), .ZN(G1345gat));
  NAND2_X1  g642(.A1(new_n838_), .A2(new_n631_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(KEYINPUT61), .B(G155gat), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n844_), .B(new_n845_), .ZN(G1346gat));
  NAND4_X1  g645(.A1(new_n802_), .A2(new_n635_), .A3(new_n640_), .A4(new_n837_), .ZN(new_n847_));
  INV_X1    g646(.A(G162gat), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  OR2_X1    g648(.A1(new_n849_), .A2(KEYINPUT122), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(KEYINPUT122), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n797_), .A2(new_n848_), .ZN(new_n852_));
  AOI22_X1  g651(.A1(new_n850_), .A2(new_n851_), .B1(new_n838_), .B2(new_n852_), .ZN(G1347gat));
  AND2_X1   g652(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n372_), .A2(new_n391_), .A3(new_n415_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n855_), .A2(new_n667_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n659_), .B1(KEYINPUT123), .B2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(KEYINPUT123), .B2(new_n856_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  AOI211_X1 g658(.A(new_n290_), .B(new_n854_), .C1(new_n802_), .C2(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n860_), .B(new_n861_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n799_), .B(KEYINPUT54), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n787_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n632_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n354_), .B1(new_n863_), .B2(new_n865_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n659_), .A2(new_n653_), .A3(new_n635_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n869_), .A2(new_n463_), .A3(new_n283_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n862_), .A2(new_n870_), .ZN(G1348gat));
  OAI21_X1  g670(.A(new_n284_), .B1(new_n868_), .B2(new_n566_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT125), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  OAI211_X1 g673(.A(KEYINPUT125), .B(new_n284_), .C1(new_n868_), .C2(new_n566_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n701_), .B1(new_n863_), .B2(new_n865_), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n566_), .A2(new_n284_), .A3(new_n855_), .ZN(new_n877_));
  AOI22_X1  g676(.A1(new_n874_), .A2(new_n875_), .B1(new_n876_), .B2(new_n877_), .ZN(G1349gat));
  NOR2_X1   g677(.A1(new_n632_), .A2(new_n287_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n866_), .A2(new_n867_), .A3(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT126), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n855_), .A2(new_n632_), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n802_), .A2(new_n881_), .A3(new_n413_), .A4(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(G183gat), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n881_), .B1(new_n876_), .B2(new_n882_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n880_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(KEYINPUT127), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT127), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n889_), .B(new_n880_), .C1(new_n885_), .C2(new_n886_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n890_), .ZN(G1350gat));
  OAI21_X1  g690(.A(G190gat), .B1(new_n868_), .B2(new_n797_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n640_), .A2(new_n288_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n868_), .B2(new_n893_), .ZN(G1351gat));
  NOR3_X1   g693(.A1(new_n413_), .A2(new_n372_), .A3(new_n635_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n866_), .A2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n463_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n666_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G204gat), .ZN(G1353gat));
  XNOR2_X1  g700(.A(KEYINPUT63), .B(G211gat), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n897_), .A2(new_n631_), .A3(new_n902_), .ZN(new_n903_));
  OAI22_X1  g702(.A1(new_n896_), .A2(new_n632_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1354gat));
  OAI21_X1  g704(.A(G218gat), .B1(new_n896_), .B2(new_n797_), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n608_), .A2(G218gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n896_), .B2(new_n907_), .ZN(G1355gat));
endmodule


