//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 1 1 1 1 1 1 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 1 1 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n799_, new_n800_, new_n801_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n819_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n842_, new_n844_, new_n845_,
    new_n847_, new_n848_, new_n849_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_;
  NAND2_X1  g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT81), .Z(new_n203_));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n204_), .B1(new_n205_), .B2(KEYINPUT1), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n206_), .B1(KEYINPUT1), .B2(new_n204_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n203_), .A2(new_n207_), .A3(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT82), .ZN(new_n211_));
  OR2_X1    g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n203_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT85), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT84), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n218_), .B1(new_n208_), .B2(KEYINPUT83), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT3), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT83), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n221_), .B1(new_n220_), .B2(KEYINPUT84), .ZN(new_n222_));
  AOI22_X1  g021(.A1(new_n219_), .A2(new_n220_), .B1(new_n208_), .B2(new_n222_), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n204_), .B(new_n212_), .C1(new_n217_), .C2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n211_), .A2(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(G127gat), .B(G134gat), .Z(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT80), .ZN(new_n227_));
  XOR2_X1   g026(.A(G113gat), .B(G120gat), .Z(new_n228_));
  XOR2_X1   g027(.A(new_n227_), .B(new_n228_), .Z(new_n229_));
  NAND2_X1  g028(.A1(new_n225_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n227_), .B(new_n228_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n231_), .A2(new_n211_), .A3(new_n224_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G225gat), .A2(G233gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n230_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT97), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n230_), .A2(KEYINPUT97), .A3(new_n232_), .A4(new_n233_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n230_), .A2(KEYINPUT4), .A3(new_n232_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n233_), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n239_), .B(new_n240_), .C1(KEYINPUT4), .C2(new_n230_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G1gat), .B(G29gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT0), .ZN(new_n244_));
  INV_X1    g043(.A(G57gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(G85gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n242_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n248_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n238_), .A2(new_n241_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G211gat), .B(G218gat), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n253_), .A2(KEYINPUT88), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(KEYINPUT88), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(G197gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(G204gat), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n257_), .A2(G204gat), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT21), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n260_), .B1(KEYINPUT87), .B2(new_n258_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n262_), .B1(KEYINPUT87), .B2(new_n258_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n256_), .B(new_n261_), .C1(new_n263_), .C2(KEYINPUT21), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n254_), .A2(KEYINPUT89), .A3(new_n255_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(KEYINPUT21), .A3(new_n263_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT89), .B1(new_n254_), .B2(new_n255_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n264_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n225_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT29), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n268_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G228gat), .A2(G233gat), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n272_), .B1(new_n268_), .B2(KEYINPUT90), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  OAI221_X1 g073(.A(new_n268_), .B1(KEYINPUT90), .B2(new_n272_), .C1(new_n269_), .C2(new_n270_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G78gat), .B(G106gat), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n274_), .A2(new_n275_), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT91), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n277_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT28), .B1(new_n225_), .B2(KEYINPUT29), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NOR3_X1   g082(.A1(new_n225_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n284_));
  XOR2_X1   g083(.A(G22gat), .B(G50gat), .Z(new_n285_));
  NOR3_X1   g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n285_), .ZN(new_n287_));
  OR3_X1    g086(.A1(new_n225_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n287_), .B1(new_n288_), .B2(new_n282_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n286_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT91), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n274_), .A2(new_n275_), .A3(new_n291_), .A4(new_n277_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n279_), .A2(new_n281_), .A3(new_n290_), .A4(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT86), .B1(new_n286_), .B2(new_n289_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n285_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT86), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n288_), .A2(new_n282_), .A3(new_n287_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n295_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  AND3_X1   g097(.A1(new_n274_), .A2(new_n275_), .A3(new_n277_), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n294_), .B(new_n298_), .C1(new_n299_), .C2(new_n280_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n293_), .A2(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(G71gat), .B(G99gat), .Z(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(G43gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G227gat), .A2(G233gat), .ZN(new_n304_));
  INV_X1    g103(.A(G15gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n303_), .B(new_n306_), .Z(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  OR2_X1    g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G169gat), .A2(G176gat), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(KEYINPUT24), .A3(new_n310_), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n309_), .A2(KEYINPUT24), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G183gat), .A2(G190gat), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT23), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(G190gat), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n318_), .A2(KEYINPUT26), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(KEYINPUT26), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n319_), .B1(KEYINPUT78), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT25), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n322_), .A2(G183gat), .ZN(new_n323_));
  OAI221_X1 g122(.A(new_n321_), .B1(KEYINPUT76), .B2(new_n323_), .C1(KEYINPUT78), .C2(new_n320_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(KEYINPUT76), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n322_), .A2(G183gat), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT77), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n322_), .A2(KEYINPUT77), .A3(G183gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n325_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  OAI211_X1 g129(.A(new_n311_), .B(new_n317_), .C1(new_n324_), .C2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n310_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT22), .B(G169gat), .ZN(new_n333_));
  INV_X1    g132(.A(G176gat), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n332_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n314_), .A2(KEYINPUT23), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n315_), .A2(G183gat), .A3(G190gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(KEYINPUT79), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT79), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n339_), .A2(new_n315_), .A3(G183gat), .A4(G190gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(G183gat), .A2(G190gat), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n335_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n331_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT30), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n344_), .A2(new_n345_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n308_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n348_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n350_), .A2(new_n307_), .A3(new_n346_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT31), .ZN(new_n352_));
  AND3_X1   g151(.A1(new_n349_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n352_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n229_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n349_), .A2(new_n351_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT31), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n349_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n357_), .A2(new_n231_), .A3(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n355_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n301_), .A2(new_n360_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n355_), .A2(new_n359_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n362_), .A2(new_n300_), .A3(new_n293_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n252_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n335_), .B1(new_n316_), .B2(new_n342_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n312_), .A2(new_n338_), .A3(new_n340_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT26), .B(G190gat), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT94), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n323_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n326_), .ZN(new_n371_));
  OAI221_X1 g170(.A(new_n311_), .B1(new_n366_), .B2(KEYINPUT95), .C1(new_n369_), .C2(new_n371_), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n366_), .A2(KEYINPUT95), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n365_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  OR2_X1    g173(.A1(new_n374_), .A2(new_n268_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G226gat), .A2(G233gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n344_), .A2(new_n268_), .ZN(new_n379_));
  AND4_X1   g178(.A1(KEYINPUT20), .A2(new_n375_), .A3(new_n378_), .A4(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT20), .B1(new_n344_), .B2(new_n268_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT93), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n374_), .A2(new_n268_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT96), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n378_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n380_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G8gat), .B(G36gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT18), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G64gat), .B(G92gat), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n390_), .B(new_n391_), .Z(new_n392_));
  NAND2_X1  g191(.A1(new_n388_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n392_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n378_), .B1(new_n383_), .B2(new_n385_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n394_), .B1(new_n395_), .B2(new_n380_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n393_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT27), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n398_), .B1(new_n388_), .B2(new_n392_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n386_), .A2(new_n378_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n375_), .A2(KEYINPUT20), .A3(new_n387_), .A4(new_n379_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n400_), .A2(new_n394_), .A3(new_n401_), .ZN(new_n402_));
  AOI22_X1  g201(.A1(new_n397_), .A2(new_n398_), .B1(new_n399_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT32), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n388_), .B1(new_n404_), .B2(new_n394_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n400_), .A2(KEYINPUT32), .A3(new_n392_), .A4(new_n401_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(new_n252_), .A3(new_n406_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n238_), .A2(KEYINPUT33), .A3(new_n241_), .A4(new_n250_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n230_), .A2(new_n232_), .A3(new_n240_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n409_), .A2(new_n248_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n231_), .B1(new_n211_), .B2(new_n224_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT4), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n240_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n239_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT99), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT99), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n410_), .A2(new_n414_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n393_), .A2(new_n396_), .A3(new_n408_), .A4(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT98), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT33), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n251_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n421_), .B1(new_n251_), .B2(new_n422_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n407_), .B1(new_n420_), .B2(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n301_), .A2(new_n362_), .ZN(new_n427_));
  AOI22_X1  g226(.A1(new_n364_), .A2(new_n403_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G229gat), .A2(G233gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G15gat), .B(G22gat), .ZN(new_n430_));
  INV_X1    g229(.A(G1gat), .ZN(new_n431_));
  INV_X1    g230(.A(G8gat), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT14), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n430_), .A2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G1gat), .B(G8gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(G43gat), .B(G50gat), .Z(new_n437_));
  XNOR2_X1  g236(.A(G29gat), .B(G36gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  OR2_X1    g238(.A1(new_n436_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n436_), .A2(new_n439_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n429_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n442_), .A2(KEYINPUT75), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(KEYINPUT75), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT15), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n439_), .B(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n436_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(new_n429_), .A3(new_n440_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n443_), .A2(new_n444_), .A3(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G113gat), .B(G141gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G169gat), .B(G197gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n449_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n452_), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n443_), .A2(new_n444_), .A3(new_n448_), .A4(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT12), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NOR3_X1   g259(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT67), .ZN(new_n463_));
  AND3_X1   g262(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n464_));
  AOI21_X1  g263(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n463_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G99gat), .A2(G106gat), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT6), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n469_), .A2(KEYINPUT67), .A3(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n462_), .A2(new_n466_), .A3(new_n471_), .ZN(new_n472_));
  AND2_X1   g271(.A1(G85gat), .A2(G92gat), .ZN(new_n473_));
  NOR2_X1   g272(.A1(G85gat), .A2(G92gat), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n472_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT8), .ZN(new_n477_));
  INV_X1    g276(.A(new_n461_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n478_), .A2(new_n469_), .A3(new_n470_), .A4(new_n459_), .ZN(new_n479_));
  XOR2_X1   g278(.A(KEYINPUT66), .B(KEYINPUT8), .Z(new_n480_));
  NAND3_X1  g279(.A1(new_n479_), .A2(new_n475_), .A3(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT9), .B1(new_n473_), .B2(new_n474_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT64), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G85gat), .A2(G92gat), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT9), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n483_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n482_), .A2(new_n486_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n483_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n488_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n489_));
  OR2_X1    g288(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n490_));
  INV_X1    g289(.A(G106gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n487_), .A2(new_n489_), .A3(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT65), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n464_), .A2(new_n465_), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n497_), .A2(new_n493_), .A3(new_n488_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(KEYINPUT65), .A3(new_n487_), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n477_), .A2(new_n481_), .B1(new_n496_), .B2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT68), .B(G71gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(G78gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G57gat), .B(G64gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT11), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(G78gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n501_), .B(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n503_), .A2(KEYINPUT11), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n505_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n458_), .B1(new_n500_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G230gat), .A2(G233gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n500_), .A2(new_n511_), .ZN(new_n514_));
  AOI21_X1  g313(.A(KEYINPUT65), .B1(new_n498_), .B2(new_n487_), .ZN(new_n515_));
  AND4_X1   g314(.A1(KEYINPUT65), .A2(new_n487_), .A3(new_n489_), .A4(new_n493_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT8), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n517_), .B1(new_n472_), .B2(new_n475_), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n479_), .A2(new_n475_), .A3(new_n480_), .ZN(new_n519_));
  OAI22_X1  g318(.A1(new_n515_), .A2(new_n516_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n520_), .A2(KEYINPUT12), .A3(new_n510_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n512_), .A2(new_n513_), .A3(new_n514_), .A4(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n520_), .B(new_n511_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n522_), .B1(new_n513_), .B2(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(G120gat), .B(G148gat), .Z(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT5), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G176gat), .B(G204gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n524_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT13), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT69), .ZN(new_n531_));
  NOR3_X1   g330(.A1(new_n428_), .A2(new_n457_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n446_), .A2(new_n520_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G232gat), .A2(G233gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT71), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT35), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n533_), .B(new_n539_), .C1(new_n520_), .C2(new_n439_), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n537_), .A2(new_n538_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G190gat), .B(G218gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G134gat), .B(G162gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n546_), .B(KEYINPUT36), .Z(new_n547_));
  NAND2_X1  g346(.A1(new_n543_), .A2(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n546_), .A2(KEYINPUT36), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n542_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT37), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G231gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n436_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(new_n511_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT73), .B(KEYINPUT17), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G127gat), .B(G155gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT16), .ZN(new_n560_));
  XOR2_X1   g359(.A(G183gat), .B(G211gat), .Z(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n558_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n558_), .A2(new_n562_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(KEYINPUT72), .B(KEYINPUT17), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n556_), .A2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n563_), .A2(new_n564_), .A3(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT74), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n553_), .A2(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n532_), .A2(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n252_), .B(KEYINPUT100), .Z(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n571_), .A2(new_n431_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT38), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT101), .ZN(new_n577_));
  INV_X1    g376(.A(new_n551_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n428_), .A2(new_n578_), .ZN(new_n579_));
  NOR3_X1   g378(.A1(new_n531_), .A2(new_n569_), .A3(new_n457_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n252_), .ZN(new_n582_));
  OAI21_X1  g381(.A(G1gat), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n577_), .B(new_n583_), .C1(new_n575_), .C2(new_n574_), .ZN(G1324gat));
  OR3_X1    g383(.A1(new_n581_), .A2(KEYINPUT102), .A3(new_n403_), .ZN(new_n585_));
  OAI21_X1  g384(.A(KEYINPUT102), .B1(new_n581_), .B2(new_n403_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(G8gat), .A3(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n588_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n403_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n571_), .A2(new_n432_), .A3(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n589_), .A2(new_n590_), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT40), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(G1325gat));
  OAI21_X1  g394(.A(G15gat), .B1(new_n581_), .B2(new_n360_), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n596_), .A2(KEYINPUT41), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(KEYINPUT41), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n571_), .A2(new_n305_), .A3(new_n362_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n597_), .A2(new_n598_), .A3(new_n599_), .ZN(G1326gat));
  INV_X1    g399(.A(new_n301_), .ZN(new_n601_));
  OAI21_X1  g400(.A(G22gat), .B1(new_n581_), .B2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT42), .ZN(new_n603_));
  INV_X1    g402(.A(new_n571_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n601_), .A2(G22gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT104), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n603_), .B1(new_n604_), .B2(new_n606_), .ZN(G1327gat));
  NOR2_X1   g406(.A1(new_n568_), .A2(new_n551_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n532_), .A2(new_n608_), .ZN(new_n609_));
  OR3_X1    g408(.A1(new_n609_), .A2(G29gat), .A3(new_n582_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT44), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n531_), .A2(new_n568_), .A3(new_n457_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n551_), .B(KEYINPUT37), .ZN(new_n614_));
  OAI211_X1 g413(.A(KEYINPUT105), .B(KEYINPUT43), .C1(new_n428_), .C2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n361_), .A2(new_n363_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n616_), .A2(new_n403_), .A3(new_n582_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n426_), .A2(new_n427_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n614_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT43), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n615_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT105), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n623_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n613_), .B1(new_n622_), .B2(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n611_), .B1(new_n625_), .B2(KEYINPUT106), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n624_), .A2(new_n615_), .A3(new_n621_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n612_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT106), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(new_n629_), .A3(KEYINPUT44), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n626_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT107), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n631_), .A2(new_n632_), .A3(new_n573_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(G29gat), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n632_), .B1(new_n631_), .B2(new_n573_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n610_), .B1(new_n634_), .B2(new_n635_), .ZN(G1328gat));
  INV_X1    g435(.A(new_n609_), .ZN(new_n637_));
  INV_X1    g436(.A(G36gat), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n637_), .A2(new_n638_), .A3(new_n591_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT45), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n403_), .B1(new_n626_), .B2(new_n630_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n640_), .B1(new_n641_), .B2(new_n638_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT46), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  OAI211_X1 g443(.A(KEYINPUT46), .B(new_n640_), .C1(new_n641_), .C2(new_n638_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(G1329gat));
  XOR2_X1   g445(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT44), .B1(new_n628_), .B2(new_n629_), .ZN(new_n648_));
  AOI211_X1 g447(.A(KEYINPUT106), .B(new_n611_), .C1(new_n627_), .C2(new_n612_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n362_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(G43gat), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n609_), .A2(G43gat), .A3(new_n360_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n647_), .B1(new_n651_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n647_), .ZN(new_n655_));
  AOI211_X1 g454(.A(new_n652_), .B(new_n655_), .C1(new_n650_), .C2(G43gat), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n654_), .A2(new_n656_), .ZN(G1330gat));
  AOI21_X1  g456(.A(G50gat), .B1(new_n637_), .B2(new_n301_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n301_), .A2(G50gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n631_), .B2(new_n659_), .ZN(G1331gat));
  AND2_X1   g459(.A1(new_n531_), .A2(new_n570_), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n661_), .A2(KEYINPUT109), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(KEYINPUT109), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n428_), .A2(new_n456_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n662_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n245_), .B1(new_n665_), .B2(new_n572_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT110), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n666_), .A2(new_n667_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n531_), .A2(new_n457_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n670_), .A2(new_n569_), .ZN(new_n671_));
  XOR2_X1   g470(.A(KEYINPUT111), .B(G57gat), .Z(new_n672_));
  NAND4_X1  g471(.A1(new_n671_), .A2(new_n579_), .A3(new_n252_), .A4(new_n672_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT112), .Z(new_n674_));
  NOR3_X1   g473(.A1(new_n668_), .A2(new_n669_), .A3(new_n674_), .ZN(G1332gat));
  NAND2_X1  g474(.A1(new_n671_), .A2(new_n579_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G64gat), .B1(new_n676_), .B2(new_n403_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT48), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n403_), .A2(G64gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n678_), .B1(new_n665_), .B2(new_n679_), .ZN(G1333gat));
  OAI21_X1  g479(.A(G71gat), .B1(new_n676_), .B2(new_n360_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT49), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n360_), .A2(G71gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n682_), .B1(new_n665_), .B2(new_n683_), .ZN(G1334gat));
  OAI21_X1  g483(.A(G78gat), .B1(new_n676_), .B2(new_n601_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT50), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n301_), .A2(new_n506_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n686_), .B1(new_n665_), .B2(new_n687_), .ZN(G1335gat));
  NOR4_X1   g487(.A1(new_n670_), .A2(new_n428_), .A3(new_n568_), .A4(new_n551_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(new_n247_), .A3(new_n573_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n670_), .A2(new_n568_), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n627_), .A2(new_n252_), .A3(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n690_), .B1(new_n692_), .B2(new_n247_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT113), .ZN(G1336gat));
  INV_X1    g493(.A(G92gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n689_), .A2(new_n695_), .A3(new_n591_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n627_), .A2(new_n591_), .A3(new_n691_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n696_), .B1(new_n697_), .B2(new_n695_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT114), .Z(G1337gat));
  NAND4_X1  g498(.A1(new_n689_), .A2(new_n490_), .A3(new_n492_), .A4(new_n362_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n627_), .A2(new_n362_), .A3(new_n691_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(G99gat), .B2(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(G1338gat));
  NAND3_X1  g505(.A1(new_n689_), .A2(new_n491_), .A3(new_n301_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT116), .Z(new_n708_));
  NAND3_X1  g507(.A1(new_n627_), .A2(new_n301_), .A3(new_n691_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(G106gat), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT52), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n709_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n708_), .A2(new_n712_), .A3(new_n713_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g514(.A1(new_n591_), .A2(new_n572_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n716_), .A2(new_n362_), .A3(new_n601_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n717_), .A2(KEYINPUT59), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n524_), .A2(new_n528_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n456_), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n520_), .A2(KEYINPUT12), .A3(new_n510_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT12), .B1(new_n520_), .B2(new_n510_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n520_), .A2(new_n510_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n721_), .A2(new_n722_), .A3(new_n723_), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n724_), .A2(KEYINPUT118), .A3(KEYINPUT55), .A4(new_n513_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT118), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT55), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n522_), .B2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n522_), .A2(new_n727_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n512_), .A2(new_n514_), .A3(new_n521_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n730_), .A2(G230gat), .A3(G233gat), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n725_), .A2(new_n728_), .A3(new_n729_), .A4(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n528_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT56), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n732_), .A2(KEYINPUT56), .A3(new_n528_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n720_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n429_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n738_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT119), .ZN(new_n740_));
  OR3_X1    g539(.A1(new_n739_), .A2(new_n740_), .A3(new_n454_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n740_), .B1(new_n739_), .B2(new_n454_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n447_), .A2(new_n738_), .A3(new_n440_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n741_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n744_), .A2(new_n455_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n529_), .A2(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n551_), .B1(new_n737_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT57), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n719_), .A2(new_n745_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n732_), .A2(KEYINPUT56), .A3(new_n528_), .ZN(new_n751_));
  AOI21_X1  g550(.A(KEYINPUT56), .B1(new_n732_), .B2(new_n528_), .ZN(new_n752_));
  OAI211_X1 g551(.A(KEYINPUT120), .B(new_n750_), .C1(new_n751_), .C2(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(KEYINPUT58), .B1(new_n753_), .B2(KEYINPUT121), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n735_), .A2(new_n736_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n756_));
  AOI22_X1  g555(.A1(new_n755_), .A2(new_n750_), .B1(KEYINPUT120), .B2(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n553_), .B1(new_n754_), .B2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n747_), .A2(new_n748_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT122), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n749_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n758_), .A2(KEYINPUT122), .A3(new_n759_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n568_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  XOR2_X1   g563(.A(KEYINPUT117), .B(KEYINPUT54), .Z(new_n765_));
  NAND3_X1  g564(.A1(new_n614_), .A2(new_n568_), .A3(new_n457_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n530_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n765_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n765_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n570_), .A2(new_n457_), .A3(new_n530_), .A4(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n718_), .B1(new_n764_), .B2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n749_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n773_), .A2(new_n758_), .A3(new_n759_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n771_), .B1(new_n774_), .B2(new_n569_), .ZN(new_n775_));
  OAI21_X1  g574(.A(KEYINPUT59), .B1(new_n775_), .B2(new_n717_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n772_), .A2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT123), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n760_), .A2(new_n761_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n780_), .A2(new_n773_), .A3(new_n763_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n771_), .B1(new_n781_), .B2(new_n569_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n718_), .ZN(new_n783_));
  OAI211_X1 g582(.A(KEYINPUT123), .B(new_n776_), .C1(new_n782_), .C2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n779_), .A2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(G113gat), .B1(new_n785_), .B2(new_n457_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n775_), .A2(new_n717_), .ZN(new_n787_));
  INV_X1    g586(.A(G113gat), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n788_), .A3(new_n456_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n786_), .A2(new_n789_), .ZN(G1340gat));
  INV_X1    g589(.A(KEYINPUT60), .ZN(new_n791_));
  INV_X1    g590(.A(G120gat), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n531_), .A2(new_n791_), .A3(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n793_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n787_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n772_), .A2(new_n531_), .A3(new_n776_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n795_), .B1(new_n797_), .B2(new_n792_), .ZN(G1341gat));
  OAI21_X1  g597(.A(G127gat), .B1(new_n785_), .B2(new_n569_), .ZN(new_n799_));
  INV_X1    g598(.A(G127gat), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n787_), .A2(new_n800_), .A3(new_n568_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(G1342gat));
  INV_X1    g601(.A(KEYINPUT124), .ZN(new_n803_));
  INV_X1    g602(.A(new_n784_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT123), .B1(new_n772_), .B2(new_n776_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n553_), .A2(G134gat), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n804_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n775_), .A2(new_n551_), .A3(new_n717_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n808_), .A2(G134gat), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n803_), .B1(new_n807_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n809_), .ZN(new_n811_));
  OAI211_X1 g610(.A(KEYINPUT124), .B(new_n811_), .C1(new_n785_), .C2(new_n806_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(G1343gat));
  NOR2_X1   g612(.A1(new_n775_), .A2(new_n361_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n716_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n456_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n531_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g619(.A1(new_n815_), .A2(new_n569_), .ZN(new_n821_));
  XOR2_X1   g620(.A(KEYINPUT61), .B(G155gat), .Z(new_n822_));
  XNOR2_X1  g621(.A(new_n821_), .B(new_n822_), .ZN(G1346gat));
  OR3_X1    g622(.A1(new_n815_), .A2(G162gat), .A3(new_n551_), .ZN(new_n824_));
  OAI21_X1  g623(.A(G162gat), .B1(new_n815_), .B2(new_n614_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(G1347gat));
  INV_X1    g625(.A(new_n782_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n572_), .A2(new_n362_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n828_), .A2(new_n403_), .A3(new_n301_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n827_), .A2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n830_), .A2(new_n456_), .A3(new_n333_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n827_), .A2(new_n456_), .A3(new_n829_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT62), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(new_n833_), .A3(G169gat), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n832_), .B2(G169gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n835_), .B2(KEYINPUT125), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT125), .ZN(new_n837_));
  AOI211_X1 g636(.A(new_n837_), .B(new_n833_), .C1(new_n832_), .C2(G169gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n831_), .B1(new_n836_), .B2(new_n838_), .ZN(G1348gat));
  AOI21_X1  g638(.A(G176gat), .B1(new_n830_), .B2(new_n531_), .ZN(new_n840_));
  NOR4_X1   g639(.A1(new_n775_), .A2(new_n403_), .A3(new_n301_), .A4(new_n828_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n531_), .A2(G176gat), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n840_), .B1(new_n841_), .B2(new_n842_), .ZN(G1349gat));
  AOI21_X1  g642(.A(G183gat), .B1(new_n841_), .B2(new_n568_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n568_), .A2(new_n371_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n844_), .B1(new_n830_), .B2(new_n845_), .ZN(G1350gat));
  INV_X1    g645(.A(new_n369_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n830_), .A2(new_n578_), .A3(new_n847_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n830_), .A2(new_n553_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(new_n318_), .ZN(G1351gat));
  NOR2_X1   g649(.A1(new_n403_), .A2(new_n252_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n814_), .A2(new_n851_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n852_), .A2(new_n457_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(new_n257_), .ZN(G1352gat));
  NAND3_X1  g653(.A1(new_n814_), .A2(new_n531_), .A3(new_n851_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  XOR2_X1   g656(.A(KEYINPUT126), .B(G204gat), .Z(new_n858_));
  AOI21_X1  g657(.A(new_n857_), .B1(new_n855_), .B2(new_n858_), .ZN(G1353gat));
  NOR2_X1   g658(.A1(new_n852_), .A2(new_n569_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n861_));
  AND2_X1   g660(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n860_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(new_n860_), .B2(new_n861_), .ZN(G1354gat));
  INV_X1    g663(.A(G218gat), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n852_), .A2(new_n865_), .A3(new_n614_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n852_), .A2(KEYINPUT127), .A3(new_n551_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(G218gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(KEYINPUT127), .B1(new_n852_), .B2(new_n551_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n866_), .B1(new_n868_), .B2(new_n869_), .ZN(G1355gat));
endmodule


