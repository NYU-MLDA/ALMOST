//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n886_, new_n888_,
    new_n889_, new_n890_, new_n891_, new_n892_, new_n893_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_;
  NOR2_X1   g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT87), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT1), .ZN(new_n205_));
  OR2_X1    g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT86), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT86), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(G141gat), .A3(G148gat), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(G141gat), .ZN(new_n212_));
  INV_X1    g011(.A(G148gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n206_), .A2(new_n211_), .A3(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n208_), .A2(new_n210_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT88), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n208_), .A2(new_n210_), .A3(KEYINPUT88), .A4(new_n216_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n212_), .A2(new_n213_), .A3(KEYINPUT3), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT3), .B1(new_n212_), .B2(new_n213_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n222_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n221_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT89), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n221_), .A2(KEYINPUT89), .A3(new_n226_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n203_), .B1(G155gat), .B2(G162gat), .ZN(new_n232_));
  AOI21_X1  g031(.A(KEYINPUT90), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  AOI211_X1 g032(.A(new_n228_), .B(new_n225_), .C1(new_n219_), .C2(new_n220_), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT89), .B1(new_n221_), .B2(new_n226_), .ZN(new_n235_));
  OAI211_X1 g034(.A(KEYINPUT90), .B(new_n232_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n215_), .B1(new_n233_), .B2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G127gat), .B(G134gat), .ZN(new_n239_));
  INV_X1    g038(.A(G113gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n239_), .B(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(G120gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n238_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G225gat), .A2(G233gat), .ZN(new_n246_));
  INV_X1    g045(.A(new_n215_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n232_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT90), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n247_), .B1(new_n250_), .B2(new_n236_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(new_n243_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n245_), .A2(new_n246_), .A3(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT0), .B(G57gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(G85gat), .ZN(new_n255_));
  XOR2_X1   g054(.A(G1gat), .B(G29gat), .Z(new_n256_));
  XOR2_X1   g055(.A(new_n255_), .B(new_n256_), .Z(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n250_), .A2(new_n236_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n243_), .B1(new_n259_), .B2(new_n215_), .ZN(new_n260_));
  AOI211_X1 g059(.A(new_n244_), .B(new_n247_), .C1(new_n250_), .C2(new_n236_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n262_));
  NOR3_X1   g061(.A1(new_n260_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n238_), .A2(new_n262_), .A3(new_n244_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n246_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n253_), .B(new_n258_), .C1(new_n263_), .C2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n245_), .A2(KEYINPUT4), .A3(new_n252_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n246_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n258_), .B1(new_n271_), .B2(new_n253_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n268_), .A2(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(KEYINPUT96), .B(KEYINPUT24), .Z(new_n274_));
  INV_X1    g073(.A(G169gat), .ZN(new_n275_));
  INV_X1    g074(.A(G176gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  OR2_X1    g076(.A1(new_n274_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G183gat), .A2(G190gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT23), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT82), .B(KEYINPUT23), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n280_), .B1(new_n281_), .B2(new_n279_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n274_), .A2(new_n277_), .A3(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT26), .B(G190gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT25), .B(G183gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n278_), .A2(new_n282_), .A3(new_n284_), .A4(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT97), .ZN(new_n289_));
  NOR2_X1   g088(.A1(G183gat), .A2(G190gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n281_), .A2(new_n279_), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n279_), .A2(KEYINPUT23), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n290_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n283_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT22), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(G169gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n275_), .A2(KEYINPUT22), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n297_), .A2(new_n298_), .A3(new_n276_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n289_), .B1(new_n295_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n299_), .ZN(new_n301_));
  NOR4_X1   g100(.A1(new_n293_), .A2(KEYINPUT97), .A3(new_n294_), .A4(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n288_), .B1(new_n300_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(G197gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(G204gat), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT92), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n304_), .A2(KEYINPUT92), .A3(G204gat), .ZN(new_n308_));
  INV_X1    g107(.A(G204gat), .ZN(new_n309_));
  AOI22_X1  g108(.A1(new_n307_), .A2(new_n308_), .B1(G197gat), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT93), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G211gat), .B(G218gat), .Z(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT21), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n316_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n313_), .B1(new_n310_), .B2(new_n316_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n309_), .A2(G197gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n319_), .A2(new_n305_), .A3(KEYINPUT91), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n320_), .B(KEYINPUT21), .C1(KEYINPUT91), .C2(new_n305_), .ZN(new_n321_));
  AOI22_X1  g120(.A1(new_n315_), .A2(new_n317_), .B1(new_n318_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n303_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT83), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n325_), .B1(new_n296_), .B2(G169gat), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n275_), .A2(KEYINPUT83), .A3(KEYINPUT22), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n326_), .A2(new_n327_), .A3(new_n276_), .A4(new_n297_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(new_n283_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT84), .ZN(new_n330_));
  INV_X1    g129(.A(new_n290_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n282_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT84), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n328_), .A2(new_n333_), .A3(new_n283_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n330_), .A2(new_n332_), .A3(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n291_), .A2(new_n292_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT26), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT81), .B1(new_n337_), .B2(G190gat), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n286_), .B(new_n338_), .C1(new_n285_), .C2(KEYINPUT81), .ZN(new_n339_));
  OR2_X1    g138(.A1(new_n277_), .A2(KEYINPUT24), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n277_), .A2(KEYINPUT24), .A3(new_n283_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n336_), .A2(new_n339_), .A3(new_n340_), .A4(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n335_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT85), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n335_), .A2(KEYINPUT85), .A3(new_n342_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(new_n346_), .A3(new_n322_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n324_), .A2(KEYINPUT20), .A3(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT95), .ZN(new_n350_));
  AND2_X1   g149(.A1(G226gat), .A2(G233gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n348_), .A2(new_n353_), .ZN(new_n354_));
  OR2_X1    g153(.A1(new_n303_), .A2(new_n323_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n346_), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT85), .B1(new_n335_), .B2(new_n342_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n323_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n355_), .A2(KEYINPUT20), .A3(new_n352_), .A4(new_n358_), .ZN(new_n359_));
  XOR2_X1   g158(.A(G8gat), .B(G36gat), .Z(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT99), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G64gat), .B(G92gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(KEYINPUT98), .B(KEYINPUT18), .Z(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n354_), .A2(new_n359_), .A3(new_n365_), .ZN(new_n366_));
  XOR2_X1   g165(.A(KEYINPUT102), .B(KEYINPUT20), .Z(new_n367_));
  NAND2_X1  g166(.A1(new_n295_), .A2(new_n299_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n322_), .A2(new_n288_), .A3(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n358_), .A2(new_n367_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n353_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n324_), .A2(new_n347_), .A3(KEYINPUT20), .A4(new_n352_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n365_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT27), .ZN(new_n374_));
  OR3_X1    g173(.A1(new_n366_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n365_), .B1(new_n354_), .B2(new_n359_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n374_), .B1(new_n366_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G78gat), .B(G106gat), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT29), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n382_), .B(new_n215_), .C1(new_n233_), .C2(new_n237_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G22gat), .B(G50gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT28), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n383_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n251_), .A2(new_n382_), .A3(new_n385_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n323_), .B1(new_n251_), .B2(new_n382_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G228gat), .A2(G233gat), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n391_), .B(new_n323_), .C1(new_n251_), .C2(new_n382_), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n389_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n389_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n381_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G15gat), .B(G43gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT31), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G227gat), .A2(G233gat), .ZN(new_n400_));
  XOR2_X1   g199(.A(new_n399_), .B(new_n400_), .Z(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT30), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n345_), .A2(new_n403_), .A3(new_n346_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n403_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n244_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G71gat), .B(G99gat), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n345_), .A2(new_n346_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT30), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(new_n404_), .A3(new_n243_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n407_), .A2(new_n409_), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n409_), .B1(new_n407_), .B2(new_n412_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n402_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NOR3_X1   g215(.A1(new_n405_), .A2(new_n244_), .A3(new_n406_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n243_), .B1(new_n411_), .B2(new_n404_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n408_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n419_), .A2(new_n413_), .A3(new_n401_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n416_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n393_), .A2(new_n394_), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n387_), .A2(new_n388_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n389_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n424_), .A2(new_n380_), .A3(new_n425_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n397_), .A2(new_n421_), .A3(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n421_), .B1(new_n397_), .B2(new_n426_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n273_), .B(new_n379_), .C1(new_n427_), .C2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT103), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n371_), .A2(new_n372_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n365_), .A2(KEYINPUT32), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n430_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n434_));
  AOI211_X1 g233(.A(KEYINPUT103), .B(new_n432_), .C1(new_n371_), .C2(new_n372_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(new_n432_), .B(KEYINPUT101), .Z(new_n437_));
  NAND3_X1  g236(.A1(new_n437_), .A2(new_n354_), .A3(new_n359_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n436_), .B(new_n438_), .C1(new_n268_), .C2(new_n272_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT100), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT33), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n267_), .A2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n366_), .A2(new_n376_), .ZN(new_n443_));
  XOR2_X1   g242(.A(KEYINPUT100), .B(KEYINPUT33), .Z(new_n444_));
  NAND4_X1  g243(.A1(new_n271_), .A2(new_n253_), .A3(new_n258_), .A4(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n269_), .A2(new_n246_), .A3(new_n264_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n245_), .A2(new_n265_), .A3(new_n252_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n446_), .A2(new_n257_), .A3(new_n447_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n442_), .A2(new_n443_), .A3(new_n445_), .A4(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n439_), .A2(new_n449_), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n416_), .A2(new_n420_), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n424_), .A2(new_n380_), .A3(new_n425_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n380_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n450_), .A2(new_n451_), .A3(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n429_), .A2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT73), .B(G134gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(G162gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G190gat), .B(G218gat), .ZN(new_n459_));
  XOR2_X1   g258(.A(new_n458_), .B(new_n459_), .Z(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G232gat), .A2(G233gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT34), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT70), .B(KEYINPUT35), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(G85gat), .B(G92gat), .Z(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT9), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT9), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(G85gat), .A3(G92gat), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT6), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n470_), .B1(G99gat), .B2(G106gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G99gat), .A2(G106gat), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n472_), .A2(KEYINPUT6), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n467_), .B(new_n469_), .C1(new_n471_), .C2(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(KEYINPUT10), .B(G99gat), .Z(new_n475_));
  XOR2_X1   g274(.A(KEYINPUT64), .B(G106gat), .Z(new_n476_));
  AND2_X1   g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n474_), .A2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT67), .B1(new_n471_), .B2(new_n473_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n472_), .A2(KEYINPUT6), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n470_), .A2(G99gat), .A3(G106gat), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT67), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n480_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n479_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(G99gat), .ZN(new_n485_));
  INV_X1    g284(.A(G106gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(new_n486_), .A3(KEYINPUT65), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT7), .ZN(new_n488_));
  NOR2_X1   g287(.A1(G99gat), .A2(G106gat), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT7), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(KEYINPUT65), .A3(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n488_), .A2(KEYINPUT66), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT66), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n489_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n489_), .A2(KEYINPUT65), .A3(new_n490_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n490_), .B1(new_n489_), .B2(KEYINPUT65), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n495_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n484_), .B1(new_n492_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n466_), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT8), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  AOI22_X1  g300(.A1(new_n498_), .A2(new_n492_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT8), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n466_), .A2(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n478_), .B1(new_n501_), .B2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G43gat), .B(G50gat), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(G29gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT71), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT71), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(G29gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(G36gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT71), .B(G29gat), .ZN(new_n515_));
  INV_X1    g314(.A(G36gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n508_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n514_), .A2(new_n517_), .A3(new_n508_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n465_), .B1(new_n506_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n463_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n464_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n498_), .A2(new_n492_), .ZN(new_n526_));
  AND3_X1   g325(.A1(new_n480_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n482_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n500_), .B1(new_n526_), .B2(new_n529_), .ZN(new_n530_));
  OAI22_X1  g329(.A1(new_n530_), .A2(new_n503_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n478_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n519_), .A2(KEYINPUT15), .A3(new_n520_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT15), .ZN(new_n535_));
  INV_X1    g334(.A(new_n520_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n535_), .B1(new_n536_), .B2(new_n518_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n534_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n533_), .A2(new_n539_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n522_), .A2(KEYINPUT72), .A3(new_n525_), .A4(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n525_), .A2(KEYINPUT72), .ZN(new_n542_));
  INV_X1    g341(.A(new_n525_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT72), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NOR3_X1   g344(.A1(new_n496_), .A2(new_n497_), .A3(new_n493_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n494_), .B1(new_n488_), .B2(new_n491_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n529_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n503_), .B1(new_n548_), .B2(new_n466_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n502_), .A2(new_n504_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n521_), .B(new_n532_), .C1(new_n549_), .C2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n465_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n538_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n542_), .B(new_n545_), .C1(new_n553_), .C2(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n461_), .B1(new_n541_), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT74), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n557_), .B1(new_n541_), .B2(new_n555_), .ZN(new_n558_));
  OAI22_X1  g357(.A1(KEYINPUT36), .A2(new_n556_), .B1(new_n558_), .B2(new_n460_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n555_), .ZN(new_n560_));
  NOR4_X1   g359(.A1(new_n553_), .A2(new_n554_), .A3(new_n544_), .A4(new_n543_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT74), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT36), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n562_), .A2(new_n563_), .A3(new_n461_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n559_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n456_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT104), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G15gat), .B(G22gat), .ZN(new_n570_));
  XOR2_X1   g369(.A(KEYINPUT75), .B(G8gat), .Z(new_n571_));
  INV_X1    g370(.A(KEYINPUT14), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n570_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(G1gat), .ZN(new_n574_));
  INV_X1    g373(.A(G1gat), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n570_), .A2(new_n572_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(G8gat), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(KEYINPUT79), .B1(new_n579_), .B2(new_n521_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(new_n521_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n582_), .A2(G229gat), .A3(G233gat), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n521_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n578_), .A2(new_n539_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G229gat), .A2(G233gat), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n587_), .B(KEYINPUT80), .Z(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n583_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G113gat), .B(G141gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(new_n275_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(new_n304_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n590_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n593_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n583_), .A2(new_n589_), .A3(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G57gat), .B(G64gat), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n598_), .A2(KEYINPUT11), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(KEYINPUT11), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G71gat), .B(G78gat), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n599_), .A2(new_n600_), .A3(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n603_), .B1(new_n600_), .B2(new_n602_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT68), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n533_), .A2(new_n605_), .A3(KEYINPUT12), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n506_), .A2(new_n604_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n506_), .A2(new_n604_), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n606_), .B(new_n607_), .C1(new_n608_), .C2(KEYINPUT12), .ZN(new_n609_));
  AND2_X1   g408(.A1(G230gat), .A2(G233gat), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n607_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n610_), .B1(new_n613_), .B2(new_n608_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G120gat), .B(G148gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(new_n309_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT5), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(new_n276_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT69), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n615_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n612_), .A2(new_n614_), .A3(new_n619_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT13), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G231gat), .A2(G233gat), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT76), .Z(new_n626_));
  XNOR2_X1  g425(.A(new_n578_), .B(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT77), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(new_n604_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(KEYINPUT16), .B(G183gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(G211gat), .ZN(new_n631_));
  XOR2_X1   g430(.A(G127gat), .B(G155gat), .Z(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT17), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT78), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n629_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT17), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n627_), .A2(new_n605_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n627_), .A2(new_n605_), .ZN(new_n639_));
  OR4_X1    g438(.A1(new_n637_), .A2(new_n638_), .A3(new_n639_), .A4(new_n633_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n636_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n569_), .A2(new_n597_), .A3(new_n624_), .A4(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G1gat), .B1(new_n643_), .B2(new_n273_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n565_), .A2(KEYINPUT37), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT37), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n559_), .A2(new_n564_), .A3(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n648_), .A2(new_n641_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n456_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n624_), .A2(new_n597_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n273_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(new_n575_), .A3(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT38), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n644_), .A2(new_n655_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT105), .Z(G1324gat));
  INV_X1    g456(.A(new_n571_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n652_), .A2(new_n658_), .A3(new_n378_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT39), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n643_), .A2(new_n379_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n661_), .B2(G8gat), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n660_), .B(G8gat), .C1(new_n643_), .C2(new_n379_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n659_), .B1(new_n662_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT40), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  OAI211_X1 g466(.A(KEYINPUT40), .B(new_n659_), .C1(new_n662_), .C2(new_n664_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1325gat));
  OAI21_X1  g468(.A(G15gat), .B1(new_n643_), .B2(new_n451_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT41), .Z(new_n671_));
  INV_X1    g470(.A(G15gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n652_), .A2(new_n672_), .A3(new_n421_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(G1326gat));
  OAI21_X1  g473(.A(G22gat), .B1(new_n643_), .B2(new_n454_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT42), .ZN(new_n676_));
  INV_X1    g475(.A(G22gat), .ZN(new_n677_));
  INV_X1    g476(.A(new_n454_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n652_), .A2(new_n677_), .A3(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n676_), .A2(new_n679_), .ZN(G1327gat));
  NOR2_X1   g479(.A1(new_n651_), .A2(new_n642_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n451_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n397_), .A2(new_n421_), .A3(new_n426_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n378_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n421_), .B1(new_n439_), .B2(new_n449_), .ZN(new_n686_));
  AOI22_X1  g485(.A1(new_n685_), .A2(new_n273_), .B1(new_n686_), .B2(new_n454_), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n682_), .A2(new_n566_), .A3(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(G29gat), .B1(new_n688_), .B2(new_n653_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n456_), .A2(new_n690_), .A3(new_n648_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n559_), .A2(new_n646_), .A3(new_n564_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n646_), .B1(new_n559_), .B2(new_n564_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n694_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n645_), .A2(KEYINPUT106), .A3(new_n647_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n699_), .B1(new_n429_), .B2(new_n455_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n693_), .B1(new_n700_), .B2(new_n690_), .ZN(new_n701_));
  OAI211_X1 g500(.A(KEYINPUT107), .B(KEYINPUT43), .C1(new_n687_), .C2(new_n699_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n692_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n703_), .A2(new_n682_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT44), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n705_), .A2(new_n273_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n689_), .B1(new_n706_), .B2(G29gat), .ZN(G1328gat));
  OAI21_X1  g506(.A(G36gat), .B1(new_n705_), .B2(new_n379_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n378_), .B(KEYINPUT108), .Z(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n688_), .A2(new_n516_), .A3(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT45), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n708_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT46), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n708_), .A2(KEYINPUT46), .A3(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1329gat));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n704_), .B(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n719_), .A2(G43gat), .A3(new_n421_), .ZN(new_n720_));
  INV_X1    g519(.A(G43gat), .ZN(new_n721_));
  INV_X1    g520(.A(new_n688_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n722_), .B2(new_n451_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n720_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT47), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n720_), .A2(new_n726_), .A3(new_n723_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(G1330gat));
  NAND3_X1  g527(.A1(new_n719_), .A2(G50gat), .A3(new_n678_), .ZN(new_n729_));
  INV_X1    g528(.A(G50gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n730_), .B1(new_n722_), .B2(new_n454_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n729_), .A2(KEYINPUT109), .A3(new_n731_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1331gat));
  NOR3_X1   g535(.A1(new_n650_), .A2(new_n597_), .A3(new_n624_), .ZN(new_n737_));
  AOI21_X1  g536(.A(G57gat), .B1(new_n737_), .B2(new_n653_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n624_), .A2(new_n597_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n569_), .A2(new_n642_), .A3(new_n739_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n740_), .A2(new_n273_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n738_), .B1(new_n741_), .B2(G57gat), .ZN(G1332gat));
  OAI21_X1  g541(.A(G64gat), .B1(new_n740_), .B2(new_n709_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT48), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n709_), .A2(G64gat), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT110), .Z(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(new_n737_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n744_), .A2(new_n747_), .ZN(G1333gat));
  OAI21_X1  g547(.A(G71gat), .B1(new_n740_), .B2(new_n451_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT49), .ZN(new_n750_));
  INV_X1    g549(.A(G71gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n737_), .A2(new_n751_), .A3(new_n421_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1334gat));
  OAI21_X1  g552(.A(G78gat), .B1(new_n740_), .B2(new_n454_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT50), .ZN(new_n755_));
  INV_X1    g554(.A(G78gat), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n737_), .A2(new_n756_), .A3(new_n678_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n755_), .A2(new_n757_), .ZN(G1335gat));
  NAND2_X1  g557(.A1(new_n739_), .A2(new_n641_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n759_), .A2(new_n687_), .A3(new_n566_), .ZN(new_n760_));
  AOI21_X1  g559(.A(G85gat), .B1(new_n760_), .B2(new_n653_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n701_), .A2(new_n702_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n759_), .B1(new_n762_), .B2(new_n691_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n764_), .A2(new_n273_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n761_), .B1(new_n765_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g565(.A(G92gat), .B1(new_n760_), .B2(new_n378_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n763_), .A2(G92gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(new_n710_), .ZN(G1337gat));
  OAI21_X1  g568(.A(G99gat), .B1(new_n764_), .B2(new_n451_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n760_), .A2(new_n475_), .A3(new_n421_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g572(.A(KEYINPUT112), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n486_), .B1(new_n763_), .B2(new_n678_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n774_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n699_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n456_), .A2(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT107), .B1(new_n779_), .B2(KEYINPUT43), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n700_), .A2(new_n693_), .A3(new_n690_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n691_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n759_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(new_n678_), .A3(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n784_), .A2(new_n776_), .A3(G106gat), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT111), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT111), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n775_), .A2(new_n787_), .A3(new_n776_), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n703_), .A2(new_n454_), .A3(new_n759_), .ZN(new_n789_));
  OAI211_X1 g588(.A(KEYINPUT112), .B(KEYINPUT52), .C1(new_n789_), .C2(new_n486_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n777_), .A2(new_n786_), .A3(new_n788_), .A4(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n760_), .A2(new_n476_), .A3(new_n678_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT53), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n791_), .A2(new_n795_), .A3(new_n792_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(G1339gat));
  INV_X1    g596(.A(new_n597_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n649_), .A2(new_n624_), .A3(new_n798_), .ZN(new_n799_));
  XOR2_X1   g598(.A(new_n799_), .B(KEYINPUT54), .Z(new_n800_));
  INV_X1    g599(.A(KEYINPUT57), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n582_), .A2(new_n588_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n586_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n802_), .B(new_n593_), .C1(new_n803_), .C2(new_n588_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n804_), .A2(new_n596_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n805_), .A2(new_n623_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n808_), .A2(new_n611_), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n609_), .A2(new_n807_), .A3(new_n610_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n620_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT56), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT113), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n597_), .B(new_n622_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n811_), .A2(new_n812_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n817_), .A2(KEYINPUT113), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n813_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n806_), .B1(new_n816_), .B2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n801_), .B1(new_n820_), .B2(new_n565_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n811_), .B(new_n812_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n822_), .A2(new_n622_), .A3(new_n805_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT58), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n824_), .A2(KEYINPUT114), .ZN(new_n825_));
  OR2_X1    g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n823_), .A2(new_n825_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n648_), .A3(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n815_), .B1(new_n813_), .B2(new_n818_), .ZN(new_n829_));
  OAI211_X1 g628(.A(KEYINPUT57), .B(new_n566_), .C1(new_n829_), .C2(new_n806_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n821_), .A2(new_n828_), .A3(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n800_), .B1(new_n831_), .B2(new_n641_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n832_), .A2(new_n678_), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n378_), .A2(new_n273_), .A3(new_n451_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT116), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n833_), .A2(new_n838_), .A3(KEYINPUT59), .A4(new_n834_), .ZN(new_n839_));
  AOI22_X1  g638(.A1(new_n837_), .A2(new_n839_), .B1(KEYINPUT117), .B2(new_n240_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n841_));
  OAI21_X1  g640(.A(G113gat), .B1(new_n798_), .B2(new_n841_), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n833_), .A2(KEYINPUT115), .A3(new_n834_), .ZN(new_n843_));
  AOI21_X1  g642(.A(KEYINPUT115), .B1(new_n833_), .B2(new_n834_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n597_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n840_), .A2(new_n842_), .B1(new_n845_), .B2(new_n240_), .ZN(G1340gat));
  OAI21_X1  g645(.A(new_n242_), .B1(new_n624_), .B2(KEYINPUT60), .ZN(new_n847_));
  OAI221_X1 g646(.A(new_n847_), .B1(KEYINPUT60), .B2(new_n242_), .C1(new_n843_), .C2(new_n844_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n624_), .B1(new_n837_), .B2(new_n839_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(new_n242_), .ZN(G1341gat));
  INV_X1    g649(.A(G127gat), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n851_), .B1(new_n837_), .B2(new_n839_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n642_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n853_));
  AOI22_X1  g652(.A1(new_n852_), .A2(new_n642_), .B1(new_n853_), .B2(new_n851_), .ZN(G1342gat));
  AOI22_X1  g653(.A1(new_n837_), .A2(new_n839_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n855_));
  XOR2_X1   g654(.A(KEYINPUT118), .B(G134gat), .Z(new_n856_));
  OAI21_X1  g655(.A(new_n565_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n857_));
  INV_X1    g656(.A(G134gat), .ZN(new_n858_));
  AOI22_X1  g657(.A1(new_n855_), .A2(new_n856_), .B1(new_n857_), .B2(new_n858_), .ZN(G1343gat));
  NOR3_X1   g658(.A1(new_n832_), .A2(new_n273_), .A3(new_n683_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n709_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(new_n798_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(new_n212_), .ZN(G1344gat));
  NOR2_X1   g662(.A1(new_n861_), .A2(new_n624_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(new_n213_), .ZN(G1345gat));
  NOR2_X1   g664(.A1(new_n861_), .A2(new_n641_), .ZN(new_n866_));
  XOR2_X1   g665(.A(KEYINPUT61), .B(G155gat), .Z(new_n867_));
  XNOR2_X1  g666(.A(new_n866_), .B(new_n867_), .ZN(G1346gat));
  INV_X1    g667(.A(new_n861_), .ZN(new_n869_));
  AND3_X1   g668(.A1(new_n869_), .A2(G162gat), .A3(new_n778_), .ZN(new_n870_));
  AOI21_X1  g669(.A(G162gat), .B1(new_n869_), .B2(new_n565_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1347gat));
  INV_X1    g671(.A(KEYINPUT62), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n709_), .A2(new_n653_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n421_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(KEYINPUT119), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n833_), .A2(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(new_n798_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n873_), .B1(new_n878_), .B2(new_n275_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n878_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n880_));
  OAI211_X1 g679(.A(KEYINPUT62), .B(G169gat), .C1(new_n877_), .C2(new_n798_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n879_), .A2(new_n880_), .A3(new_n881_), .ZN(G1348gat));
  NOR2_X1   g681(.A1(new_n877_), .A2(new_n624_), .ZN(new_n883_));
  XOR2_X1   g682(.A(KEYINPUT120), .B(G176gat), .Z(new_n884_));
  XNOR2_X1  g683(.A(new_n883_), .B(new_n884_), .ZN(G1349gat));
  NOR2_X1   g684(.A1(new_n877_), .A2(new_n641_), .ZN(new_n886_));
  MUX2_X1   g685(.A(G183gat), .B(new_n286_), .S(new_n886_), .Z(G1350gat));
  INV_X1    g686(.A(new_n648_), .ZN(new_n888_));
  OAI21_X1  g687(.A(G190gat), .B1(new_n877_), .B2(new_n888_), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n889_), .A2(KEYINPUT121), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n889_), .A2(KEYINPUT121), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n565_), .A2(new_n285_), .ZN(new_n892_));
  XOR2_X1   g691(.A(new_n892_), .B(KEYINPUT122), .Z(new_n893_));
  OAI22_X1  g692(.A1(new_n890_), .A2(new_n891_), .B1(new_n877_), .B2(new_n893_), .ZN(G1351gat));
  INV_X1    g693(.A(new_n874_), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n832_), .A2(new_n683_), .A3(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n597_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(KEYINPUT123), .B(G197gat), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n897_), .B(new_n898_), .ZN(G1352gat));
  INV_X1    g698(.A(new_n624_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n896_), .A2(new_n900_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g701(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n642_), .A2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(KEYINPUT124), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  NOR4_X1   g705(.A1(new_n832_), .A2(new_n683_), .A3(new_n895_), .A4(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT125), .ZN(new_n908_));
  OR2_X1    g707(.A1(new_n904_), .A2(KEYINPUT124), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n907_), .A2(new_n908_), .A3(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n908_), .B1(new_n907_), .B2(new_n909_), .ZN(new_n912_));
  OAI22_X1  g711(.A1(new_n911_), .A2(new_n912_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n913_));
  INV_X1    g712(.A(new_n912_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n914_), .A2(new_n915_), .A3(new_n910_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n913_), .A2(new_n916_), .ZN(G1354gat));
  AOI21_X1  g716(.A(G218gat), .B1(new_n896_), .B2(new_n565_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n648_), .A2(G218gat), .ZN(new_n919_));
  XOR2_X1   g718(.A(new_n919_), .B(KEYINPUT126), .Z(new_n920_));
  AOI21_X1  g719(.A(new_n918_), .B1(new_n896_), .B2(new_n920_), .ZN(G1355gat));
endmodule


