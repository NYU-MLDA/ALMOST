//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0 1 1 0 0 1 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1 0 0 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0 1 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n881_, new_n882_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n908_, new_n909_, new_n910_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n932_;
  INV_X1    g000(.A(KEYINPUT23), .ZN(new_n202_));
  NAND3_X1  g001(.A1(new_n202_), .A2(G183gat), .A3(G190gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n203_), .A2(KEYINPUT80), .ZN(new_n204_));
  INV_X1    g003(.A(G183gat), .ZN(new_n205_));
  INV_X1    g004(.A(G190gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT23), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(KEYINPUT80), .A3(new_n203_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n205_), .A2(new_n206_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n204_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(KEYINPUT79), .A2(G169gat), .ZN(new_n213_));
  AOI21_X1  g012(.A(G176gat), .B1(new_n213_), .B2(KEYINPUT22), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT22), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(KEYINPUT79), .A3(G169gat), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n212_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n210_), .A2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT25), .B(G183gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT26), .B(G190gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n207_), .A2(new_n203_), .ZN(new_n222_));
  INV_X1    g021(.A(G169gat), .ZN(new_n223_));
  INV_X1    g022(.A(G176gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n225_), .A2(KEYINPUT24), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(KEYINPUT24), .A3(new_n211_), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n221_), .A2(new_n222_), .A3(new_n226_), .A4(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n218_), .A2(KEYINPUT81), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT81), .B1(new_n218_), .B2(new_n228_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT30), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT83), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G227gat), .A2(G233gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT82), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G15gat), .B(G43gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G71gat), .B(G99gat), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n239_), .B(new_n240_), .Z(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n235_), .A2(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n242_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  XOR2_X1   g044(.A(G127gat), .B(G134gat), .Z(new_n246_));
  XOR2_X1   g045(.A(G113gat), .B(G120gat), .Z(new_n247_));
  XOR2_X1   g046(.A(new_n246_), .B(new_n247_), .Z(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT31), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n243_), .A2(new_n245_), .A3(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n249_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(G141gat), .A2(G148gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT85), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT85), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n257_), .B1(G141gat), .B2(G148gat), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT3), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n256_), .A2(KEYINPUT86), .A3(new_n258_), .A4(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G141gat), .A2(G148gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT2), .ZN(new_n262_));
  OAI22_X1  g061(.A1(new_n255_), .A2(new_n259_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT84), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n261_), .B(new_n265_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n260_), .B(new_n264_), .C1(new_n266_), .C2(KEYINPUT2), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n258_), .A2(new_n259_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT86), .B1(new_n269_), .B2(new_n256_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT87), .B1(new_n267_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G155gat), .A2(G162gat), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(G155gat), .A2(G162gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n261_), .B(KEYINPUT84), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n263_), .B1(new_n276_), .B2(new_n262_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT87), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT86), .ZN(new_n279_));
  INV_X1    g078(.A(new_n256_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n279_), .B1(new_n280_), .B2(new_n268_), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n277_), .A2(new_n278_), .A3(new_n281_), .A4(new_n260_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n271_), .A2(new_n275_), .A3(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n255_), .B1(new_n273_), .B2(KEYINPUT1), .ZN(new_n284_));
  INV_X1    g083(.A(new_n275_), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n276_), .B(new_n284_), .C1(new_n285_), .C2(KEYINPUT1), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n283_), .A2(new_n286_), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n287_), .A2(KEYINPUT29), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT28), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n287_), .A2(KEYINPUT29), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT28), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G22gat), .B(G50gat), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n289_), .A2(new_n292_), .A3(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n294_), .B1(new_n289_), .B2(new_n292_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(G233gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT88), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n299_), .A2(G228gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(G228gat), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n298_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT89), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(G78gat), .ZN(new_n304_));
  INV_X1    g103(.A(G106gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n287_), .A2(KEYINPUT29), .ZN(new_n307_));
  NOR2_X1   g106(.A1(G197gat), .A2(G204gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT91), .B(G197gat), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n308_), .B1(new_n309_), .B2(G204gat), .ZN(new_n310_));
  OR2_X1    g109(.A1(new_n310_), .A2(KEYINPUT21), .ZN(new_n311_));
  XOR2_X1   g110(.A(G211gat), .B(G218gat), .Z(new_n312_));
  OR2_X1    g111(.A1(new_n309_), .A2(G204gat), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT21), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n314_), .B1(G197gat), .B2(G204gat), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n312_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n312_), .A2(KEYINPUT21), .ZN(new_n317_));
  AOI22_X1  g116(.A1(new_n311_), .A2(new_n316_), .B1(new_n310_), .B2(new_n317_), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n318_), .A2(KEYINPUT90), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n306_), .B1(new_n307_), .B2(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n307_), .A2(new_n319_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n304_), .B(G106gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n295_), .A2(new_n297_), .A3(new_n320_), .A4(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n320_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n295_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n325_), .B1(new_n326_), .B2(new_n296_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n324_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT99), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G226gat), .A2(G233gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT19), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n222_), .A2(new_n209_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT22), .B(G169gat), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n212_), .B1(new_n334_), .B2(new_n224_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT94), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n221_), .A2(new_n227_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT92), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n204_), .A2(new_n208_), .A3(new_n226_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT92), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n221_), .A2(new_n341_), .A3(new_n227_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n339_), .A2(new_n340_), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT93), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n339_), .A2(new_n340_), .A3(KEYINPUT93), .A4(new_n342_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n337_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n332_), .B1(new_n347_), .B2(new_n318_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n311_), .A2(new_n316_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n317_), .A2(new_n310_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n351_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n348_), .A2(KEYINPUT20), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n231_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n354_), .A2(new_n318_), .A3(new_n229_), .ZN(new_n355_));
  OAI211_X1 g154(.A(KEYINPUT20), .B(new_n355_), .C1(new_n347_), .C2(new_n318_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n332_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G8gat), .B(G36gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT18), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G64gat), .B(G92gat), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n359_), .B(new_n360_), .Z(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT32), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n353_), .A2(new_n357_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n318_), .A2(new_n343_), .A3(new_n336_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n352_), .A2(KEYINPUT20), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(new_n332_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n367_), .B1(new_n356_), .B2(new_n332_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT98), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n345_), .A2(new_n346_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n351_), .B1(new_n370_), .B2(new_n337_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n332_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n371_), .A2(KEYINPUT20), .A3(new_n372_), .A4(new_n355_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT98), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n369_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n362_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n364_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G1gat), .B(G29gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(G85gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(KEYINPUT0), .B(G57gat), .ZN(new_n381_));
  XOR2_X1   g180(.A(new_n380_), .B(new_n381_), .Z(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT4), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT95), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n283_), .A2(new_n385_), .A3(new_n286_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n248_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n283_), .A2(new_n385_), .A3(new_n286_), .A4(new_n248_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n384_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G225gat), .A2(G233gat), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n287_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n248_), .A2(new_n384_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n392_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n390_), .A2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n392_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n383_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n388_), .A2(new_n389_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n391_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n400_), .B(new_n382_), .C1(new_n390_), .C2(new_n395_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n398_), .A2(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n330_), .B1(new_n378_), .B2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n374_), .B1(new_n373_), .B2(new_n367_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n356_), .ZN(new_n405_));
  AOI21_X1  g204(.A(KEYINPUT98), .B1(new_n405_), .B2(new_n372_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n377_), .B1(new_n404_), .B2(new_n406_), .ZN(new_n407_));
  AND4_X1   g206(.A1(new_n330_), .A2(new_n402_), .A3(new_n407_), .A4(new_n363_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n403_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n401_), .A2(KEYINPUT33), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n399_), .A2(KEYINPUT4), .ZN(new_n411_));
  INV_X1    g210(.A(new_n395_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT33), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n413_), .A2(new_n414_), .A3(new_n400_), .A4(new_n382_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n410_), .A2(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n391_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT96), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n411_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT96), .B1(new_n390_), .B2(new_n417_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n382_), .B1(new_n399_), .B2(new_n392_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n420_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n361_), .B1(new_n353_), .B2(new_n357_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n353_), .A2(new_n357_), .A3(new_n361_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n423_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT97), .B1(new_n416_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n410_), .A2(new_n415_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n426_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n430_), .A2(new_n424_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT97), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n429_), .A2(new_n431_), .A3(new_n432_), .A4(new_n423_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n428_), .A2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n329_), .B1(new_n409_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT27), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n436_), .B1(new_n430_), .B2(new_n424_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n361_), .B1(new_n369_), .B2(new_n375_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n426_), .A2(KEYINPUT27), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n437_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n328_), .A2(new_n402_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n441_), .A2(new_n442_), .A3(KEYINPUT100), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT100), .ZN(new_n444_));
  INV_X1    g243(.A(new_n402_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(new_n324_), .A3(new_n327_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n444_), .B1(new_n446_), .B2(new_n440_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n443_), .A2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n254_), .B1(new_n435_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n253_), .A2(new_n445_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n441_), .A2(new_n328_), .ZN(new_n451_));
  OR2_X1    g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n449_), .A2(new_n452_), .ZN(new_n453_));
  XOR2_X1   g252(.A(G29gat), .B(G36gat), .Z(new_n454_));
  XOR2_X1   g253(.A(G43gat), .B(G50gat), .Z(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT15), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G15gat), .B(G22gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G1gat), .A2(G8gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT14), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G1gat), .B(G8gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n457_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n456_), .ZN(new_n465_));
  OR2_X1    g264(.A1(new_n465_), .A2(new_n463_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G229gat), .A2(G233gat), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n464_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n465_), .B(new_n463_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n467_), .ZN(new_n470_));
  AND3_X1   g269(.A1(new_n469_), .A2(KEYINPUT77), .A3(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT77), .B1(new_n469_), .B2(new_n470_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n468_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G113gat), .B(G141gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G169gat), .B(G197gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n474_), .B(new_n475_), .Z(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n473_), .A2(new_n477_), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n468_), .B(new_n476_), .C1(new_n471_), .C2(new_n472_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n478_), .A2(KEYINPUT78), .A3(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT78), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n473_), .A2(new_n481_), .A3(new_n477_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n453_), .A2(KEYINPUT101), .A3(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT101), .B1(new_n453_), .B2(new_n484_), .ZN(new_n486_));
  OR2_X1    g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n488_));
  XOR2_X1   g287(.A(KEYINPUT65), .B(G92gat), .Z(new_n489_));
  INV_X1    g288(.A(G85gat), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n488_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G85gat), .B(G92gat), .ZN(new_n492_));
  INV_X1    g291(.A(G92gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n492_), .B1(KEYINPUT9), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n491_), .A2(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(KEYINPUT10), .B(G99gat), .Z(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(new_n305_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G99gat), .A2(G106gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT6), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n495_), .A2(new_n497_), .A3(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT8), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT68), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT67), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n506_), .A2(KEYINPUT6), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT6), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n508_), .A2(KEYINPUT67), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n498_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT7), .ZN(new_n511_));
  INV_X1    g310(.A(G99gat), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n512_), .A3(new_n305_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT68), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(new_n514_), .A3(new_n502_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n508_), .A2(KEYINPUT67), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n506_), .A2(KEYINPUT6), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n516_), .A2(new_n517_), .A3(G99gat), .A4(G106gat), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n505_), .A2(new_n510_), .A3(new_n515_), .A4(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n492_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n501_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  XOR2_X1   g320(.A(KEYINPUT66), .B(KEYINPUT8), .Z(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n503_), .A2(new_n504_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n523_), .B1(new_n499_), .B2(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n500_), .B1(new_n521_), .B2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G57gat), .B(G64gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT11), .ZN(new_n528_));
  XOR2_X1   g327(.A(G71gat), .B(G78gat), .Z(new_n529_));
  OR2_X1    g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n527_), .A2(KEYINPUT11), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n528_), .A2(new_n529_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n530_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n526_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT12), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n500_), .B(new_n533_), .C1(new_n521_), .C2(new_n525_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G230gat), .A2(G233gat), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n500_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n519_), .A2(new_n520_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT8), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT69), .ZN(new_n544_));
  INV_X1    g343(.A(new_n525_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n543_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT69), .B1(new_n521_), .B2(new_n525_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n541_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n534_), .A2(KEYINPUT12), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n537_), .B(new_n540_), .C1(new_n548_), .C2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT70), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n544_), .B1(new_n543_), .B2(new_n545_), .ZN(new_n552_));
  NOR3_X1   g351(.A1(new_n521_), .A2(KEYINPUT69), .A3(new_n525_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n500_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n549_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT70), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n556_), .A2(new_n557_), .A3(new_n537_), .A4(new_n540_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n535_), .A2(new_n538_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n539_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n551_), .A2(new_n558_), .A3(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G120gat), .B(G148gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT5), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G176gat), .B(G204gat), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n564_), .B(new_n565_), .Z(new_n566_));
  NAND2_X1  g365(.A1(new_n562_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n566_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n551_), .A2(new_n558_), .A3(new_n561_), .A4(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT13), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT71), .ZN(new_n573_));
  AOI21_X1  g372(.A(KEYINPUT13), .B1(new_n567_), .B2(new_n569_), .ZN(new_n574_));
  OR3_X1    g373(.A1(new_n572_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n573_), .B1(new_n572_), .B2(new_n574_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT34), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT35), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(KEYINPUT35), .ZN(new_n581_));
  INV_X1    g380(.A(new_n526_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n581_), .B1(new_n582_), .B2(new_n456_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT72), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n580_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n457_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n583_), .B1(new_n586_), .B2(new_n548_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  OAI221_X1 g387(.A(new_n583_), .B1(new_n584_), .B2(new_n580_), .C1(new_n586_), .C2(new_n548_), .ZN(new_n589_));
  XOR2_X1   g388(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n590_));
  NAND3_X1  g389(.A1(new_n588_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT74), .B(KEYINPUT36), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n592_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G190gat), .B(G218gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G134gat), .B(G162gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n593_), .A2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n593_), .A2(new_n596_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n591_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT37), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT37), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n601_), .B(new_n591_), .C1(new_n597_), .C2(new_n598_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G231gat), .A2(G233gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n463_), .B(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(new_n534_), .ZN(new_n606_));
  XOR2_X1   g405(.A(G127gat), .B(G155gat), .Z(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT16), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G183gat), .B(G211gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT17), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n606_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT75), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n610_), .B(KEYINPUT17), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n615_), .A2(KEYINPUT76), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n615_), .A2(KEYINPUT76), .ZN(new_n617_));
  OR3_X1    g416(.A1(new_n616_), .A2(new_n617_), .A3(new_n606_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n614_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n577_), .A2(new_n603_), .A3(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n487_), .A2(KEYINPUT102), .A3(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n621_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT102), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n445_), .A2(G1gat), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n622_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT38), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n622_), .A2(KEYINPUT38), .A3(new_n625_), .A4(new_n626_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n599_), .B(KEYINPUT103), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT104), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n453_), .A2(new_n632_), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n577_), .A2(new_n483_), .A3(new_n620_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(G1gat), .B1(new_n635_), .B2(new_n445_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n629_), .A2(new_n630_), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT105), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n629_), .A2(KEYINPUT105), .A3(new_n630_), .A4(new_n636_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1324gat));
  INV_X1    g440(.A(new_n635_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(new_n440_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(G8gat), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT39), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n643_), .A2(new_n646_), .A3(G8gat), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n441_), .A2(G8gat), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n622_), .A2(new_n625_), .A3(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n648_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n651_), .B1(new_n648_), .B2(new_n650_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1325gat));
  OAI21_X1  g453(.A(G15gat), .B1(new_n635_), .B2(new_n254_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT41), .Z(new_n656_));
  OR3_X1    g455(.A1(new_n623_), .A2(G15gat), .A3(new_n254_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1326gat));
  XNOR2_X1  g457(.A(new_n328_), .B(KEYINPUT107), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(G22gat), .B1(new_n635_), .B2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT42), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n660_), .A2(G22gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n662_), .B1(new_n623_), .B2(new_n663_), .ZN(G1327gat));
  NOR3_X1   g463(.A1(new_n577_), .A2(new_n631_), .A3(new_n619_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n487_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(G29gat), .B1(new_n667_), .B2(new_n402_), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n577_), .A2(new_n483_), .A3(new_n619_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT43), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n670_), .B1(new_n453_), .B2(new_n603_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n603_), .ZN(new_n672_));
  AOI211_X1 g471(.A(KEYINPUT43), .B(new_n672_), .C1(new_n449_), .C2(new_n452_), .ZN(new_n673_));
  OAI211_X1 g472(.A(KEYINPUT44), .B(new_n669_), .C1(new_n671_), .C2(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT108), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n671_), .A2(new_n673_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(new_n669_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n675_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n402_), .A2(G29gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n668_), .B1(new_n681_), .B2(new_n682_), .ZN(G1328gat));
  INV_X1    g482(.A(G36gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n441_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n675_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT46), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n441_), .A2(G36gat), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n665_), .B(new_n688_), .C1(new_n485_), .C2(new_n486_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT45), .Z(new_n690_));
  OR3_X1    g489(.A1(new_n686_), .A2(new_n687_), .A3(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n687_), .B1(new_n686_), .B2(new_n690_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1329gat));
  NAND4_X1  g492(.A1(new_n675_), .A2(G43gat), .A3(new_n253_), .A4(new_n679_), .ZN(new_n694_));
  INV_X1    g493(.A(G43gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n695_), .B1(new_n666_), .B2(new_n254_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n694_), .A2(new_n696_), .A3(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n694_), .B2(new_n696_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1330gat));
  INV_X1    g499(.A(G50gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n701_), .B1(new_n666_), .B2(new_n660_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n329_), .A2(G50gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n680_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT110), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  OAI211_X1 g505(.A(KEYINPUT110), .B(new_n702_), .C1(new_n680_), .C2(new_n703_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1331gat));
  INV_X1    g507(.A(new_n577_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n709_), .A2(new_n484_), .A3(new_n620_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n633_), .A2(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(G57gat), .B1(new_n711_), .B2(new_n445_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n603_), .A2(new_n620_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(new_n577_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT111), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n484_), .B1(new_n449_), .B2(new_n452_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  OR2_X1    g516(.A1(new_n445_), .A2(G57gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n712_), .B1(new_n717_), .B2(new_n718_), .ZN(G1332gat));
  OAI21_X1  g518(.A(G64gat), .B1(new_n711_), .B2(new_n441_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT48), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n441_), .A2(G64gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n717_), .B2(new_n722_), .ZN(G1333gat));
  OAI21_X1  g522(.A(G71gat), .B1(new_n711_), .B2(new_n254_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT49), .ZN(new_n725_));
  OR3_X1    g524(.A1(new_n717_), .A2(G71gat), .A3(new_n254_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT112), .ZN(G1334gat));
  OAI21_X1  g527(.A(G78gat), .B1(new_n711_), .B2(new_n660_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT50), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n660_), .A2(G78gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n717_), .B2(new_n731_), .ZN(G1335gat));
  XOR2_X1   g531(.A(new_n599_), .B(KEYINPUT103), .Z(new_n733_));
  AND4_X1   g532(.A1(new_n577_), .A2(new_n716_), .A3(new_n620_), .A4(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(new_n490_), .A3(new_n402_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n709_), .A2(new_n484_), .A3(new_n619_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n676_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n402_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n739_), .B2(new_n490_), .ZN(G1336gat));
  AOI21_X1  g539(.A(G92gat), .B1(new_n734_), .B2(new_n440_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n441_), .A2(new_n489_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n737_), .B2(new_n742_), .ZN(G1337gat));
  AOI21_X1  g542(.A(new_n512_), .B1(new_n737_), .B2(new_n253_), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n734_), .A2(new_n253_), .A3(new_n496_), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g546(.A1(new_n734_), .A2(new_n305_), .A3(new_n329_), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n329_), .B(new_n736_), .C1(new_n671_), .C2(new_n673_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(G106gat), .ZN(new_n750_));
  AOI21_X1  g549(.A(KEYINPUT114), .B1(new_n750_), .B2(KEYINPUT52), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT114), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT52), .ZN(new_n753_));
  AOI211_X1 g552(.A(new_n752_), .B(new_n753_), .C1(new_n749_), .C2(G106gat), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n751_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT113), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n756_), .B1(new_n750_), .B2(KEYINPUT52), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n749_), .A2(KEYINPUT113), .A3(new_n753_), .A4(G106gat), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n748_), .B1(new_n755_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT53), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n762_), .B(new_n748_), .C1(new_n755_), .C2(new_n759_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1339gat));
  INV_X1    g563(.A(KEYINPUT121), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n253_), .A2(new_n402_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n766_), .A2(new_n451_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n550_), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n537_), .B(new_n538_), .C1(new_n548_), .C2(new_n549_), .ZN(new_n770_));
  AOI22_X1  g569(.A1(new_n769_), .A2(KEYINPUT55), .B1(new_n560_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT55), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n551_), .A2(new_n558_), .A3(new_n772_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n771_), .A2(new_n773_), .A3(KEYINPUT117), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT117), .B1(new_n771_), .B2(new_n773_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n566_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT56), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT117), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n551_), .A2(new_n772_), .A3(new_n558_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n770_), .A2(new_n560_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n780_), .B1(new_n772_), .B2(new_n550_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n778_), .B1(new_n779_), .B2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n771_), .A2(new_n773_), .A3(KEYINPUT117), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n568_), .A2(new_n777_), .ZN(new_n785_));
  AOI22_X1  g584(.A1(new_n776_), .A2(new_n777_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n484_), .A2(new_n569_), .ZN(new_n787_));
  OAI21_X1  g586(.A(KEYINPUT118), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT118), .ZN(new_n789_));
  INV_X1    g588(.A(new_n787_), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT56), .B1(new_n784_), .B2(new_n566_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n785_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n789_), .B(new_n790_), .C1(new_n791_), .C2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n464_), .A2(new_n466_), .A3(new_n470_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n476_), .B1(new_n469_), .B2(new_n467_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n479_), .A2(new_n797_), .ZN(new_n798_));
  XOR2_X1   g597(.A(new_n798_), .B(KEYINPUT119), .Z(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n570_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n788_), .A2(new_n794_), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n631_), .A2(KEYINPUT57), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n776_), .A2(new_n777_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n792_), .A2(KEYINPUT120), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT120), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n784_), .A2(new_n805_), .A3(new_n785_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n803_), .A2(new_n804_), .A3(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n799_), .A2(new_n569_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n807_), .A2(KEYINPUT58), .A3(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n603_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT58), .B1(new_n807_), .B2(new_n809_), .ZN(new_n812_));
  OAI22_X1  g611(.A1(new_n801_), .A2(new_n802_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n788_), .A2(new_n794_), .A3(new_n800_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT57), .B1(new_n814_), .B2(new_n631_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n620_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n572_), .A2(new_n484_), .A3(new_n574_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n817_), .A2(new_n600_), .A3(new_n619_), .A4(new_n602_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n819_));
  OR3_X1    g618(.A1(new_n818_), .A2(new_n819_), .A3(KEYINPUT54), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(KEYINPUT54), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n818_), .A2(KEYINPUT116), .A3(KEYINPUT54), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n819_), .B1(new_n818_), .B2(KEYINPUT54), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n820_), .A2(new_n823_), .A3(new_n824_), .A4(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n768_), .B1(new_n816_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT59), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n765_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n826_), .ZN(new_n830_));
  AOI22_X1  g629(.A1(KEYINPUT120), .A2(new_n792_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n808_), .B1(new_n831_), .B2(new_n806_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n672_), .B1(new_n832_), .B2(KEYINPUT58), .ZN(new_n833_));
  INV_X1    g632(.A(new_n812_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n802_), .ZN(new_n835_));
  AOI22_X1  g634(.A1(new_n833_), .A2(new_n834_), .B1(new_n814_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT57), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(new_n801_), .B2(new_n733_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n830_), .B1(new_n839_), .B2(new_n620_), .ZN(new_n840_));
  OAI211_X1 g639(.A(KEYINPUT121), .B(KEYINPUT59), .C1(new_n840_), .C2(new_n768_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n829_), .A2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n619_), .B1(new_n836_), .B2(new_n838_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n828_), .B(new_n767_), .C1(new_n843_), .C2(new_n830_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT122), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n816_), .A2(new_n826_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n847_), .A2(KEYINPUT122), .A3(new_n828_), .A4(new_n767_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n842_), .A2(new_n849_), .A3(new_n484_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(G113gat), .ZN(new_n851_));
  INV_X1    g650(.A(new_n827_), .ZN(new_n852_));
  OR2_X1    g651(.A1(new_n483_), .A2(G113gat), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n851_), .B1(new_n852_), .B2(new_n853_), .ZN(G1340gat));
  INV_X1    g653(.A(G120gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n709_), .B2(KEYINPUT60), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n827_), .B(new_n856_), .C1(KEYINPUT60), .C2(new_n855_), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n842_), .A2(new_n577_), .A3(new_n849_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n855_), .ZN(G1341gat));
  NAND2_X1  g658(.A1(new_n619_), .A2(G127gat), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n842_), .A2(new_n849_), .A3(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(G127gat), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(new_n852_), .B2(new_n620_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT123), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n862_), .A2(KEYINPUT123), .A3(new_n864_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1342gat));
  NAND3_X1  g668(.A1(new_n842_), .A2(new_n849_), .A3(new_n603_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(G134gat), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n632_), .A2(G134gat), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n852_), .B2(new_n872_), .ZN(G1343gat));
  INV_X1    g672(.A(KEYINPUT124), .ZN(new_n874_));
  NOR4_X1   g673(.A1(new_n253_), .A2(new_n328_), .A3(new_n440_), .A4(new_n445_), .ZN(new_n875_));
  AND3_X1   g674(.A1(new_n847_), .A2(new_n874_), .A3(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n874_), .B1(new_n847_), .B2(new_n875_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n484_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g678(.A1(new_n876_), .A2(new_n877_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n880_), .A2(new_n709_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(KEYINPUT125), .B(G148gat), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n881_), .B(new_n882_), .ZN(G1345gat));
  NOR2_X1   g682(.A1(new_n880_), .A2(new_n620_), .ZN(new_n884_));
  XOR2_X1   g683(.A(KEYINPUT61), .B(G155gat), .Z(new_n885_));
  XNOR2_X1  g684(.A(new_n884_), .B(new_n885_), .ZN(G1346gat));
  OAI21_X1  g685(.A(G162gat), .B1(new_n880_), .B2(new_n672_), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n632_), .A2(G162gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n880_), .B2(new_n888_), .ZN(G1347gat));
  NOR2_X1   g688(.A1(new_n450_), .A2(new_n441_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n659_), .ZN(new_n892_));
  AND2_X1   g691(.A1(new_n847_), .A2(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n223_), .B1(new_n893_), .B2(new_n484_), .ZN(new_n894_));
  OR2_X1    g693(.A1(new_n894_), .A2(KEYINPUT126), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(KEYINPUT126), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n895_), .A2(KEYINPUT62), .A3(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n894_), .A2(KEYINPUT126), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n893_), .A2(new_n484_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  AOI22_X1  g700(.A1(new_n898_), .A2(new_n899_), .B1(new_n334_), .B2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n897_), .A2(new_n902_), .ZN(G1348gat));
  AOI21_X1  g702(.A(G176gat), .B1(new_n893_), .B2(new_n577_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n840_), .A2(new_n329_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n891_), .A2(new_n224_), .A3(new_n709_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n904_), .B1(new_n905_), .B2(new_n906_), .ZN(G1349gat));
  NAND3_X1  g706(.A1(new_n905_), .A2(new_n619_), .A3(new_n890_), .ZN(new_n908_));
  OR2_X1    g707(.A1(new_n620_), .A2(new_n219_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  AOI22_X1  g709(.A1(new_n908_), .A2(new_n205_), .B1(new_n893_), .B2(new_n910_), .ZN(G1350gat));
  INV_X1    g710(.A(new_n893_), .ZN(new_n912_));
  OAI21_X1  g711(.A(G190gat), .B1(new_n912_), .B2(new_n672_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n632_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n893_), .A2(new_n220_), .A3(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n913_), .A2(new_n915_), .ZN(G1351gat));
  NOR4_X1   g715(.A1(new_n840_), .A2(new_n441_), .A3(new_n253_), .A4(new_n446_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n484_), .ZN(new_n918_));
  INV_X1    g717(.A(G197gat), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n918_), .B1(KEYINPUT127), .B2(new_n919_), .ZN(new_n920_));
  XOR2_X1   g719(.A(KEYINPUT127), .B(G197gat), .Z(new_n921_));
  AOI21_X1  g720(.A(new_n920_), .B1(new_n918_), .B2(new_n921_), .ZN(G1352gat));
  NAND2_X1  g721(.A1(new_n917_), .A2(new_n577_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g723(.A1(new_n917_), .A2(new_n619_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n926_));
  AND2_X1   g725(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n925_), .A2(new_n926_), .A3(new_n927_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n928_), .B1(new_n925_), .B2(new_n926_), .ZN(G1354gat));
  INV_X1    g728(.A(G218gat), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n917_), .A2(new_n930_), .A3(new_n914_), .ZN(new_n931_));
  AND2_X1   g730(.A1(new_n917_), .A2(new_n603_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n932_), .B2(new_n930_), .ZN(G1355gat));
endmodule


