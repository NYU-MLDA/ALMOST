//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 1 0 1 0 1 1 1 1 0 0 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n855_, new_n856_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_;
  INV_X1    g000(.A(KEYINPUT9), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT65), .B(G85gat), .ZN(new_n203_));
  INV_X1    g002(.A(G92gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(new_n202_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT66), .ZN(new_n206_));
  NAND3_X1  g005(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT67), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT67), .B1(G85gat), .B2(G92gat), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n209_), .B1(new_n207_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n206_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G99gat), .A2(G106gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT6), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT10), .B(G99gat), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n212_), .B(new_n214_), .C1(G106gat), .C2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G99gat), .ZN(new_n217_));
  INV_X1    g016(.A(G106gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(new_n218_), .A3(KEYINPUT68), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT68), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n220_), .B1(G99gat), .B2(G106gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT7), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT69), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT69), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT7), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n219_), .A2(new_n221_), .A3(new_n223_), .A4(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(new_n214_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT8), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G85gat), .B(G92gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n229_), .A2(new_n230_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT71), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT6), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT70), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT70), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT6), .ZN(new_n238_));
  AND3_X1   g037(.A1(new_n236_), .A2(new_n238_), .A3(new_n213_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n213_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n234_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n213_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n237_), .A2(KEYINPUT6), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n235_), .A2(KEYINPUT70), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n242_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n236_), .A2(new_n238_), .A3(new_n213_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(KEYINPUT71), .A3(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n228_), .A2(new_n241_), .A3(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n230_), .B1(new_n248_), .B2(new_n232_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n233_), .B1(new_n249_), .B2(KEYINPUT72), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT72), .ZN(new_n251_));
  AOI211_X1 g050(.A(new_n251_), .B(new_n230_), .C1(new_n248_), .C2(new_n232_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n216_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(G71gat), .B(G78gat), .Z(new_n254_));
  XNOR2_X1  g053(.A(G57gat), .B(G64gat), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n254_), .B1(KEYINPUT11), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(KEYINPUT11), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n253_), .B(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT73), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n259_), .B1(new_n260_), .B2(KEYINPUT12), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G230gat), .A2(G233gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT64), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n253_), .A2(new_n258_), .ZN(new_n265_));
  XOR2_X1   g064(.A(KEYINPUT73), .B(KEYINPUT12), .Z(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n261_), .A2(new_n264_), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n259_), .A2(new_n263_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(G120gat), .B(G148gat), .Z(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(G204gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT5), .B(G176gat), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n272_), .B(new_n273_), .Z(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n270_), .A2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n268_), .A2(new_n269_), .A3(new_n274_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT13), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n276_), .A2(KEYINPUT13), .A3(new_n277_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G127gat), .B(G155gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT16), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(G183gat), .ZN(new_n286_));
  INV_X1    g085(.A(G211gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n289_), .A2(KEYINPUT79), .A3(KEYINPUT17), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G15gat), .B(G22gat), .ZN(new_n291_));
  INV_X1    g090(.A(G1gat), .ZN(new_n292_));
  INV_X1    g091(.A(G8gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT14), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n291_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G1gat), .B(G8gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G231gat), .A2(G233gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(new_n258_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n290_), .A2(new_n301_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n290_), .B(new_n301_), .C1(KEYINPUT17), .C2(new_n289_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT80), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT37), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G232gat), .A2(G233gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT34), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT35), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT75), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G29gat), .B(G36gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G43gat), .B(G50gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n216_), .B(new_n316_), .C1(new_n250_), .C2(new_n252_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n310_), .A2(new_n311_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n309_), .A2(KEYINPUT35), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n317_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n316_), .B(KEYINPUT15), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(KEYINPUT71), .B1(new_n245_), .B2(new_n246_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n226_), .A2(new_n227_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n231_), .B1(new_n326_), .B2(new_n247_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n251_), .B1(new_n327_), .B2(new_n230_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n249_), .A2(KEYINPUT72), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n328_), .A2(new_n329_), .A3(new_n233_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n323_), .B1(new_n330_), .B2(new_n216_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n313_), .B1(new_n321_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n253_), .A2(new_n322_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n333_), .A2(new_n312_), .A3(new_n317_), .A4(new_n320_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G190gat), .B(G218gat), .ZN(new_n335_));
  INV_X1    g134(.A(G134gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT74), .ZN(new_n338_));
  INV_X1    g137(.A(G162gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n340_), .B(KEYINPUT36), .Z(new_n341_));
  AND3_X1   g140(.A1(new_n332_), .A2(new_n334_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT77), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n340_), .A2(KEYINPUT36), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n345_), .B1(new_n332_), .B2(new_n334_), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n342_), .A2(new_n343_), .B1(new_n346_), .B2(KEYINPUT76), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n332_), .A2(new_n334_), .A3(new_n341_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT77), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n307_), .B1(new_n347_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n342_), .A2(new_n307_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n332_), .A2(new_n334_), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n352_), .A2(new_n344_), .B1(KEYINPUT76), .B2(KEYINPUT37), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT78), .B1(new_n350_), .B2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n352_), .A2(KEYINPUT76), .A3(new_n344_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n332_), .A2(new_n341_), .A3(new_n334_), .A4(new_n343_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n349_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT37), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT78), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(new_n354_), .A3(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n306_), .B1(new_n356_), .B2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n283_), .A2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT81), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT93), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G226gat), .A2(G233gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT20), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G211gat), .B(G218gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT21), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT21), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n287_), .A2(G218gat), .ZN(new_n376_));
  INV_X1    g175(.A(G218gat), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n377_), .A2(G211gat), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n375_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G197gat), .B(G204gat), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n374_), .A2(new_n379_), .A3(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n373_), .A2(new_n380_), .A3(KEYINPUT21), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G169gat), .A2(G176gat), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT22), .B(G169gat), .ZN(new_n388_));
  INV_X1    g187(.A(G176gat), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n387_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G183gat), .A2(G190gat), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT23), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n393_), .B(new_n394_), .C1(G183gat), .C2(G190gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n390_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT26), .B(G190gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT25), .B(G183gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  AND2_X1   g198(.A1(new_n393_), .A2(new_n394_), .ZN(new_n400_));
  INV_X1    g199(.A(G169gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n389_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(KEYINPUT24), .A3(new_n386_), .ZN(new_n403_));
  OR3_X1    g202(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n399_), .A2(new_n400_), .A3(new_n403_), .A4(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT94), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n404_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n408_), .A2(KEYINPUT94), .A3(new_n403_), .A4(new_n399_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n385_), .A2(new_n396_), .A3(new_n407_), .A4(new_n409_), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n382_), .A2(KEYINPUT87), .A3(new_n383_), .ZN(new_n411_));
  AOI21_X1  g210(.A(KEYINPUT87), .B1(new_n382_), .B2(new_n383_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n400_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT82), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT25), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n415_), .B1(new_n416_), .B2(G183gat), .ZN(new_n417_));
  OAI211_X1 g216(.A(new_n397_), .B(new_n417_), .C1(new_n398_), .C2(new_n415_), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n414_), .A2(new_n418_), .B1(new_n395_), .B2(new_n390_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n413_), .A2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n372_), .A2(new_n410_), .A3(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n407_), .A2(new_n396_), .A3(new_n409_), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT95), .B1(new_n423_), .B2(new_n384_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT87), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n384_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n382_), .A2(KEYINPUT87), .A3(new_n383_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n371_), .B1(new_n429_), .B2(new_n419_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n423_), .A2(KEYINPUT95), .A3(new_n384_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n425_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT96), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n432_), .A2(new_n433_), .A3(new_n370_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n433_), .B1(new_n432_), .B2(new_n370_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n422_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G8gat), .B(G36gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT18), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(G64gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(new_n204_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n436_), .A2(new_n441_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n440_), .B(new_n422_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT100), .B(KEYINPUT27), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT27), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n405_), .A2(new_n396_), .A3(new_n382_), .A4(new_n383_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT20), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n448_), .B1(new_n413_), .B2(new_n420_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT99), .ZN(new_n450_));
  OR3_X1    g249(.A1(new_n449_), .A2(new_n450_), .A3(new_n369_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n450_), .B1(new_n449_), .B2(new_n369_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n425_), .A2(new_n430_), .A3(new_n369_), .A4(new_n431_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n451_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n446_), .B1(new_n454_), .B2(new_n441_), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n444_), .A2(new_n445_), .B1(new_n443_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  XOR2_X1   g256(.A(G155gat), .B(G162gat), .Z(new_n458_));
  OR2_X1    g257(.A1(G141gat), .A2(G148gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT3), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G141gat), .A2(G148gat), .ZN(new_n461_));
  XOR2_X1   g260(.A(new_n461_), .B(KEYINPUT2), .Z(new_n462_));
  OAI21_X1  g261(.A(new_n458_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT1), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n458_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n465_), .A2(new_n459_), .A3(new_n461_), .A4(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n463_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT29), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G228gat), .A2(G233gat), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT86), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n427_), .A2(new_n471_), .A3(new_n428_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT88), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n470_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n470_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n475_), .A2(new_n471_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n413_), .A2(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n469_), .B1(new_n474_), .B2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n384_), .B1(new_n469_), .B2(KEYINPUT88), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(new_n475_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G78gat), .B(G106gat), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT89), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n478_), .A2(new_n480_), .A3(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n483_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n485_));
  OAI22_X1  g284(.A1(new_n484_), .A2(new_n485_), .B1(KEYINPUT89), .B2(new_n482_), .ZN(new_n486_));
  OR2_X1    g285(.A1(new_n468_), .A2(KEYINPUT29), .ZN(new_n487_));
  XOR2_X1   g286(.A(G22gat), .B(G50gat), .Z(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT28), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n487_), .B(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n486_), .A2(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n482_), .A2(KEYINPUT90), .ZN(new_n492_));
  INV_X1    g291(.A(new_n469_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n472_), .A2(new_n473_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(new_n475_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n413_), .A2(new_n476_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n493_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n480_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n492_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n478_), .B(new_n480_), .C1(KEYINPUT90), .C2(new_n482_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n490_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n499_), .A2(new_n500_), .A3(KEYINPUT91), .A4(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT91), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n491_), .A2(new_n502_), .A3(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n419_), .B(KEYINPUT83), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G227gat), .A2(G233gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n508_), .B(KEYINPUT84), .Z(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT30), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n507_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n507_), .A2(new_n510_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G15gat), .B(G43gat), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT85), .ZN(new_n516_));
  XOR2_X1   g315(.A(G127gat), .B(G134gat), .Z(new_n517_));
  XOR2_X1   g316(.A(G113gat), .B(G120gat), .Z(new_n518_));
  XOR2_X1   g317(.A(new_n517_), .B(new_n518_), .Z(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT31), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n516_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n522_), .B1(new_n521_), .B2(new_n520_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G71gat), .B(G99gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n513_), .A2(new_n514_), .ZN(new_n527_));
  OR3_X1    g326(.A1(new_n515_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(G1gat), .B(G29gat), .Z(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT0), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(G57gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(G85gat), .ZN(new_n532_));
  INV_X1    g331(.A(G57gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n530_), .B(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(G85gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n532_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G225gat), .A2(G233gat), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT4), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT97), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n463_), .A2(new_n541_), .A3(new_n467_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n520_), .A2(new_n542_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n519_), .A2(new_n541_), .A3(new_n463_), .A4(new_n467_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n540_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(KEYINPUT98), .B(KEYINPUT4), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n468_), .A2(new_n519_), .A3(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n539_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n543_), .A2(new_n544_), .A3(new_n538_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n537_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n548_), .A2(new_n537_), .A3(new_n549_), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n526_), .B1(new_n527_), .B2(new_n515_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n528_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  NOR3_X1   g354(.A1(new_n457_), .A2(new_n506_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n431_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n419_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(KEYINPUT20), .ZN(new_n559_));
  NOR3_X1   g358(.A1(new_n557_), .A2(new_n559_), .A3(new_n424_), .ZN(new_n560_));
  OAI21_X1  g359(.A(KEYINPUT96), .B1(new_n560_), .B2(new_n369_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n432_), .A2(new_n433_), .A3(new_n370_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n440_), .B1(new_n563_), .B2(new_n422_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n422_), .ZN(new_n565_));
  AOI211_X1 g364(.A(new_n441_), .B(new_n565_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n445_), .B1(new_n564_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n443_), .A2(new_n455_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n506_), .A2(new_n567_), .A3(new_n568_), .A4(new_n553_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT101), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n456_), .A2(KEYINPUT101), .A3(new_n506_), .A4(new_n553_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n440_), .A2(KEYINPUT32), .ZN(new_n573_));
  AOI22_X1  g372(.A1(new_n551_), .A2(new_n552_), .B1(new_n454_), .B2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n574_), .B1(new_n436_), .B2(new_n573_), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n550_), .A2(KEYINPUT33), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n550_), .A2(KEYINPUT33), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n545_), .A2(new_n539_), .A3(new_n547_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n543_), .A2(new_n544_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n537_), .B1(new_n538_), .B2(new_n579_), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n576_), .B(new_n577_), .C1(new_n578_), .C2(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n575_), .B1(new_n444_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n506_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n571_), .A2(new_n572_), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n528_), .A2(new_n554_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n556_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n297_), .B(new_n316_), .Z(new_n588_));
  NAND2_X1  g387(.A1(G229gat), .A2(G233gat), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n322_), .A2(new_n297_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n297_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n590_), .B1(new_n592_), .B2(new_n316_), .ZN(new_n593_));
  AOI22_X1  g392(.A1(new_n588_), .A2(new_n590_), .B1(new_n591_), .B2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G113gat), .B(G141gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(new_n401_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(G197gat), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n594_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n594_), .A2(new_n597_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NOR3_X1   g400(.A1(new_n365_), .A2(new_n587_), .A3(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n553_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n602_), .A2(new_n292_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT38), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(KEYINPUT102), .B1(new_n282_), .B2(new_n601_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n304_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT102), .ZN(new_n609_));
  INV_X1    g408(.A(new_n601_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n280_), .A2(new_n609_), .A3(new_n281_), .A4(new_n610_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n607_), .A2(new_n608_), .A3(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n342_), .A2(new_n346_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n587_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(G1gat), .B1(new_n615_), .B2(new_n553_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n604_), .A2(new_n605_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n606_), .A2(new_n616_), .A3(new_n617_), .ZN(G1324gat));
  NAND3_X1  g417(.A1(new_n602_), .A2(new_n293_), .A3(new_n457_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n612_), .A2(new_n457_), .A3(new_n614_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n620_), .A2(G8gat), .A3(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n621_), .B1(new_n620_), .B2(G8gat), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n619_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g424(.A(G15gat), .B1(new_n615_), .B2(new_n586_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT41), .Z(new_n627_));
  INV_X1    g426(.A(G15gat), .ZN(new_n628_));
  INV_X1    g427(.A(new_n586_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n602_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n627_), .A2(new_n630_), .ZN(G1326gat));
  OAI21_X1  g430(.A(G22gat), .B1(new_n615_), .B2(new_n583_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT42), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n583_), .A2(G22gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT104), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n602_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n633_), .A2(new_n636_), .ZN(G1327gat));
  INV_X1    g436(.A(new_n613_), .ZN(new_n638_));
  NOR4_X1   g437(.A1(new_n282_), .A2(new_n305_), .A3(new_n601_), .A4(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n585_), .A2(new_n586_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n556_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n639_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(G29gat), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(new_n644_), .A3(new_n603_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT105), .ZN(new_n646_));
  AOI221_X4 g445(.A(KEYINPUT78), .B1(new_n351_), .B2(new_n353_), .C1(new_n359_), .C2(KEYINPUT37), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n361_), .B1(new_n360_), .B2(new_n354_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n646_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n356_), .A2(KEYINPUT105), .A3(new_n362_), .ZN(new_n650_));
  AOI22_X1  g449(.A1(new_n569_), .A2(new_n570_), .B1(new_n583_), .B2(new_n582_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n629_), .B1(new_n651_), .B2(new_n572_), .ZN(new_n652_));
  OAI211_X1 g451(.A(new_n649_), .B(new_n650_), .C1(new_n652_), .C2(new_n556_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n356_), .A2(new_n362_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n654_), .A2(KEYINPUT43), .ZN(new_n655_));
  AOI22_X1  g454(.A1(new_n653_), .A2(KEYINPUT43), .B1(new_n642_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT44), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n607_), .A2(new_n306_), .A3(new_n611_), .ZN(new_n658_));
  NOR4_X1   g457(.A1(new_n656_), .A2(KEYINPUT106), .A3(new_n657_), .A4(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT106), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n649_), .A2(new_n650_), .ZN(new_n661_));
  OAI21_X1  g460(.A(KEYINPUT43), .B1(new_n661_), .B2(new_n587_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n642_), .A2(new_n655_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n658_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n660_), .B1(new_n664_), .B2(KEYINPUT44), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n659_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n662_), .A2(new_n663_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n658_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(new_n657_), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n667_), .A2(new_n603_), .A3(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT107), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G29gat), .B1(new_n672_), .B2(new_n673_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n645_), .B1(new_n675_), .B2(new_n676_), .ZN(G1328gat));
  INV_X1    g476(.A(G36gat), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n643_), .A2(new_n678_), .A3(new_n457_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT45), .Z(new_n680_));
  INV_X1    g479(.A(KEYINPUT108), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n457_), .B1(new_n664_), .B2(KEYINPUT44), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n668_), .A2(KEYINPUT44), .A3(new_n669_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT106), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n664_), .A2(new_n660_), .A3(KEYINPUT44), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n682_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n681_), .B1(new_n686_), .B2(new_n678_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n456_), .B1(new_n670_), .B2(new_n657_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n688_), .B1(new_n665_), .B2(new_n659_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(KEYINPUT108), .A3(G36gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n680_), .B1(new_n687_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT46), .ZN(new_n692_));
  AND3_X1   g491(.A1(new_n691_), .A2(KEYINPUT109), .A3(new_n692_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n692_), .A2(KEYINPUT109), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n692_), .A2(KEYINPUT109), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n691_), .A2(new_n694_), .A3(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n693_), .A2(new_n696_), .ZN(G1329gat));
  AOI21_X1  g496(.A(G43gat), .B1(new_n643_), .B2(new_n629_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n671_), .A2(G43gat), .A3(new_n629_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n699_), .B1(new_n666_), .B2(new_n700_), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n701_), .A2(KEYINPUT110), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(KEYINPUT110), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n702_), .A2(new_n703_), .A3(KEYINPUT47), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT47), .B1(new_n702_), .B2(new_n703_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1330gat));
  AOI21_X1  g505(.A(G50gat), .B1(new_n643_), .B2(new_n506_), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n671_), .A2(G50gat), .A3(new_n506_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n667_), .B2(new_n708_), .ZN(G1331gat));
  NOR2_X1   g508(.A1(new_n587_), .A2(new_n610_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT111), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n654_), .A2(new_n305_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n711_), .A2(new_n283_), .A3(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(new_n533_), .A3(new_n603_), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n614_), .A2(new_n282_), .A3(new_n305_), .A4(new_n601_), .ZN(new_n715_));
  OAI21_X1  g514(.A(G57gat), .B1(new_n715_), .B2(new_n553_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1332gat));
  OAI21_X1  g516(.A(G64gat), .B1(new_n715_), .B2(new_n456_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT48), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n456_), .A2(G64gat), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT112), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n713_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n719_), .A2(new_n722_), .ZN(G1333gat));
  OAI21_X1  g522(.A(G71gat), .B1(new_n715_), .B2(new_n586_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT49), .ZN(new_n725_));
  INV_X1    g524(.A(G71gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n713_), .A2(new_n726_), .A3(new_n629_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(new_n728_));
  XOR2_X1   g527(.A(new_n728_), .B(KEYINPUT113), .Z(G1334gat));
  OAI21_X1  g528(.A(G78gat), .B1(new_n715_), .B2(new_n583_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT50), .ZN(new_n731_));
  INV_X1    g530(.A(G78gat), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n713_), .A2(new_n732_), .A3(new_n506_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1335gat));
  NOR4_X1   g533(.A1(new_n711_), .A2(new_n283_), .A3(new_n305_), .A4(new_n638_), .ZN(new_n735_));
  AOI21_X1  g534(.A(G85gat), .B1(new_n735_), .B2(new_n603_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n282_), .A2(new_n306_), .A3(new_n601_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n656_), .A2(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n553_), .A2(new_n203_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n736_), .B1(new_n738_), .B2(new_n739_), .ZN(G1336gat));
  NAND3_X1  g539(.A1(new_n735_), .A2(new_n204_), .A3(new_n457_), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n656_), .A2(new_n456_), .A3(new_n737_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n741_), .B1(new_n204_), .B2(new_n742_), .ZN(G1337gat));
  AOI21_X1  g542(.A(new_n217_), .B1(new_n738_), .B2(new_n629_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n586_), .A2(new_n215_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n735_), .B2(new_n745_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g546(.A1(new_n735_), .A2(new_n218_), .A3(new_n506_), .ZN(new_n748_));
  AOI211_X1 g547(.A(new_n583_), .B(new_n737_), .C1(new_n662_), .C2(new_n663_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT114), .ZN(new_n750_));
  OAI21_X1  g549(.A(G106gat), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n737_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n668_), .A2(new_n506_), .A3(new_n752_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n753_), .A2(KEYINPUT114), .ZN(new_n754_));
  OAI21_X1  g553(.A(KEYINPUT115), .B1(new_n751_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT52), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n218_), .B1(new_n753_), .B2(KEYINPUT114), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT115), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n749_), .A2(new_n750_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n757_), .A2(new_n758_), .A3(new_n759_), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n755_), .A2(new_n756_), .A3(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n756_), .B1(new_n755_), .B2(new_n760_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n748_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT53), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT53), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n765_), .B(new_n748_), .C1(new_n761_), .C2(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1339gat));
  XNOR2_X1  g566(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n768_));
  OR3_X1    g567(.A1(new_n364_), .A2(new_n610_), .A3(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n768_), .B1(new_n364_), .B2(new_n610_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n597_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n589_), .B1(new_n592_), .B2(new_n316_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n591_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n598_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n777_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT119), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n277_), .A2(new_n610_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT117), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n780_), .A2(KEYINPUT117), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n268_), .A2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n261_), .A2(KEYINPUT55), .A3(new_n267_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n264_), .A2(KEYINPUT118), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n786_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n261_), .A2(KEYINPUT55), .A3(new_n267_), .A4(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n784_), .A2(new_n787_), .A3(new_n789_), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n790_), .A2(KEYINPUT56), .A3(new_n275_), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT56), .B1(new_n790_), .B2(new_n275_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n781_), .B(new_n782_), .C1(new_n791_), .C2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n779_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n638_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT57), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n613_), .B1(new_n779_), .B2(new_n793_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT57), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n277_), .A2(new_n776_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n800_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT58), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n654_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  OAI211_X1 g602(.A(KEYINPUT58), .B(new_n800_), .C1(new_n791_), .C2(new_n792_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n797_), .A2(new_n799_), .A3(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n771_), .B1(new_n806_), .B2(new_n304_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n457_), .A2(new_n506_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n808_), .A2(new_n603_), .A3(new_n629_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(G113gat), .B1(new_n810_), .B2(new_n610_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n809_), .A2(KEYINPUT59), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n805_), .B1(KEYINPUT57), .B2(new_n798_), .ZN(new_n813_));
  OR2_X1    g612(.A1(new_n813_), .A2(KEYINPUT121), .ZN(new_n814_));
  INV_X1    g613(.A(new_n799_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n815_), .B1(new_n813_), .B2(KEYINPUT121), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n305_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n812_), .B1(new_n817_), .B2(new_n771_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n304_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n771_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n809_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT120), .B1(new_n823_), .B2(KEYINPUT59), .ZN(new_n824_));
  OAI211_X1 g623(.A(KEYINPUT120), .B(KEYINPUT59), .C1(new_n807_), .C2(new_n809_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n818_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n610_), .A2(G113gat), .ZN(new_n829_));
  XOR2_X1   g628(.A(new_n829_), .B(KEYINPUT122), .Z(new_n830_));
  AOI21_X1  g629(.A(new_n811_), .B1(new_n828_), .B2(new_n830_), .ZN(G1340gat));
  INV_X1    g630(.A(G120gat), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT60), .B1(new_n282_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n283_), .B1(new_n810_), .B2(new_n834_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n818_), .B(new_n835_), .C1(new_n824_), .C2(new_n826_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(G120gat), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n810_), .A2(new_n834_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(KEYINPUT60), .B2(new_n838_), .ZN(G1341gat));
  OAI21_X1  g638(.A(G127gat), .B1(new_n827_), .B2(new_n304_), .ZN(new_n840_));
  OR3_X1    g639(.A1(new_n823_), .A2(G127gat), .A3(new_n306_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(G1342gat));
  OAI21_X1  g641(.A(new_n336_), .B1(new_n823_), .B2(new_n638_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT123), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  OAI211_X1 g644(.A(KEYINPUT123), .B(new_n336_), .C1(new_n823_), .C2(new_n638_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n654_), .A2(new_n336_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n847_), .B1(new_n828_), .B2(new_n848_), .ZN(G1343gat));
  NOR4_X1   g648(.A1(new_n457_), .A2(new_n629_), .A3(new_n583_), .A4(new_n553_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n851_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n610_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n282_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT124), .B(G148gat), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(G1345gat));
  INV_X1    g656(.A(KEYINPUT125), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n858_), .B1(new_n852_), .B2(new_n305_), .ZN(new_n859_));
  NOR4_X1   g658(.A1(new_n807_), .A2(KEYINPUT125), .A3(new_n306_), .A4(new_n851_), .ZN(new_n860_));
  OAI21_X1  g659(.A(KEYINPUT61), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  AOI22_X1  g660(.A1(new_n795_), .A2(new_n796_), .B1(new_n804_), .B2(new_n803_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n608_), .B1(new_n862_), .B2(new_n799_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n305_), .B(new_n850_), .C1(new_n863_), .C2(new_n771_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(KEYINPUT125), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n852_), .A2(new_n858_), .A3(new_n305_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT61), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n865_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n861_), .A2(G155gat), .A3(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(G155gat), .B1(new_n861_), .B2(new_n868_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1346gat));
  AOI21_X1  g670(.A(G162gat), .B1(new_n852_), .B2(new_n613_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n661_), .A2(new_n339_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n872_), .B1(new_n852_), .B2(new_n873_), .ZN(G1347gat));
  INV_X1    g673(.A(KEYINPUT62), .ZN(new_n875_));
  OR2_X1    g674(.A1(new_n456_), .A2(new_n555_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(KEYINPUT126), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(new_n506_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n878_), .B1(new_n817_), .B2(new_n771_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(new_n601_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n875_), .B1(new_n880_), .B2(new_n401_), .ZN(new_n881_));
  OAI211_X1 g680(.A(KEYINPUT62), .B(G169gat), .C1(new_n879_), .C2(new_n601_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n388_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n881_), .A2(new_n882_), .A3(new_n883_), .ZN(G1348gat));
  INV_X1    g683(.A(new_n879_), .ZN(new_n885_));
  AOI21_X1  g684(.A(G176gat), .B1(new_n885_), .B2(new_n282_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n807_), .A2(new_n506_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n877_), .A2(new_n283_), .A3(new_n389_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n886_), .B1(new_n887_), .B2(new_n888_), .ZN(G1349gat));
  NOR3_X1   g688(.A1(new_n879_), .A2(new_n304_), .A3(new_n398_), .ZN(new_n890_));
  INV_X1    g689(.A(G183gat), .ZN(new_n891_));
  INV_X1    g690(.A(new_n877_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n887_), .A2(new_n305_), .A3(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n890_), .B1(new_n891_), .B2(new_n893_), .ZN(G1350gat));
  OAI21_X1  g693(.A(G190gat), .B1(new_n879_), .B2(new_n654_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n613_), .A2(new_n397_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n879_), .B2(new_n896_), .ZN(G1351gat));
  NOR4_X1   g696(.A1(new_n629_), .A2(new_n456_), .A3(new_n583_), .A4(new_n603_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n821_), .A2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n610_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n282_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G204gat), .ZN(G1353gat));
  XOR2_X1   g703(.A(KEYINPUT63), .B(G211gat), .Z(new_n905_));
  NAND3_X1  g704(.A1(new_n900_), .A2(new_n608_), .A3(new_n905_), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n906_), .A2(KEYINPUT127), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n906_), .A2(KEYINPUT127), .ZN(new_n908_));
  AOI211_X1 g707(.A(KEYINPUT63), .B(G211gat), .C1(new_n900_), .C2(new_n608_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n907_), .A2(new_n908_), .A3(new_n909_), .ZN(G1354gat));
  OAI21_X1  g709(.A(G218gat), .B1(new_n899_), .B2(new_n654_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n613_), .A2(new_n377_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n899_), .B2(new_n912_), .ZN(G1355gat));
endmodule


