//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 1 1 1 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 0 1 0 1 0 1 1 1 1 0 0 0 0 0 1 0 0 0 1 0 0 0 1 0 0 1 1 0 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n612_, new_n613_, new_n614_, new_n616_,
    new_n617_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n750_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n804_, new_n806_, new_n807_, new_n808_, new_n809_, new_n811_,
    new_n812_, new_n813_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n823_, new_n824_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(G204gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(G197gat), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n204_), .A2(KEYINPUT93), .ZN(new_n205_));
  OR2_X1    g004(.A1(new_n203_), .A2(G197gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(KEYINPUT93), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G211gat), .B(G218gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT21), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n208_), .A2(new_n211_), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n210_), .B1(new_n206_), .B2(new_n204_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT92), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n209_), .B1(new_n208_), .B2(KEYINPUT21), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n212_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT94), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n218_), .B(KEYINPUT89), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT2), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n222_));
  OR2_X1    g021(.A1(G141gat), .A2(G148gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n223_), .B1(KEYINPUT90), .B2(KEYINPUT3), .ZN(new_n224_));
  OR3_X1    g023(.A1(new_n223_), .A2(KEYINPUT90), .A3(KEYINPUT3), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n221_), .A2(new_n222_), .A3(new_n224_), .A4(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(G155gat), .B(G162gat), .Z(new_n227_));
  INV_X1    g026(.A(KEYINPUT1), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n230_));
  AND3_X1   g029(.A1(new_n219_), .A2(new_n223_), .A3(new_n230_), .ZN(new_n231_));
  AOI22_X1  g030(.A1(new_n226_), .A2(new_n227_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT29), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G228gat), .A2(G233gat), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n235_), .B(KEYINPUT91), .Z(new_n236_));
  NOR2_X1   g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n217_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n216_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n236_), .B1(new_n234_), .B2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  XOR2_X1   g040(.A(G22gat), .B(G50gat), .Z(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n232_), .A2(new_n233_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT28), .ZN(new_n245_));
  XOR2_X1   g044(.A(G78gat), .B(G106gat), .Z(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n243_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n243_), .A2(new_n247_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G127gat), .B(G134gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G113gat), .B(G120gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(new_n232_), .B(new_n254_), .Z(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT4), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G225gat), .A2(G233gat), .ZN(new_n257_));
  OR3_X1    g056(.A1(new_n232_), .A2(KEYINPUT4), .A3(new_n254_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G1gat), .B(G29gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(G85gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT0), .B(G57gat), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n261_), .B(new_n262_), .Z(new_n263_));
  INV_X1    g062(.A(new_n257_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n263_), .B1(new_n255_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n259_), .A2(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT97), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n257_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n255_), .A2(new_n264_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n263_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT33), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n267_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT20), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G183gat), .A2(G190gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT23), .ZN(new_n278_));
  NOR2_X1   g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT24), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(G169gat), .ZN(new_n283_));
  INV_X1    g082(.A(G176gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT24), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n285_), .A2(new_n279_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT86), .B(G190gat), .ZN(new_n287_));
  MUX2_X1   g086(.A(G190gat), .B(new_n287_), .S(KEYINPUT26), .Z(new_n288_));
  INV_X1    g087(.A(G183gat), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n289_), .A2(KEYINPUT85), .ZN(new_n290_));
  XOR2_X1   g089(.A(new_n290_), .B(KEYINPUT25), .Z(new_n291_));
  OAI211_X1 g090(.A(new_n282_), .B(new_n286_), .C1(new_n288_), .C2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n287_), .A2(new_n289_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n278_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(G169gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n292_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT87), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n276_), .B1(new_n300_), .B2(new_n216_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n278_), .B1(G183gat), .B2(G190gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(new_n296_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT95), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n285_), .A2(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n279_), .B1(new_n285_), .B2(new_n304_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT26), .B(G190gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT25), .B(G183gat), .ZN(new_n308_));
  AOI22_X1  g107(.A1(new_n305_), .A2(new_n306_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT96), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n282_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n303_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n301_), .B1(new_n216_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G226gat), .A2(G233gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT19), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n314_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n313_), .A2(new_n216_), .ZN(new_n319_));
  OAI211_X1 g118(.A(KEYINPUT20), .B(new_n319_), .C1(new_n300_), .C2(new_n216_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n318_), .B1(new_n317_), .B2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G8gat), .B(G36gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT18), .ZN(new_n323_));
  XOR2_X1   g122(.A(G64gat), .B(G92gat), .Z(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n321_), .B(new_n325_), .ZN(new_n326_));
  AOI211_X1 g125(.A(new_n275_), .B(new_n326_), .C1(new_n274_), .C2(new_n273_), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n217_), .A2(new_n313_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(new_n301_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n316_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n330_), .B1(new_n316_), .B2(new_n320_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n325_), .A2(KEYINPUT32), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n270_), .A2(new_n271_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n273_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  AOI211_X1 g136(.A(new_n334_), .B(new_n337_), .C1(new_n321_), .C2(new_n333_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n251_), .B1(new_n327_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT98), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  OAI211_X1 g140(.A(KEYINPUT98), .B(new_n251_), .C1(new_n327_), .C2(new_n338_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT27), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n326_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT99), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n343_), .B1(new_n321_), .B2(new_n325_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n346_), .B1(new_n332_), .B2(new_n325_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n337_), .A2(new_n250_), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n341_), .B(new_n342_), .C1(new_n348_), .C2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G227gat), .A2(G233gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(G15gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n300_), .B(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT31), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G71gat), .B(G99gat), .ZN(new_n355_));
  INV_X1    g154(.A(G43gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT88), .B(KEYINPUT30), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n359_), .B(new_n254_), .Z(new_n360_));
  OR2_X1    g159(.A1(new_n354_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n354_), .A2(new_n360_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n350_), .A2(new_n363_), .ZN(new_n364_));
  NOR3_X1   g163(.A1(new_n363_), .A2(new_n250_), .A3(new_n336_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n345_), .A2(new_n347_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT100), .ZN(new_n367_));
  OR2_X1    g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n366_), .A2(new_n367_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n364_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G230gat), .A2(G233gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT64), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT73), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G99gat), .A2(G106gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT6), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT6), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n377_), .A2(G99gat), .A3(G106gat), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n376_), .A2(new_n378_), .A3(KEYINPUT70), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT70), .B1(new_n376_), .B2(new_n378_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(G99gat), .ZN(new_n382_));
  INV_X1    g181(.A(G106gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT68), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT7), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT7), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT68), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n384_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n382_), .A2(new_n383_), .B1(new_n387_), .B2(KEYINPUT68), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT71), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n384_), .A2(new_n388_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT71), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT68), .B(KEYINPUT7), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n392_), .B(new_n393_), .C1(new_n394_), .C2(new_n384_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n381_), .A2(new_n391_), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(G85gat), .ZN(new_n397_));
  INV_X1    g196(.A(G92gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G85gat), .A2(G92gat), .ZN(new_n400_));
  AND2_X1   g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n396_), .A2(KEYINPUT72), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT8), .ZN(new_n403_));
  AOI21_X1  g202(.A(KEYINPUT72), .B1(new_n396_), .B2(new_n401_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n374_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n396_), .A2(new_n401_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT72), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n408_), .A2(KEYINPUT73), .A3(KEYINPUT8), .A4(new_n402_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT8), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n376_), .A2(new_n378_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(KEYINPUT66), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n392_), .B1(new_n394_), .B2(new_n384_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n410_), .B(new_n401_), .C1(new_n412_), .C2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT69), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n405_), .A2(new_n409_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT9), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n399_), .B1(new_n417_), .B2(new_n400_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT65), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n400_), .A2(new_n419_), .A3(new_n417_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n419_), .B1(new_n400_), .B2(new_n417_), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n418_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  XOR2_X1   g221(.A(KEYINPUT10), .B(G99gat), .Z(new_n423_));
  AOI211_X1 g222(.A(new_n422_), .B(new_n412_), .C1(new_n383_), .C2(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT67), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n416_), .A2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G57gat), .B(G64gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT11), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(KEYINPUT74), .ZN(new_n429_));
  XOR2_X1   g228(.A(G71gat), .B(G78gat), .Z(new_n430_));
  OAI21_X1  g229(.A(new_n430_), .B1(KEYINPUT11), .B2(new_n427_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n429_), .B(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n373_), .B1(new_n426_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n426_), .A2(new_n433_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n426_), .A2(KEYINPUT75), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n435_), .A2(new_n436_), .A3(KEYINPUT12), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n432_), .B1(new_n416_), .B2(new_n425_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT75), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n439_), .B1(new_n416_), .B2(new_n425_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT12), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n438_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n434_), .B1(new_n437_), .B2(new_n442_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n416_), .A2(new_n425_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n432_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n373_), .B1(new_n445_), .B2(new_n435_), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT76), .B1(new_n443_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n434_), .ZN(new_n448_));
  NOR3_X1   g247(.A1(new_n438_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n449_));
  AOI221_X4 g248(.A(new_n432_), .B1(new_n439_), .B2(KEYINPUT12), .C1(new_n416_), .C2(new_n425_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n448_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n446_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT76), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n451_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G120gat), .B(G148gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT5), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G176gat), .B(G204gat), .ZN(new_n457_));
  XOR2_X1   g256(.A(new_n456_), .B(new_n457_), .Z(new_n458_));
  NAND3_X1  g257(.A1(new_n447_), .A2(new_n454_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n437_), .A2(new_n442_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n446_), .B1(new_n460_), .B2(new_n448_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n458_), .ZN(new_n462_));
  AOI21_X1  g261(.A(KEYINPUT77), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT77), .ZN(new_n464_));
  NOR4_X1   g263(.A1(new_n443_), .A2(new_n464_), .A3(new_n446_), .A4(new_n458_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n459_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT78), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n451_), .A2(new_n452_), .A3(new_n462_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(new_n464_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n461_), .A2(KEYINPUT77), .A3(new_n462_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n472_), .A2(KEYINPUT78), .A3(new_n459_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n468_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT13), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n468_), .A2(KEYINPUT13), .A3(new_n473_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  XOR2_X1   g277(.A(G29gat), .B(G36gat), .Z(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT80), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G43gat), .B(G50gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT15), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G1gat), .B(G8gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT82), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G15gat), .B(G22gat), .ZN(new_n486_));
  INV_X1    g285(.A(G8gat), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n485_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n485_), .A2(new_n489_), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n483_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n491_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n492_), .B1(new_n482_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G229gat), .A2(G233gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n482_), .B(new_n493_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n497_), .A2(G229gat), .A3(G233gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  XOR2_X1   g298(.A(G113gat), .B(G141gat), .Z(new_n500_));
  XNOR2_X1  g299(.A(G169gat), .B(G197gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n499_), .B(new_n502_), .Z(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n478_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n371_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G231gat), .A2(G233gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n493_), .B(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(new_n432_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(new_n439_), .ZN(new_n510_));
  XOR2_X1   g309(.A(G127gat), .B(G155gat), .Z(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G183gat), .B(G211gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n510_), .A2(KEYINPUT17), .A3(new_n515_), .ZN(new_n516_));
  XOR2_X1   g315(.A(KEYINPUT84), .B(KEYINPUT17), .Z(new_n517_));
  XNOR2_X1  g316(.A(new_n515_), .B(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n509_), .A2(new_n518_), .ZN(new_n519_));
  OR2_X1    g318(.A1(new_n516_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT35), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT79), .B(KEYINPUT34), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G232gat), .A2(G233gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  AOI22_X1  g324(.A1(new_n444_), .A2(new_n482_), .B1(new_n522_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n426_), .A2(new_n483_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT81), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n426_), .A2(KEYINPUT81), .A3(new_n483_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n526_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n525_), .A2(new_n522_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G190gat), .B(G218gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G134gat), .B(G162gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n536_), .A2(KEYINPUT36), .ZN(new_n537_));
  INV_X1    g336(.A(new_n532_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n526_), .A2(new_n529_), .A3(new_n538_), .A4(new_n530_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n533_), .A2(new_n537_), .A3(new_n539_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n533_), .A2(new_n539_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n536_), .B(KEYINPUT36), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n540_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n521_), .A2(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n506_), .A2(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n202_), .B1(new_n545_), .B2(new_n336_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT103), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n543_), .A2(KEYINPUT37), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT37), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n540_), .B(new_n549_), .C1(new_n541_), .C2(new_n542_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(new_n521_), .ZN(new_n553_));
  NOR4_X1   g352(.A1(new_n506_), .A2(G1gat), .A3(new_n553_), .A4(new_n337_), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n554_), .B(KEYINPUT101), .Z(new_n555_));
  AND3_X1   g354(.A1(new_n555_), .A2(KEYINPUT102), .A3(KEYINPUT38), .ZN(new_n556_));
  AOI21_X1  g355(.A(KEYINPUT102), .B1(new_n555_), .B2(KEYINPUT38), .ZN(new_n557_));
  OAI221_X1 g356(.A(new_n547_), .B1(KEYINPUT38), .B2(new_n555_), .C1(new_n556_), .C2(new_n557_), .ZN(G1324gat));
  INV_X1    g357(.A(new_n348_), .ZN(new_n559_));
  NOR3_X1   g358(.A1(new_n506_), .A2(new_n559_), .A3(new_n544_), .ZN(new_n560_));
  OR3_X1    g359(.A1(new_n560_), .A2(KEYINPUT39), .A3(new_n487_), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT39), .B1(new_n560_), .B2(new_n487_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n506_), .A2(new_n553_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n559_), .A2(G8gat), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n561_), .A2(new_n562_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n565_), .B(new_n566_), .Z(G1325gat));
  INV_X1    g366(.A(G15gat), .ZN(new_n568_));
  INV_X1    g367(.A(new_n363_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n568_), .B1(new_n545_), .B2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT41), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n563_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(G1326gat));
  INV_X1    g372(.A(G22gat), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n574_), .B1(new_n545_), .B2(new_n250_), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n575_), .B(KEYINPUT42), .Z(new_n576_));
  NAND3_X1  g375(.A1(new_n563_), .A2(new_n574_), .A3(new_n250_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(G1327gat));
  NOR2_X1   g377(.A1(new_n521_), .A2(new_n543_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n506_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT106), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(G29gat), .B1(new_n583_), .B2(new_n336_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n371_), .A2(KEYINPUT105), .A3(KEYINPUT43), .A4(new_n551_), .ZN(new_n585_));
  OR2_X1    g384(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n586_));
  NAND2_X1  g385(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n587_));
  AOI22_X1  g386(.A1(new_n350_), .A2(new_n363_), .B1(new_n369_), .B2(new_n368_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n586_), .B(new_n587_), .C1(new_n588_), .C2(new_n552_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n585_), .A2(new_n589_), .A3(new_n520_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT44), .ZN(new_n591_));
  INV_X1    g390(.A(new_n505_), .ZN(new_n592_));
  OR3_X1    g391(.A1(new_n590_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n591_), .B1(new_n590_), .B2(new_n592_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n336_), .A2(G29gat), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n584_), .B1(new_n596_), .B2(new_n597_), .ZN(G1328gat));
  NOR2_X1   g397(.A1(new_n559_), .A2(G36gat), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n583_), .A2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n583_), .A2(new_n601_), .A3(new_n599_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(G36gat), .B1(new_n595_), .B2(new_n559_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT46), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n605_), .A2(KEYINPUT46), .A3(new_n606_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(G1329gat));
  AND2_X1   g410(.A1(new_n583_), .A2(new_n569_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n569_), .A2(G43gat), .ZN(new_n613_));
  OAI22_X1  g412(.A1(new_n612_), .A2(G43gat), .B1(new_n595_), .B2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g414(.A(G50gat), .B1(new_n583_), .B2(new_n250_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n250_), .A2(G50gat), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n616_), .B1(new_n596_), .B2(new_n617_), .ZN(G1331gat));
  INV_X1    g417(.A(new_n478_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n619_), .A2(new_n503_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n371_), .A2(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n621_), .A2(new_n553_), .ZN(new_n622_));
  INV_X1    g421(.A(G57gat), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(new_n623_), .A3(new_n336_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n621_), .A2(new_n544_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT108), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n627_), .A2(new_n336_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n624_), .B1(new_n628_), .B2(new_n623_), .ZN(G1332gat));
  INV_X1    g428(.A(G64gat), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n622_), .A2(new_n630_), .A3(new_n348_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT48), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n627_), .A2(new_n348_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n632_), .B1(new_n633_), .B2(G64gat), .ZN(new_n634_));
  AOI211_X1 g433(.A(KEYINPUT48), .B(new_n630_), .C1(new_n627_), .C2(new_n348_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n631_), .B1(new_n634_), .B2(new_n635_), .ZN(G1333gat));
  INV_X1    g435(.A(G71gat), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n622_), .A2(new_n637_), .A3(new_n569_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT49), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n627_), .A2(new_n569_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n639_), .B1(new_n640_), .B2(G71gat), .ZN(new_n641_));
  AOI211_X1 g440(.A(KEYINPUT49), .B(new_n637_), .C1(new_n627_), .C2(new_n569_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n638_), .B1(new_n641_), .B2(new_n642_), .ZN(G1334gat));
  INV_X1    g442(.A(G78gat), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n622_), .A2(new_n644_), .A3(new_n250_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n627_), .A2(new_n250_), .ZN(new_n646_));
  XOR2_X1   g445(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n647_));
  AND3_X1   g446(.A1(new_n646_), .A2(G78gat), .A3(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n647_), .B1(new_n646_), .B2(G78gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n645_), .B1(new_n648_), .B2(new_n649_), .ZN(G1335gat));
  NOR2_X1   g449(.A1(new_n621_), .A2(new_n580_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT110), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(G85gat), .B1(new_n653_), .B2(new_n336_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n585_), .A2(new_n589_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n620_), .A2(new_n520_), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n656_), .A2(KEYINPUT111), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(KEYINPUT111), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n655_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n659_), .B(KEYINPUT112), .Z(new_n660_));
  NOR2_X1   g459(.A1(new_n337_), .A2(new_n397_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n654_), .B1(new_n660_), .B2(new_n661_), .ZN(G1336gat));
  AOI21_X1  g461(.A(G92gat), .B1(new_n653_), .B2(new_n348_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n559_), .A2(new_n398_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n660_), .B2(new_n664_), .ZN(G1337gat));
  AOI21_X1  g464(.A(new_n382_), .B1(new_n659_), .B2(new_n569_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n569_), .A2(new_n423_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n666_), .B1(new_n653_), .B2(new_n667_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g468(.A(KEYINPUT52), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n659_), .A2(new_n250_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n671_), .B2(G106gat), .ZN(new_n672_));
  AOI211_X1 g471(.A(KEYINPUT52), .B(new_n383_), .C1(new_n659_), .C2(new_n250_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n250_), .A2(new_n383_), .ZN(new_n674_));
  OAI22_X1  g473(.A1(new_n672_), .A2(new_n673_), .B1(new_n652_), .B2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT53), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT53), .ZN(new_n677_));
  OAI221_X1 g476(.A(new_n677_), .B1(new_n652_), .B2(new_n674_), .C1(new_n672_), .C2(new_n673_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(G1339gat));
  AOI211_X1 g478(.A(new_n520_), .B(new_n503_), .C1(new_n548_), .C2(new_n550_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n476_), .A2(new_n680_), .A3(new_n477_), .ZN(new_n681_));
  OR2_X1    g480(.A1(KEYINPUT113), .A2(KEYINPUT54), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(KEYINPUT113), .A2(KEYINPUT54), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT114), .Z(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n683_), .A2(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n681_), .A2(new_n682_), .A3(new_n685_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(KEYINPUT55), .B1(new_n443_), .B2(KEYINPUT115), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT115), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT55), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n451_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n445_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n373_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n690_), .A2(new_n693_), .A3(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(new_n458_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT56), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT56), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n697_), .A2(new_n700_), .A3(new_n458_), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n699_), .A2(new_n503_), .A3(new_n472_), .A4(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT116), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  AOI22_X1  g503(.A1(new_n698_), .A2(KEYINPUT56), .B1(new_n470_), .B2(new_n471_), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n705_), .A2(KEYINPUT116), .A3(new_n503_), .A4(new_n701_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n499_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n494_), .A2(G229gat), .A3(G233gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n502_), .B1(new_n497_), .B2(new_n495_), .ZN(new_n709_));
  AOI22_X1  g508(.A1(new_n707_), .A2(new_n502_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n473_), .ZN(new_n711_));
  AOI21_X1  g510(.A(KEYINPUT78), .B1(new_n472_), .B2(new_n459_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n710_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n704_), .A2(new_n706_), .A3(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n543_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT57), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n714_), .A2(KEYINPUT57), .A3(new_n543_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n699_), .A2(new_n472_), .A3(new_n701_), .A4(new_n710_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT58), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n705_), .A2(KEYINPUT58), .A3(new_n701_), .A4(new_n710_), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n721_), .A2(new_n551_), .A3(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n717_), .A2(new_n718_), .A3(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n689_), .B1(new_n725_), .B2(new_n520_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n559_), .A2(new_n569_), .A3(new_n251_), .A4(new_n336_), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT59), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n729_), .B1(new_n726_), .B2(KEYINPUT117), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n728_), .B(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(G113gat), .B1(new_n731_), .B2(new_n504_), .ZN(new_n732_));
  OR3_X1    g531(.A1(new_n728_), .A2(G113gat), .A3(new_n504_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1340gat));
  OAI21_X1  g533(.A(G120gat), .B1(new_n731_), .B2(new_n619_), .ZN(new_n735_));
  INV_X1    g534(.A(G120gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n736_), .B1(new_n619_), .B2(KEYINPUT60), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n737_), .B1(KEYINPUT60), .B2(new_n736_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n735_), .B1(new_n728_), .B2(new_n738_), .ZN(G1341gat));
  OAI21_X1  g538(.A(G127gat), .B1(new_n731_), .B2(new_n520_), .ZN(new_n740_));
  OR3_X1    g539(.A1(new_n728_), .A2(G127gat), .A3(new_n520_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1342gat));
  OAI21_X1  g541(.A(G134gat), .B1(new_n731_), .B2(new_n552_), .ZN(new_n743_));
  OR3_X1    g542(.A1(new_n728_), .A2(G134gat), .A3(new_n543_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1343gat));
  NAND3_X1  g544(.A1(new_n363_), .A2(new_n250_), .A3(new_n336_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n726_), .A2(new_n348_), .A3(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(new_n503_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n478_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g550(.A1(new_n747_), .A2(new_n521_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(KEYINPUT61), .B(G155gat), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n752_), .B(new_n753_), .ZN(G1346gat));
  INV_X1    g553(.A(new_n747_), .ZN(new_n755_));
  OAI21_X1  g554(.A(G162gat), .B1(new_n755_), .B2(new_n552_), .ZN(new_n756_));
  OR2_X1    g555(.A1(new_n543_), .A2(G162gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n756_), .B1(new_n755_), .B2(new_n757_), .ZN(G1347gat));
  AOI21_X1  g557(.A(new_n723_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n521_), .B1(new_n759_), .B2(new_n718_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n348_), .B(new_n365_), .C1(new_n760_), .C2(new_n689_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT118), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n762_), .A2(new_n763_), .A3(new_n503_), .ZN(new_n764_));
  OAI21_X1  g563(.A(KEYINPUT118), .B1(new_n761_), .B2(new_n504_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n764_), .A2(G169gat), .A3(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT62), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT119), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n761_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n689_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n714_), .A2(KEYINPUT57), .A3(new_n543_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT57), .B1(new_n714_), .B2(new_n543_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n771_), .A2(new_n772_), .A3(new_n723_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n770_), .B1(new_n773_), .B2(new_n521_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n774_), .A2(KEYINPUT119), .A3(new_n348_), .A4(new_n365_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n769_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(KEYINPUT22), .B(G169gat), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n503_), .A2(new_n778_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT120), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n767_), .B1(new_n777_), .B2(new_n780_), .ZN(G1348gat));
  NAND3_X1  g580(.A1(new_n762_), .A2(G176gat), .A3(new_n478_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n543_), .ZN(new_n783_));
  AOI22_X1  g582(.A1(new_n703_), .A2(new_n702_), .B1(new_n474_), .B2(new_n710_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n784_), .B2(new_n706_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n724_), .B1(new_n785_), .B2(KEYINPUT57), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n520_), .B1(new_n786_), .B2(new_n771_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n559_), .B1(new_n787_), .B2(new_n770_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT119), .B1(new_n788_), .B2(new_n365_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n365_), .ZN(new_n790_));
  NOR4_X1   g589(.A1(new_n726_), .A2(new_n768_), .A3(new_n559_), .A4(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n478_), .B1(new_n789_), .B2(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT121), .B1(new_n792_), .B2(new_n284_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n619_), .B1(new_n769_), .B2(new_n775_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT121), .ZN(new_n795_));
  NOR3_X1   g594(.A1(new_n794_), .A2(new_n795_), .A3(G176gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n782_), .B1(new_n793_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT122), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT122), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n799_), .B(new_n782_), .C1(new_n793_), .C2(new_n796_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(G1349gat));
  OAI21_X1  g600(.A(new_n289_), .B1(new_n761_), .B2(new_n520_), .ZN(new_n802_));
  OR2_X1    g601(.A1(new_n520_), .A2(new_n308_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n777_), .B2(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT123), .ZN(G1350gat));
  NAND3_X1  g604(.A1(new_n776_), .A2(new_n783_), .A3(new_n307_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n776_), .A2(new_n551_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n807_), .A2(KEYINPUT124), .A3(G190gat), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT124), .B1(new_n807_), .B2(G190gat), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n806_), .B1(new_n808_), .B2(new_n809_), .ZN(G1351gat));
  NAND4_X1  g609(.A1(new_n788_), .A2(new_n363_), .A3(new_n250_), .A4(new_n337_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n811_), .A2(new_n504_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(KEYINPUT125), .B(G197gat), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n812_), .B(new_n813_), .ZN(G1352gat));
  NOR2_X1   g613(.A1(new_n811_), .A2(new_n619_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(new_n203_), .ZN(G1353gat));
  NOR2_X1   g615(.A1(new_n811_), .A2(new_n520_), .ZN(new_n817_));
  XOR2_X1   g616(.A(KEYINPUT63), .B(G211gat), .Z(new_n818_));
  AND3_X1   g617(.A1(new_n817_), .A2(KEYINPUT126), .A3(new_n818_), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n817_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT126), .B1(new_n817_), .B2(new_n818_), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n819_), .A2(new_n820_), .A3(new_n821_), .ZN(G1354gat));
  OAI21_X1  g621(.A(G218gat), .B1(new_n811_), .B2(new_n552_), .ZN(new_n823_));
  OR2_X1    g622(.A1(new_n543_), .A2(G218gat), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n823_), .B1(new_n811_), .B2(new_n824_), .ZN(G1355gat));
endmodule


