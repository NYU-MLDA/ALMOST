//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 0 0 1 0 1 1 0 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 1 1 0 0 0 1 1 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n913_, new_n915_, new_n916_, new_n918_, new_n919_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n944_, new_n945_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n977_, new_n978_, new_n979_;
  OR2_X1    g000(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n202_));
  INV_X1    g001(.A(G106gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n202_), .A2(new_n203_), .A3(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT64), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT64), .ZN(new_n207_));
  NAND4_X1  g006(.A1(new_n202_), .A2(new_n207_), .A3(new_n203_), .A4(new_n204_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  OR2_X1    g008(.A1(G85gat), .A2(G92gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G85gat), .A2(G92gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n210_), .A2(KEYINPUT9), .A3(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G99gat), .A2(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT6), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT6), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(G99gat), .A3(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n211_), .A2(KEYINPUT9), .ZN(new_n218_));
  AND3_X1   g017(.A1(new_n212_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n209_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT66), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n210_), .A2(new_n211_), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n214_), .A2(new_n216_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT7), .ZN(new_n224_));
  INV_X1    g023(.A(G99gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(new_n225_), .A3(new_n203_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n222_), .B1(new_n223_), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT8), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n217_), .A2(new_n227_), .A3(new_n226_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT8), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(new_n232_), .A3(new_n222_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n230_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n209_), .A2(new_n219_), .A3(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n221_), .A2(new_n234_), .A3(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT12), .ZN(new_n238_));
  INV_X1    g037(.A(G64gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(G57gat), .ZN(new_n240_));
  INV_X1    g039(.A(G57gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(G64gat), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n240_), .A2(new_n242_), .A3(KEYINPUT11), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT65), .B(G71gat), .ZN(new_n245_));
  INV_X1    g044(.A(G78gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n245_), .A2(new_n246_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n244_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(KEYINPUT65), .B(G71gat), .Z(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(G78gat), .ZN(new_n252_));
  AOI21_X1  g051(.A(KEYINPUT11), .B1(new_n240_), .B2(new_n242_), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n252_), .B(new_n247_), .C1(new_n253_), .C2(new_n243_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n238_), .B1(new_n250_), .B2(new_n254_), .ZN(new_n255_));
  AOI22_X1  g054(.A1(new_n230_), .A2(new_n233_), .B1(new_n209_), .B2(new_n219_), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n250_), .A2(new_n254_), .ZN(new_n257_));
  AOI22_X1  g056(.A1(new_n237_), .A2(new_n255_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G230gat), .A2(G233gat), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n238_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n258_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n259_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n256_), .A2(new_n257_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n256_), .A2(new_n257_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n262_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(G120gat), .B(G148gat), .Z(new_n267_));
  XNOR2_X1  g066(.A(G176gat), .B(G204gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n261_), .A2(new_n266_), .A3(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n271_), .B1(new_n261_), .B2(new_n266_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(KEYINPUT68), .A2(KEYINPUT13), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  AND2_X1   g076(.A1(KEYINPUT68), .A2(KEYINPUT13), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n275_), .B1(new_n278_), .B2(new_n276_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(G29gat), .B(G36gat), .Z(new_n281_));
  XOR2_X1   g080(.A(G43gat), .B(G50gat), .Z(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G29gat), .B(G36gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G43gat), .B(G50gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n283_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT69), .B(KEYINPUT15), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G15gat), .B(G22gat), .ZN(new_n290_));
  INV_X1    g089(.A(G1gat), .ZN(new_n291_));
  INV_X1    g090(.A(G8gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT14), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n290_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G1gat), .B(G8gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n289_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n287_), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G229gat), .A2(G233gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n297_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n296_), .B(new_n298_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n300_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n301_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G113gat), .B(G141gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G169gat), .B(G197gat), .ZN(new_n307_));
  XOR2_X1   g106(.A(new_n306_), .B(new_n307_), .Z(new_n308_));
  NOR2_X1   g107(.A1(new_n308_), .A2(KEYINPUT75), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n305_), .B(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  AND3_X1   g112(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n314_));
  AOI21_X1  g113(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(G183gat), .ZN(new_n317_));
  INV_X1    g116(.A(G190gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n313_), .B1(new_n316_), .B2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT22), .B(G169gat), .ZN(new_n321_));
  INV_X1    g120(.A(G176gat), .ZN(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT79), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(G169gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT22), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT22), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(G169gat), .ZN(new_n327_));
  AND4_X1   g126(.A1(KEYINPUT79), .A2(new_n325_), .A3(new_n327_), .A4(new_n322_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n320_), .B1(new_n323_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT78), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT24), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n331_), .A2(new_n324_), .A3(new_n322_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n330_), .B1(new_n316_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G183gat), .A2(G190gat), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT23), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n337_));
  AND4_X1   g136(.A1(new_n330_), .A2(new_n332_), .A3(new_n336_), .A4(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n333_), .A2(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(G169gat), .A2(G176gat), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT77), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n341_), .A2(new_n342_), .A3(KEYINPUT24), .A4(new_n312_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n312_), .A2(KEYINPUT24), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT77), .B1(new_n344_), .B2(new_n340_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT26), .B(G190gat), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT76), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n347_), .B1(new_n317_), .B2(KEYINPUT25), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT25), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(G183gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n317_), .A2(KEYINPUT25), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n347_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n343_), .B(new_n345_), .C1(new_n349_), .C2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n329_), .B1(new_n339_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT80), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n329_), .B(KEYINPUT80), .C1(new_n339_), .C2(new_n354_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  XOR2_X1   g158(.A(G71gat), .B(G99gat), .Z(new_n360_));
  XNOR2_X1  g159(.A(G15gat), .B(G43gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n359_), .B(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G127gat), .B(G134gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G113gat), .B(G120gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n363_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n366_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n358_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n318_), .A2(KEYINPUT26), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT26), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(G190gat), .ZN(new_n372_));
  AND3_X1   g171(.A1(new_n348_), .A2(new_n370_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n351_), .A2(new_n352_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT76), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n341_), .A2(KEYINPUT24), .A3(new_n312_), .ZN(new_n376_));
  AOI22_X1  g175(.A1(new_n373_), .A2(new_n375_), .B1(KEYINPUT77), .B2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n332_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT78), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n332_), .A2(new_n336_), .A3(new_n330_), .A4(new_n337_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n377_), .A2(new_n381_), .A3(new_n343_), .ZN(new_n382_));
  AOI21_X1  g181(.A(KEYINPUT80), .B1(new_n382_), .B2(new_n329_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n369_), .A2(new_n383_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n384_), .A2(new_n362_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n362_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n368_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n367_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G227gat), .A2(G233gat), .ZN(new_n389_));
  XOR2_X1   g188(.A(new_n389_), .B(KEYINPUT81), .Z(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT30), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT31), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n388_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n367_), .A2(new_n387_), .A3(new_n392_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT85), .B(G50gat), .ZN(new_n398_));
  NAND3_X1  g197(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT83), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(KEYINPUT83), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(G141gat), .A2(G148gat), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT3), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G141gat), .A2(G148gat), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT2), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n403_), .A2(new_n406_), .A3(new_n409_), .A4(new_n410_), .ZN(new_n411_));
  AND2_X1   g210(.A1(G155gat), .A2(G162gat), .ZN(new_n412_));
  NOR2_X1   g211(.A1(G155gat), .A2(G162gat), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT1), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n413_), .B1(new_n412_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G155gat), .A2(G162gat), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n417_), .A2(KEYINPUT82), .A3(KEYINPUT1), .ZN(new_n418_));
  AOI21_X1  g217(.A(KEYINPUT82), .B1(new_n417_), .B2(KEYINPUT1), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n416_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  XOR2_X1   g219(.A(G141gat), .B(G148gat), .Z(new_n421_));
  AOI22_X1  g220(.A1(new_n411_), .A2(new_n414_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT29), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT84), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n401_), .A2(new_n402_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n406_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n414_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n420_), .A2(new_n421_), .ZN(new_n428_));
  AND4_X1   g227(.A1(KEYINPUT84), .A2(new_n427_), .A3(new_n428_), .A4(new_n423_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n398_), .B1(new_n424_), .B2(new_n429_), .ZN(new_n430_));
  XOR2_X1   g229(.A(KEYINPUT28), .B(G22gat), .Z(new_n431_));
  NAND3_X1  g230(.A1(new_n427_), .A2(new_n428_), .A3(new_n423_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT84), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n422_), .A2(KEYINPUT84), .A3(new_n423_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n398_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n434_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n430_), .A2(new_n431_), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G228gat), .A2(G233gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n427_), .A2(new_n428_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT29), .ZN(new_n441_));
  OR2_X1    g240(.A1(G197gat), .A2(G204gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G197gat), .A2(G204gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(KEYINPUT21), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT21), .ZN(new_n445_));
  AND2_X1   g244(.A1(G197gat), .A2(G204gat), .ZN(new_n446_));
  NOR2_X1   g245(.A1(G197gat), .A2(G204gat), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n445_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT87), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G211gat), .B(G218gat), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n444_), .A2(new_n448_), .A3(new_n449_), .A4(new_n450_), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n444_), .A2(new_n448_), .A3(new_n450_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT87), .B1(new_n444_), .B2(new_n450_), .ZN(new_n453_));
  OAI211_X1 g252(.A(KEYINPUT86), .B(new_n451_), .C1(new_n452_), .C2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n439_), .B1(new_n441_), .B2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n423_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n439_), .ZN(new_n458_));
  NOR3_X1   g257(.A1(new_n457_), .A2(new_n454_), .A3(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT88), .B1(new_n456_), .B2(new_n459_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n438_), .A2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n431_), .B1(new_n430_), .B2(new_n437_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n441_), .A2(new_n455_), .A3(new_n439_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n458_), .B1(new_n457_), .B2(new_n454_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT88), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n464_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  XOR2_X1   g266(.A(G78gat), .B(G106gat), .Z(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n468_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n464_), .A2(new_n465_), .A3(new_n466_), .A4(new_n470_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n461_), .A2(new_n463_), .A3(new_n469_), .A4(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n469_), .A2(new_n471_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n438_), .A2(new_n460_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n473_), .B1(new_n474_), .B2(new_n462_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n472_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT27), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G8gat), .B(G36gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT18), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G64gat), .B(G92gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n451_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n357_), .A2(new_n358_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT20), .ZN(new_n485_));
  INV_X1    g284(.A(new_n483_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n374_), .A2(KEYINPUT89), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT89), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n351_), .A2(new_n352_), .A3(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n346_), .A3(new_n489_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n344_), .A2(new_n340_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n378_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n321_), .A2(new_n322_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n320_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n485_), .B1(new_n486_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n484_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G226gat), .A2(G233gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT19), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n486_), .B1(new_n369_), .B2(new_n383_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n500_), .ZN(new_n503_));
  OAI211_X1 g302(.A(KEYINPUT20), .B(new_n503_), .C1(new_n486_), .C2(new_n496_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n482_), .B1(new_n501_), .B2(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n503_), .B1(new_n484_), .B2(new_n497_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n504_), .B1(new_n359_), .B2(new_n486_), .ZN(new_n509_));
  NOR3_X1   g308(.A1(new_n508_), .A2(new_n509_), .A3(new_n481_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n477_), .B1(new_n507_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n440_), .A2(new_n368_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n422_), .A2(new_n366_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G225gat), .A2(G233gat), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n514_), .B(KEYINPUT90), .Z(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n512_), .A2(new_n513_), .A3(new_n516_), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n512_), .A2(new_n513_), .A3(KEYINPUT4), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT4), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n440_), .A2(new_n519_), .A3(new_n368_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(new_n515_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n517_), .B1(new_n518_), .B2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G1gat), .B(G29gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(G85gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT0), .B(G57gat), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n524_), .B(new_n525_), .Z(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n522_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT95), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n517_), .B(new_n526_), .C1(new_n518_), .C2(new_n521_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n522_), .A2(KEYINPUT95), .A3(new_n527_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n476_), .A2(new_n511_), .A3(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT92), .B(KEYINPUT20), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  AOI22_X1  g335(.A1(new_n490_), .A2(new_n492_), .B1(new_n320_), .B2(new_n494_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n483_), .B1(new_n537_), .B2(KEYINPUT93), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n493_), .A2(KEYINPUT93), .A3(new_n495_), .ZN(new_n539_));
  OAI211_X1 g338(.A(KEYINPUT94), .B(new_n536_), .C1(new_n538_), .C2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n502_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT93), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n496_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n537_), .A2(KEYINPUT93), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(new_n483_), .A3(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(KEYINPUT94), .B1(new_n545_), .B2(new_n536_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n500_), .B1(new_n541_), .B2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n484_), .A2(new_n503_), .A3(new_n497_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n482_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n501_), .A2(new_n482_), .A3(new_n506_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT27), .ZN(new_n551_));
  OAI21_X1  g350(.A(KEYINPUT96), .B1(new_n549_), .B2(new_n551_), .ZN(new_n552_));
  AOI22_X1  g351(.A1(new_n498_), .A2(new_n500_), .B1(new_n502_), .B2(new_n505_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n477_), .B1(new_n553_), .B2(new_n482_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT96), .ZN(new_n555_));
  INV_X1    g354(.A(new_n548_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n536_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT94), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n559_), .A2(new_n502_), .A3(new_n540_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n556_), .B1(new_n560_), .B2(new_n500_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n554_), .B(new_n555_), .C1(new_n561_), .C2(new_n482_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n534_), .B1(new_n552_), .B2(new_n562_), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n531_), .A2(new_n532_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n547_), .A2(new_n548_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n482_), .A2(KEYINPUT32), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n553_), .A2(new_n566_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n564_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT33), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n520_), .A2(new_n516_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n512_), .A2(new_n513_), .A3(KEYINPUT4), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n526_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n512_), .A2(new_n513_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT91), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n512_), .A2(new_n513_), .A3(KEYINPUT91), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n577_), .A2(new_n515_), .A3(new_n578_), .ZN(new_n579_));
  AOI22_X1  g378(.A1(new_n571_), .A2(new_n530_), .B1(new_n574_), .B2(new_n579_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n530_), .A2(new_n571_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n481_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n580_), .A2(new_n581_), .A3(new_n550_), .A4(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n476_), .B1(new_n570_), .B2(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n397_), .B1(new_n563_), .B2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n552_), .A2(new_n562_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n564_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n476_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n586_), .A2(new_n587_), .A3(new_n588_), .A4(new_n511_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n311_), .B1(new_n585_), .B2(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(G127gat), .B(G155gat), .Z(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT16), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G183gat), .B(G211gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT17), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n594_), .A2(new_n595_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G231gat), .A2(G233gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n296_), .B(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(new_n257_), .ZN(new_n600_));
  AOI211_X1 g399(.A(new_n596_), .B(new_n597_), .C1(new_n600_), .C2(KEYINPUT74), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n601_), .B1(KEYINPUT74), .B2(new_n600_), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n596_), .B(KEYINPUT73), .Z(new_n603_));
  OR2_X1    g402(.A1(new_n603_), .A2(new_n600_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT37), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n237_), .A2(new_n289_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT35), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G232gat), .A2(G233gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT34), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  AOI22_X1  g411(.A1(new_n256_), .A2(new_n287_), .B1(new_n609_), .B2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n608_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n233_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n232_), .B1(new_n231_), .B2(new_n222_), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n220_), .B(new_n287_), .C1(new_n615_), .C2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT70), .ZN(new_n618_));
  AOI211_X1 g417(.A(new_n609_), .B(new_n612_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n614_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n611_), .A2(KEYINPUT35), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n608_), .B(new_n613_), .C1(new_n618_), .C2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G190gat), .B(G218gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G134gat), .B(G162gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT36), .Z(new_n627_));
  AOI21_X1  g426(.A(new_n607_), .B1(new_n623_), .B2(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n626_), .A2(KEYINPUT36), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n620_), .A2(new_n622_), .A3(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT71), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT71), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n620_), .A2(new_n632_), .A3(new_n622_), .A4(new_n629_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n628_), .A2(new_n631_), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n630_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n627_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n636_), .B1(new_n623_), .B2(KEYINPUT72), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT72), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n620_), .A2(new_n638_), .A3(new_n622_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n635_), .B1(new_n637_), .B2(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n634_), .B1(new_n640_), .B2(KEYINPUT37), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  AND4_X1   g441(.A1(new_n280_), .A2(new_n590_), .A3(new_n606_), .A4(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n643_), .A2(new_n291_), .A3(new_n564_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n640_), .B1(new_n585_), .B2(new_n589_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n280_), .A2(KEYINPUT97), .A3(new_n310_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT97), .B1(new_n280_), .B2(new_n310_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n645_), .A2(new_n649_), .A3(new_n606_), .ZN(new_n650_));
  OAI21_X1  g449(.A(G1gat), .B1(new_n650_), .B2(new_n533_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n644_), .A2(new_n651_), .ZN(new_n652_));
  MUX2_X1   g451(.A(new_n644_), .B(new_n652_), .S(KEYINPUT38), .Z(G1324gat));
  NAND2_X1  g452(.A1(new_n586_), .A2(new_n511_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n643_), .A2(new_n292_), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n654_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G8gat), .B1(new_n650_), .B2(new_n656_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n657_), .A2(KEYINPUT39), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(KEYINPUT39), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n655_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT40), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n660_), .B(new_n661_), .ZN(G1325gat));
  OAI21_X1  g461(.A(G15gat), .B1(new_n650_), .B2(new_n397_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT41), .Z(new_n664_));
  INV_X1    g463(.A(G15gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n643_), .A2(new_n665_), .A3(new_n396_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(G1326gat));
  OAI21_X1  g466(.A(G22gat), .B1(new_n650_), .B2(new_n588_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT42), .ZN(new_n669_));
  INV_X1    g468(.A(G22gat), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n643_), .A2(new_n670_), .A3(new_n476_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(G1327gat));
  INV_X1    g471(.A(new_n280_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n605_), .A2(new_n640_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n590_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(G29gat), .B1(new_n677_), .B2(new_n564_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n648_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n679_), .A2(new_n646_), .A3(new_n605_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n641_), .B2(KEYINPUT98), .ZN(new_n683_));
  AOI211_X1 g482(.A(new_n642_), .B(new_n683_), .C1(new_n585_), .C2(new_n589_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n683_), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n476_), .A2(new_n533_), .A3(new_n511_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n561_), .A2(new_n566_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n569_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n583_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  AOI22_X1  g488(.A1(new_n686_), .A2(new_n586_), .B1(new_n689_), .B2(new_n588_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n589_), .B1(new_n690_), .B2(new_n396_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n685_), .B1(new_n691_), .B2(new_n641_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n681_), .B1(new_n684_), .B2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT99), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT99), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n696_), .B(new_n681_), .C1(new_n684_), .C2(new_n692_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n694_), .A2(new_n695_), .A3(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n686_), .A2(new_n586_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n689_), .A2(new_n588_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n396_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n589_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n641_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(new_n683_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n691_), .A2(new_n641_), .A3(new_n685_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n680_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT44), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n698_), .A2(new_n707_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n564_), .A2(G29gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n678_), .B1(new_n708_), .B2(new_n709_), .ZN(G1328gat));
  INV_X1    g509(.A(KEYINPUT46), .ZN(new_n711_));
  INV_X1    g510(.A(G36gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n656_), .B1(new_n706_), .B2(KEYINPUT44), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n698_), .B2(new_n713_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n656_), .A2(KEYINPUT100), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n656_), .A2(KEYINPUT100), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(new_n712_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(KEYINPUT101), .B(KEYINPUT45), .ZN(new_n719_));
  OR3_X1    g518(.A1(new_n718_), .A2(new_n676_), .A3(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n718_), .B2(new_n676_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n711_), .B1(new_n714_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n722_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n654_), .B1(new_n693_), .B2(new_n695_), .ZN(new_n725_));
  AOI21_X1  g524(.A(KEYINPUT44), .B1(new_n693_), .B2(KEYINPUT99), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n697_), .B2(new_n726_), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n724_), .B(KEYINPUT46), .C1(new_n727_), .C2(new_n712_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n723_), .A2(new_n728_), .ZN(G1329gat));
  INV_X1    g528(.A(G43gat), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n397_), .A2(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n695_), .B1(new_n706_), .B2(new_n696_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n697_), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n707_), .B(new_n731_), .C1(new_n732_), .C2(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n730_), .B1(new_n676_), .B2(new_n397_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT47), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT47), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n734_), .A2(new_n738_), .A3(new_n735_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(G1330gat));
  INV_X1    g539(.A(G50gat), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n588_), .A2(new_n741_), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n707_), .B(new_n742_), .C1(new_n732_), .C2(new_n733_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n741_), .B1(new_n676_), .B2(new_n588_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT102), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n743_), .A2(KEYINPUT102), .A3(new_n744_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1331gat));
  NOR2_X1   g548(.A1(new_n605_), .A2(new_n310_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n645_), .A2(new_n673_), .A3(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n751_), .A2(G57gat), .A3(new_n564_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n752_), .A2(KEYINPUT103), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n752_), .A2(KEYINPUT103), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n310_), .B1(new_n585_), .B2(new_n589_), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n280_), .A2(new_n641_), .A3(new_n605_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(G57gat), .B1(new_n757_), .B2(new_n564_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n753_), .A2(new_n754_), .A3(new_n758_), .ZN(G1332gat));
  AOI21_X1  g558(.A(new_n239_), .B1(new_n751_), .B2(new_n717_), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT48), .Z(new_n761_));
  NAND3_X1  g560(.A1(new_n757_), .A2(new_n239_), .A3(new_n717_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(G1333gat));
  INV_X1    g562(.A(G71gat), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n757_), .A2(new_n764_), .A3(new_n396_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT49), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n751_), .A2(new_n396_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n767_), .B2(G71gat), .ZN(new_n768_));
  AOI211_X1 g567(.A(KEYINPUT49), .B(new_n764_), .C1(new_n751_), .C2(new_n396_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n765_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT104), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n770_), .B(new_n771_), .ZN(G1334gat));
  AOI21_X1  g571(.A(new_n246_), .B1(new_n751_), .B2(new_n476_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(KEYINPUT105), .B(KEYINPUT50), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n773_), .B(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n757_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n476_), .A2(new_n246_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT106), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n775_), .B1(new_n776_), .B2(new_n778_), .ZN(G1335gat));
  NOR2_X1   g578(.A1(new_n684_), .A2(new_n692_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n673_), .A2(new_n311_), .A3(new_n605_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT107), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(G85gat), .B1(new_n784_), .B2(new_n533_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n280_), .A2(new_n674_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n755_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(G85gat), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n788_), .A3(new_n564_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n785_), .A2(new_n789_), .ZN(G1336gat));
  AOI21_X1  g589(.A(G92gat), .B1(new_n787_), .B2(new_n654_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n717_), .A2(G92gat), .ZN(new_n792_));
  XOR2_X1   g591(.A(new_n792_), .B(KEYINPUT108), .Z(new_n793_));
  INV_X1    g592(.A(new_n784_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n791_), .B1(new_n793_), .B2(new_n794_), .ZN(G1337gat));
  INV_X1    g594(.A(KEYINPUT110), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n796_), .A2(KEYINPUT51), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n396_), .A2(new_n202_), .A3(new_n204_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n755_), .A2(new_n786_), .A3(new_n798_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT109), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n783_), .B(new_n396_), .C1(new_n684_), .C2(new_n692_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(G99gat), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n797_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n796_), .A2(KEYINPUT51), .ZN(new_n804_));
  XOR2_X1   g603(.A(new_n804_), .B(KEYINPUT111), .Z(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n803_), .B(new_n806_), .ZN(G1338gat));
  OAI211_X1 g606(.A(new_n783_), .B(new_n476_), .C1(new_n684_), .C2(new_n692_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(G106gat), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n755_), .A2(new_n203_), .A3(new_n476_), .A4(new_n786_), .ZN(new_n812_));
  XOR2_X1   g611(.A(new_n812_), .B(KEYINPUT112), .Z(new_n813_));
  NAND3_X1  g612(.A1(new_n808_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n811_), .A2(new_n813_), .A3(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT53), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n811_), .A2(new_n813_), .A3(new_n817_), .A4(new_n814_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(G1339gat));
  NAND3_X1  g618(.A1(new_n297_), .A2(new_n299_), .A3(new_n303_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n308_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n302_), .A2(new_n300_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n820_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n823_), .A2(new_n824_), .ZN(new_n826_));
  OAI22_X1  g625(.A1(new_n825_), .A2(new_n826_), .B1(new_n821_), .B2(new_n305_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n827_), .A2(new_n273_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n259_), .B1(new_n258_), .B2(new_n260_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n261_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n258_), .A2(KEYINPUT55), .A3(new_n259_), .A4(new_n260_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n271_), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT56), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT56), .ZN(new_n836_));
  AOI211_X1 g635(.A(new_n836_), .B(new_n271_), .C1(new_n831_), .C2(new_n832_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n828_), .B1(new_n835_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT58), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n828_), .B(KEYINPUT58), .C1(new_n835_), .C2(new_n837_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n641_), .A3(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n637_), .A2(new_n639_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n630_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n275_), .A2(new_n827_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n310_), .A2(new_n272_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n236_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n235_), .B1(new_n209_), .B2(new_n219_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n255_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n850_), .A2(new_n260_), .A3(new_n263_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n830_), .B1(new_n851_), .B2(new_n262_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n851_), .A2(new_n262_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n832_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n834_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n836_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n833_), .A2(KEYINPUT56), .A3(new_n834_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n847_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n846_), .B1(new_n859_), .B2(KEYINPUT114), .ZN(new_n860_));
  INV_X1    g659(.A(new_n847_), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n861_), .B(KEYINPUT114), .C1(new_n835_), .C2(new_n837_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n844_), .B1(new_n860_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT57), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n842_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n861_), .B1(new_n835_), .B2(new_n837_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT114), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n845_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n640_), .B1(new_n869_), .B2(new_n862_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n870_), .A2(KEYINPUT57), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n605_), .B1(new_n866_), .B2(new_n871_), .ZN(new_n872_));
  AND3_X1   g671(.A1(new_n280_), .A2(new_n750_), .A3(KEYINPUT113), .ZN(new_n873_));
  AOI21_X1  g672(.A(KEYINPUT113), .B1(new_n280_), .B2(new_n750_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n642_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(KEYINPUT54), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n872_), .A2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n656_), .A2(new_n564_), .A3(new_n588_), .A4(new_n396_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n877_), .A2(new_n878_), .A3(new_n880_), .ZN(new_n881_));
  AND3_X1   g680(.A1(new_n840_), .A2(new_n641_), .A3(new_n841_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n882_), .B1(new_n870_), .B2(KEYINPUT57), .ZN(new_n883_));
  OAI21_X1  g682(.A(KEYINPUT116), .B1(new_n870_), .B2(KEYINPUT57), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT116), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n864_), .A2(new_n885_), .A3(new_n865_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n883_), .A2(new_n884_), .A3(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n605_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n879_), .B1(new_n888_), .B2(new_n876_), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n881_), .B(new_n310_), .C1(new_n889_), .C2(new_n878_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(G113gat), .ZN(new_n891_));
  INV_X1    g690(.A(G113gat), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n889_), .A2(new_n892_), .A3(new_n310_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n893_), .ZN(G1340gat));
  OAI211_X1 g693(.A(new_n881_), .B(new_n673_), .C1(new_n889_), .C2(new_n878_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(G120gat), .ZN(new_n896_));
  INV_X1    g695(.A(G120gat), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n897_), .B1(new_n280_), .B2(KEYINPUT60), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n889_), .B(new_n898_), .C1(KEYINPUT60), .C2(new_n897_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n896_), .A2(new_n899_), .ZN(G1341gat));
  OAI211_X1 g699(.A(new_n881_), .B(new_n606_), .C1(new_n889_), .C2(new_n878_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(G127gat), .ZN(new_n902_));
  INV_X1    g701(.A(G127gat), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n889_), .A2(new_n903_), .A3(new_n606_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n904_), .ZN(G1342gat));
  OAI211_X1 g704(.A(new_n881_), .B(new_n641_), .C1(new_n889_), .C2(new_n878_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(G134gat), .ZN(new_n907_));
  INV_X1    g706(.A(G134gat), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n889_), .A2(new_n908_), .A3(new_n640_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n907_), .A2(new_n909_), .ZN(G1343gat));
  NAND2_X1  g709(.A1(new_n888_), .A2(new_n876_), .ZN(new_n911_));
  NOR4_X1   g710(.A1(new_n717_), .A2(new_n533_), .A3(new_n588_), .A4(new_n396_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n911_), .A2(new_n310_), .A3(new_n912_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g713(.A1(new_n911_), .A2(new_n673_), .A3(new_n912_), .ZN(new_n915_));
  XOR2_X1   g714(.A(KEYINPUT117), .B(G148gat), .Z(new_n916_));
  XNOR2_X1  g715(.A(new_n915_), .B(new_n916_), .ZN(G1345gat));
  NAND3_X1  g716(.A1(new_n911_), .A2(new_n606_), .A3(new_n912_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(KEYINPUT61), .B(G155gat), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n918_), .B(new_n919_), .ZN(G1346gat));
  AND2_X1   g719(.A1(new_n911_), .A2(new_n912_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(new_n640_), .ZN(new_n922_));
  INV_X1    g721(.A(G162gat), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n641_), .A2(G162gat), .ZN(new_n924_));
  XOR2_X1   g723(.A(new_n924_), .B(KEYINPUT118), .Z(new_n925_));
  AOI22_X1  g724(.A1(new_n922_), .A2(new_n923_), .B1(new_n921_), .B2(new_n925_), .ZN(G1347gat));
  AOI21_X1  g725(.A(new_n476_), .B1(new_n872_), .B2(new_n876_), .ZN(new_n927_));
  AND2_X1   g726(.A1(new_n717_), .A2(new_n587_), .ZN(new_n928_));
  AND2_X1   g727(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n310_), .A2(new_n321_), .ZN(new_n930_));
  XOR2_X1   g729(.A(new_n930_), .B(KEYINPUT121), .Z(new_n931_));
  NAND2_X1  g730(.A1(new_n929_), .A2(new_n931_), .ZN(new_n932_));
  OAI211_X1 g731(.A(new_n587_), .B(new_n310_), .C1(new_n715_), .C2(new_n716_), .ZN(new_n933_));
  XOR2_X1   g732(.A(new_n933_), .B(KEYINPUT119), .Z(new_n934_));
  AOI21_X1  g733(.A(new_n324_), .B1(new_n927_), .B2(new_n934_), .ZN(new_n935_));
  AND2_X1   g734(.A1(KEYINPUT120), .A2(KEYINPUT62), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(KEYINPUT120), .B(KEYINPUT62), .ZN(new_n938_));
  OAI211_X1 g737(.A(new_n932_), .B(new_n937_), .C1(new_n935_), .C2(new_n938_), .ZN(G1348gat));
  NAND3_X1  g738(.A1(new_n928_), .A2(G176gat), .A3(new_n673_), .ZN(new_n940_));
  AOI211_X1 g739(.A(new_n476_), .B(new_n940_), .C1(new_n876_), .C2(new_n888_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n929_), .A2(new_n673_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n941_), .B1(new_n942_), .B2(new_n322_), .ZN(G1349gat));
  NAND4_X1  g742(.A1(new_n911_), .A2(new_n588_), .A3(new_n606_), .A4(new_n928_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n605_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n945_));
  AOI22_X1  g744(.A1(new_n317_), .A2(new_n944_), .B1(new_n929_), .B2(new_n945_), .ZN(G1350gat));
  NAND2_X1  g745(.A1(new_n927_), .A2(new_n928_), .ZN(new_n947_));
  OAI21_X1  g746(.A(G190gat), .B1(new_n947_), .B2(new_n642_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n640_), .A2(new_n346_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n949_), .B(KEYINPUT122), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n948_), .B1(new_n947_), .B2(new_n950_), .ZN(G1351gat));
  NAND3_X1  g750(.A1(new_n397_), .A2(new_n533_), .A3(new_n476_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n952_), .B(KEYINPUT123), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n717_), .A2(new_n953_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n954_), .B1(new_n888_), .B2(new_n876_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(KEYINPUT124), .A2(G197gat), .ZN(new_n956_));
  OR2_X1    g755(.A1(KEYINPUT124), .A2(G197gat), .ZN(new_n957_));
  AOI22_X1  g756(.A1(new_n955_), .A2(new_n310_), .B1(new_n956_), .B2(new_n957_), .ZN(new_n958_));
  INV_X1    g757(.A(new_n955_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(new_n959_), .A2(new_n311_), .ZN(new_n960_));
  AOI21_X1  g759(.A(new_n958_), .B1(new_n960_), .B2(new_n957_), .ZN(G1352gat));
  INV_X1    g760(.A(KEYINPUT125), .ZN(new_n962_));
  AND2_X1   g761(.A1(new_n962_), .A2(G204gat), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n962_), .A2(G204gat), .ZN(new_n964_));
  OAI211_X1 g763(.A(new_n955_), .B(new_n673_), .C1(new_n963_), .C2(new_n964_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n959_), .A2(new_n280_), .ZN(new_n966_));
  OAI21_X1  g765(.A(new_n965_), .B1(new_n966_), .B2(new_n964_), .ZN(G1353gat));
  AOI21_X1  g766(.A(new_n605_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n968_));
  NOR2_X1   g767(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n969_), .B(KEYINPUT126), .ZN(new_n970_));
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n971_));
  OR2_X1    g770(.A1(new_n970_), .A2(new_n971_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n970_), .A2(new_n971_), .ZN(new_n973_));
  AOI22_X1  g772(.A1(new_n955_), .A2(new_n968_), .B1(new_n972_), .B2(new_n973_), .ZN(new_n974_));
  AND2_X1   g773(.A1(new_n955_), .A2(new_n968_), .ZN(new_n975_));
  AOI21_X1  g774(.A(new_n974_), .B1(new_n975_), .B2(new_n973_), .ZN(G1354gat));
  OAI21_X1  g775(.A(G218gat), .B1(new_n959_), .B2(new_n642_), .ZN(new_n977_));
  INV_X1    g776(.A(G218gat), .ZN(new_n978_));
  NAND3_X1  g777(.A1(new_n955_), .A2(new_n978_), .A3(new_n640_), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n977_), .A2(new_n979_), .ZN(G1355gat));
endmodule


