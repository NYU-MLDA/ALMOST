//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 1 1 1 0 0 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1 1 1 0 0 0 0 1 0 0 0 0 0 1 0 0 1 1 0 1 1 1 0 1 0 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n818_, new_n819_, new_n820_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n930_,
    new_n931_, new_n932_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n978_, new_n979_, new_n981_, new_n982_, new_n984_, new_n985_,
    new_n987_, new_n989_, new_n990_, new_n991_, new_n993_, new_n994_,
    new_n995_;
  OAI21_X1  g000(.A(KEYINPUT86), .B1(G155gat), .B2(G162gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NOR3_X1   g002(.A1(KEYINPUT86), .A2(G155gat), .A3(G162gat), .ZN(new_n204_));
  AND3_X1   g003(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n205_));
  AOI21_X1  g004(.A(KEYINPUT1), .B1(G155gat), .B2(G162gat), .ZN(new_n206_));
  OAI22_X1  g005(.A1(new_n203_), .A2(new_n204_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(G141gat), .B(G148gat), .Z(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n210_));
  INV_X1    g009(.A(G141gat), .ZN(new_n211_));
  INV_X1    g010(.A(G148gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n213_), .A2(new_n216_), .A3(new_n217_), .A4(new_n218_), .ZN(new_n219_));
  AND2_X1   g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT86), .ZN(new_n221_));
  INV_X1    g020(.A(G155gat), .ZN(new_n222_));
  INV_X1    g021(.A(G162gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n220_), .B1(new_n224_), .B2(new_n202_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n219_), .A2(new_n225_), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n209_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G127gat), .B(G134gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G113gat), .B(G120gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  NOR3_X1   g029(.A1(new_n227_), .A2(KEYINPUT4), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G225gat), .A2(G233gat), .ZN(new_n233_));
  XOR2_X1   g032(.A(new_n233_), .B(KEYINPUT102), .Z(new_n234_));
  NAND2_X1  g033(.A1(new_n209_), .A2(new_n226_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT100), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(new_n236_), .A3(new_n230_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n209_), .A2(KEYINPUT100), .A3(new_n226_), .ZN(new_n238_));
  XOR2_X1   g037(.A(new_n228_), .B(new_n229_), .Z(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(KEYINPUT100), .B1(new_n209_), .B2(new_n226_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n237_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n242_), .A2(KEYINPUT101), .A3(KEYINPUT4), .ZN(new_n243_));
  AOI21_X1  g042(.A(KEYINPUT101), .B1(new_n242_), .B2(KEYINPUT4), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n232_), .B(new_n234_), .C1(new_n243_), .C2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n242_), .A2(new_n233_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G1gat), .B(G29gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT0), .ZN(new_n248_));
  INV_X1    g047(.A(G57gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(G85gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n245_), .A2(new_n246_), .A3(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT104), .ZN(new_n256_));
  INV_X1    g055(.A(new_n246_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n242_), .A2(KEYINPUT4), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT101), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n242_), .A2(KEYINPUT101), .A3(KEYINPUT4), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n231_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n257_), .B1(new_n262_), .B2(new_n234_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n256_), .B1(new_n263_), .B2(new_n253_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n245_), .A2(new_n246_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(KEYINPUT104), .A3(new_n252_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n255_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G8gat), .B(G36gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT18), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G64gat), .B(G92gat), .ZN(new_n270_));
  XOR2_X1   g069(.A(new_n269_), .B(new_n270_), .Z(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT32), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(G204gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT89), .B1(new_n274_), .B2(G197gat), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT89), .ZN(new_n276_));
  INV_X1    g075(.A(G197gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(new_n277_), .A3(G204gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(G197gat), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n275_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT21), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT90), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n280_), .A2(KEYINPUT90), .A3(KEYINPUT21), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G211gat), .B(G218gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT91), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT91), .ZN(new_n288_));
  INV_X1    g087(.A(G211gat), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n289_), .A2(G218gat), .ZN(new_n290_));
  INV_X1    g089(.A(G218gat), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n291_), .A2(G211gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n288_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G197gat), .B(G204gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT21), .ZN(new_n295_));
  AOI22_X1  g094(.A1(new_n287_), .A2(new_n293_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n287_), .A2(new_n293_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n294_), .A2(new_n295_), .ZN(new_n298_));
  AOI22_X1  g097(.A1(new_n285_), .A2(new_n296_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT25), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(G183gat), .ZN(new_n301_));
  INV_X1    g100(.A(G183gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT25), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT96), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT26), .B(G190gat), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT96), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n301_), .A2(new_n303_), .A3(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n305_), .A2(new_n306_), .A3(new_n308_), .ZN(new_n309_));
  NOR3_X1   g108(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT23), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT82), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT82), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(KEYINPUT23), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n312_), .A2(new_n314_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n311_), .A2(KEYINPUT23), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n310_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  OR2_X1    g118(.A1(G169gat), .A2(G176gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G169gat), .A2(G176gat), .ZN(new_n321_));
  AND3_X1   g120(.A1(new_n321_), .A2(KEYINPUT97), .A3(KEYINPUT24), .ZN(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT97), .B1(new_n321_), .B2(KEYINPUT24), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n320_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n309_), .A2(new_n319_), .A3(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT22), .B(G169gat), .ZN(new_n326_));
  INV_X1    g125(.A(G176gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(new_n321_), .B(KEYINPUT98), .Z(new_n329_));
  NOR2_X1   g128(.A1(new_n311_), .A2(new_n313_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n314_), .A2(new_n316_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n331_), .B1(new_n332_), .B2(new_n312_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(G183gat), .A2(G190gat), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n328_), .B(new_n329_), .C1(new_n333_), .C2(new_n334_), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n325_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n299_), .A2(new_n336_), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n317_), .A2(new_n318_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n321_), .B(new_n328_), .C1(new_n338_), .C2(new_n334_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n320_), .A2(KEYINPUT24), .A3(new_n321_), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT80), .B1(new_n302_), .B2(KEYINPUT25), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n306_), .A2(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(KEYINPUT80), .B1(new_n301_), .B2(new_n303_), .ZN(new_n343_));
  OAI211_X1 g142(.A(KEYINPUT81), .B(new_n340_), .C1(new_n342_), .C2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT82), .B(KEYINPUT23), .ZN(new_n345_));
  AOI211_X1 g144(.A(new_n310_), .B(new_n330_), .C1(new_n345_), .C2(new_n311_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT25), .B(G183gat), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n306_), .B(new_n341_), .C1(new_n348_), .C2(KEYINPUT80), .ZN(new_n349_));
  AOI21_X1  g148(.A(KEYINPUT81), .B1(new_n349_), .B2(new_n340_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n339_), .B1(new_n347_), .B2(new_n350_), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n280_), .A2(KEYINPUT90), .A3(KEYINPUT21), .ZN(new_n352_));
  AOI21_X1  g151(.A(KEYINPUT90), .B1(new_n280_), .B2(KEYINPUT21), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n296_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n297_), .A2(new_n298_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n351_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G226gat), .A2(G233gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n337_), .A2(new_n357_), .A3(KEYINPUT20), .A4(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT20), .B1(new_n299_), .B2(new_n336_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n351_), .A2(new_n356_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n273_), .B(new_n361_), .C1(new_n364_), .C2(new_n360_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n360_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n360_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n337_), .A2(new_n357_), .A3(KEYINPUT20), .A4(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n366_), .A2(new_n368_), .A3(new_n272_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n365_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT103), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT33), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n254_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n271_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n368_), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n351_), .A2(new_n356_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT20), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n325_), .A2(new_n335_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n377_), .B1(new_n356_), .B2(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n367_), .B1(new_n376_), .B2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n374_), .B1(new_n375_), .B2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n366_), .A2(new_n368_), .A3(new_n271_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n381_), .A2(KEYINPUT99), .A3(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT99), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n366_), .A2(new_n368_), .A3(new_n271_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n271_), .B1(new_n366_), .B2(new_n368_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n384_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n253_), .B1(new_n242_), .B2(new_n234_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n233_), .B(new_n232_), .C1(new_n243_), .C2(new_n244_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n373_), .A2(new_n383_), .A3(new_n387_), .A4(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n372_), .B1(new_n254_), .B2(new_n371_), .ZN(new_n392_));
  OAI22_X1  g191(.A1(new_n267_), .A2(new_n370_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n239_), .B(KEYINPUT31), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT85), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT30), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n351_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G15gat), .B(G43gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G71gat), .B(G99gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G227gat), .A2(G233gat), .ZN(new_n403_));
  XOR2_X1   g202(.A(new_n403_), .B(KEYINPUT83), .Z(new_n404_));
  XNOR2_X1  g203(.A(new_n402_), .B(new_n404_), .ZN(new_n405_));
  OAI211_X1 g204(.A(KEYINPUT30), .B(new_n339_), .C1(new_n347_), .C2(new_n350_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n399_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT84), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n399_), .A2(KEYINPUT84), .A3(new_n405_), .A4(new_n406_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n405_), .B1(new_n399_), .B2(new_n406_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n397_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n414_));
  AOI211_X1 g213(.A(new_n412_), .B(new_n396_), .C1(new_n409_), .C2(new_n410_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G78gat), .B(G106gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT88), .B(G233gat), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n419_), .A2(G228gat), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n420_), .A2(KEYINPUT92), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(KEYINPUT92), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n235_), .A2(KEYINPUT29), .ZN(new_n424_));
  AOI211_X1 g223(.A(new_n421_), .B(new_n423_), .C1(new_n356_), .C2(new_n424_), .ZN(new_n425_));
  AND4_X1   g224(.A1(KEYINPUT92), .A2(new_n356_), .A3(new_n424_), .A4(new_n420_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n418_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT93), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT29), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n227_), .A2(KEYINPUT87), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT87), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n431_), .B1(new_n235_), .B2(KEYINPUT29), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT28), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT28), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n430_), .A2(new_n435_), .A3(new_n432_), .ZN(new_n436_));
  XOR2_X1   g235(.A(G22gat), .B(G50gat), .Z(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n434_), .A2(new_n436_), .A3(new_n438_), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n430_), .A2(new_n435_), .A3(new_n432_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n435_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n437_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  AOI22_X1  g241(.A1(new_n427_), .A2(new_n428_), .B1(new_n439_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n421_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n424_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n444_), .B(new_n422_), .C1(new_n299_), .C2(new_n445_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n356_), .A2(KEYINPUT92), .A3(new_n424_), .A4(new_n420_), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n446_), .A2(new_n447_), .A3(new_n417_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n417_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT94), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT94), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n446_), .A2(new_n447_), .A3(new_n417_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n427_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n443_), .A2(new_n450_), .A3(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n443_), .B1(new_n450_), .B2(new_n453_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n416_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n414_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n415_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n461_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n442_), .A2(new_n439_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n463_), .B1(KEYINPUT93), .B2(new_n449_), .ZN(new_n464_));
  NOR3_X1   g263(.A1(new_n448_), .A2(new_n449_), .A3(KEYINPUT94), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n451_), .B1(new_n427_), .B2(new_n452_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n464_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n467_), .A2(new_n416_), .A3(new_n454_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n462_), .A2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(KEYINPUT104), .B1(new_n265_), .B2(new_n252_), .ZN(new_n470_));
  AOI211_X1 g269(.A(new_n256_), .B(new_n253_), .C1(new_n245_), .C2(new_n246_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n254_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT27), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n385_), .A2(new_n473_), .ZN(new_n474_));
  OAI211_X1 g273(.A(new_n374_), .B(new_n361_), .C1(new_n364_), .C2(new_n360_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n381_), .A2(new_n382_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(new_n473_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n472_), .A2(new_n479_), .ZN(new_n480_));
  AOI22_X1  g279(.A1(new_n393_), .A2(new_n458_), .B1(new_n469_), .B2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G29gat), .B(G36gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G43gat), .B(G50gat), .ZN(new_n483_));
  XOR2_X1   g282(.A(new_n482_), .B(new_n483_), .Z(new_n484_));
  XOR2_X1   g283(.A(G1gat), .B(G8gat), .Z(new_n485_));
  INV_X1    g284(.A(G1gat), .ZN(new_n486_));
  INV_X1    g285(.A(G8gat), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT14), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(G22gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(G15gat), .ZN(new_n490_));
  INV_X1    g289(.A(G15gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(G22gat), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n488_), .A2(new_n490_), .A3(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT74), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT74), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n488_), .A2(new_n495_), .A3(new_n490_), .A4(new_n492_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n485_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n494_), .A2(new_n485_), .A3(new_n496_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n484_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n499_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n482_), .B(new_n483_), .ZN(new_n502_));
  NOR3_X1   g301(.A1(new_n501_), .A2(new_n502_), .A3(new_n497_), .ZN(new_n503_));
  OAI211_X1 g302(.A(G229gat), .B(G233gat), .C1(new_n500_), .C2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n484_), .A2(KEYINPUT15), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT15), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n502_), .A2(new_n506_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n505_), .A2(new_n498_), .A3(new_n507_), .A4(new_n499_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n502_), .B1(new_n501_), .B2(new_n497_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G229gat), .A2(G233gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT76), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n508_), .A2(KEYINPUT77), .A3(new_n509_), .A4(new_n511_), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n504_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n508_), .A2(new_n509_), .A3(new_n511_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT77), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  XOR2_X1   g315(.A(G113gat), .B(G141gat), .Z(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT78), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G169gat), .B(G197gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n513_), .A2(KEYINPUT79), .A3(new_n516_), .A4(new_n520_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n516_), .A2(new_n512_), .A3(new_n504_), .A4(new_n520_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT79), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n521_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n513_), .A2(new_n516_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n520_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n525_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G230gat), .A2(G233gat), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT68), .ZN(new_n533_));
  INV_X1    g332(.A(G99gat), .ZN(new_n534_));
  INV_X1    g333(.A(G106gat), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n535_), .A3(KEYINPUT7), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT7), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n537_), .B1(G99gat), .B2(G106gat), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n533_), .B1(new_n539_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n536_), .A2(new_n538_), .ZN(new_n545_));
  AND3_X1   g344(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n546_), .A2(new_n540_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n545_), .A2(new_n547_), .A3(KEYINPUT68), .ZN(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT69), .B(KEYINPUT8), .ZN(new_n549_));
  AND2_X1   g348(.A1(G85gat), .A2(G92gat), .ZN(new_n550_));
  NOR2_X1   g349(.A1(G85gat), .A2(G92gat), .ZN(new_n551_));
  NOR3_X1   g350(.A1(new_n549_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n544_), .A2(new_n548_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n545_), .A2(new_n547_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n550_), .A2(new_n551_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT8), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT9), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n550_), .A2(KEYINPUT67), .A3(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n547_), .A2(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT64), .ZN(new_n563_));
  NAND2_X1  g362(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n562_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n564_), .ZN(new_n566_));
  OAI21_X1  g365(.A(KEYINPUT64), .B1(new_n566_), .B2(new_n561_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT65), .B(G106gat), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n560_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(KEYINPUT67), .B(KEYINPUT9), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n571_), .A2(KEYINPUT66), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(KEYINPUT66), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n572_), .A2(new_n573_), .A3(new_n555_), .ZN(new_n574_));
  AOI22_X1  g373(.A1(new_n553_), .A2(new_n557_), .B1(new_n570_), .B2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT70), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G57gat), .B(G64gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G71gat), .B(G78gat), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n577_), .A2(new_n578_), .A3(KEYINPUT11), .ZN(new_n579_));
  INV_X1    g378(.A(G64gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(G57gat), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n249_), .A2(G64gat), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n581_), .A2(new_n582_), .A3(KEYINPUT11), .ZN(new_n583_));
  AND2_X1   g382(.A1(G71gat), .A2(G78gat), .ZN(new_n584_));
  NOR2_X1   g383(.A1(G71gat), .A2(G78gat), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(KEYINPUT11), .B1(new_n581_), .B2(new_n582_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n576_), .B(new_n579_), .C1(new_n587_), .C2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT11), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n249_), .A2(G64gat), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n580_), .A2(G57gat), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n591_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(new_n583_), .A3(new_n586_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n576_), .B1(new_n595_), .B2(new_n579_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n590_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n575_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n575_), .A2(new_n597_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n532_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT12), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n602_), .B1(new_n575_), .B2(new_n597_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n595_), .A2(KEYINPUT12), .A3(new_n579_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT8), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n606_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n548_), .A2(new_n552_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n607_), .B1(new_n608_), .B2(new_n544_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n570_), .A2(new_n574_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n605_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n603_), .A2(new_n531_), .A3(new_n611_), .A4(new_n598_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n601_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G120gat), .B(G148gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT5), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G176gat), .B(G204gat), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n615_), .B(new_n616_), .Z(new_n617_));
  NAND2_X1  g416(.A1(new_n613_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n617_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n601_), .A2(new_n612_), .A3(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n621_), .A2(KEYINPUT13), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(KEYINPUT13), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n481_), .A2(new_n530_), .A3(new_n625_), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n505_), .B(new_n507_), .C1(new_n609_), .C2(new_n610_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT71), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G232gat), .A2(G233gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT34), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(KEYINPUT35), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n631_), .A2(KEYINPUT35), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n553_), .A2(new_n557_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n570_), .A2(new_n574_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(KEYINPUT72), .B1(new_n636_), .B2(new_n484_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT72), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n575_), .A2(new_n638_), .A3(new_n502_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n633_), .B1(new_n637_), .B2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n629_), .A2(new_n632_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n632_), .B1(new_n629_), .B2(new_n640_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(G190gat), .B(G218gat), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT73), .ZN(new_n645_));
  XNOR2_X1  g444(.A(G134gat), .B(G162gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT36), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n642_), .A2(new_n643_), .A3(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n647_), .B(new_n648_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n629_), .A2(new_n640_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n631_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT35), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n652_), .A2(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n651_), .B1(new_n656_), .B2(new_n641_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n650_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(KEYINPUT37), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n656_), .A2(new_n648_), .A3(new_n647_), .A4(new_n641_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n642_), .A2(new_n643_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n660_), .B1(new_n661_), .B2(new_n651_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT37), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n659_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n498_), .A2(new_n499_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(G231gat), .A2(G233gat), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT75), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n666_), .B(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n595_), .A2(new_n579_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT17), .ZN(new_n672_));
  XOR2_X1   g471(.A(G127gat), .B(G155gat), .Z(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT16), .ZN(new_n674_));
  XNOR2_X1  g473(.A(G183gat), .B(G211gat), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n674_), .B(new_n675_), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n671_), .A2(new_n672_), .A3(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n669_), .A2(new_n670_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n676_), .B(new_n672_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n597_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n669_), .B2(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n682_), .B1(new_n681_), .B2(new_n669_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n679_), .A2(new_n683_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n665_), .A2(new_n684_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n626_), .A2(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n686_), .A2(new_n486_), .A3(new_n472_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT38), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n481_), .A2(new_n658_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n625_), .A2(new_n530_), .A3(new_n684_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(G1gat), .B1(new_n691_), .B2(new_n267_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n688_), .A2(new_n692_), .ZN(G1324gat));
  NAND3_X1  g492(.A1(new_n686_), .A2(new_n487_), .A3(new_n479_), .ZN(new_n694_));
  AOI22_X1  g493(.A1(new_n475_), .A2(new_n474_), .B1(new_n477_), .B2(new_n473_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G8gat), .B1(new_n691_), .B2(new_n695_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n696_), .A2(KEYINPUT39), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n696_), .A2(KEYINPUT39), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n694_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g499(.A(G15gat), .B1(new_n691_), .B2(new_n416_), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n701_), .A2(KEYINPUT41), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(KEYINPUT41), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n686_), .A2(new_n491_), .A3(new_n461_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n702_), .A2(new_n703_), .A3(new_n704_), .ZN(G1326gat));
  NOR2_X1   g504(.A1(new_n455_), .A2(new_n456_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(G22gat), .B1(new_n691_), .B2(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT42), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n686_), .A2(new_n489_), .A3(new_n706_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1327gat));
  INV_X1    g510(.A(new_n684_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n662_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n626_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(G29gat), .B1(new_n715_), .B2(new_n472_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n659_), .A2(new_n664_), .ZN(new_n717_));
  OAI21_X1  g516(.A(KEYINPUT43), .B1(new_n481_), .B2(new_n717_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n467_), .A2(new_n416_), .A3(new_n454_), .ZN(new_n719_));
  AOI22_X1  g518(.A1(new_n467_), .A2(new_n454_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n267_), .B(new_n695_), .C1(new_n719_), .C2(new_n720_), .ZN(new_n721_));
  AND4_X1   g520(.A1(new_n373_), .A2(new_n383_), .A3(new_n387_), .A4(new_n390_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n392_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n370_), .ZN(new_n724_));
  AOI22_X1  g523(.A1(new_n722_), .A2(new_n723_), .B1(new_n472_), .B2(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n721_), .B1(new_n725_), .B2(new_n457_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n726_), .A2(new_n727_), .A3(new_n665_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n718_), .A2(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n624_), .A2(new_n529_), .A3(new_n684_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT105), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n734_), .A2(G29gat), .A3(new_n472_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n729_), .A2(KEYINPUT44), .A3(new_n731_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n716_), .B1(new_n735_), .B2(new_n736_), .ZN(G1328gat));
  NOR3_X1   g536(.A1(new_n714_), .A2(G36gat), .A3(new_n695_), .ZN(new_n738_));
  XOR2_X1   g537(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n739_));
  XNOR2_X1  g538(.A(new_n738_), .B(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(G36gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(KEYINPUT44), .B1(new_n729_), .B2(new_n731_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n743_), .A2(new_n695_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n742_), .B1(new_n744_), .B2(new_n736_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n741_), .A2(KEYINPUT46), .A3(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT46), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n748_), .B1(new_n740_), .B2(new_n745_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1329gat));
  NAND3_X1  g549(.A1(new_n734_), .A2(G43gat), .A3(new_n461_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n736_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n714_), .A2(new_n416_), .ZN(new_n753_));
  OAI22_X1  g552(.A1(new_n751_), .A2(new_n752_), .B1(G43gat), .B2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g554(.A(G50gat), .B1(new_n715_), .B2(new_n706_), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n734_), .A2(G50gat), .A3(new_n706_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n757_), .B2(new_n736_), .ZN(G1331gat));
  NOR3_X1   g557(.A1(new_n624_), .A2(new_n529_), .A3(new_n684_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n689_), .A2(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(G57gat), .B1(new_n760_), .B2(new_n267_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n393_), .A2(new_n458_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n529_), .B1(new_n762_), .B2(new_n721_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n624_), .B1(new_n763_), .B2(KEYINPUT107), .ZN(new_n764_));
  AOI21_X1  g563(.A(KEYINPUT107), .B1(new_n726_), .B2(new_n530_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n764_), .A2(new_n685_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n472_), .A2(new_n249_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n761_), .B1(new_n767_), .B2(new_n768_), .ZN(G1332gat));
  INV_X1    g568(.A(new_n760_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n479_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(G64gat), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT109), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n771_), .A2(new_n774_), .A3(G64gat), .ZN(new_n775_));
  XOR2_X1   g574(.A(KEYINPUT108), .B(KEYINPUT48), .Z(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n773_), .A2(new_n775_), .A3(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n773_), .B2(new_n775_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n479_), .A2(new_n580_), .ZN(new_n780_));
  OAI22_X1  g579(.A1(new_n778_), .A2(new_n779_), .B1(new_n767_), .B2(new_n780_), .ZN(G1333gat));
  OAI21_X1  g580(.A(G71gat), .B1(new_n760_), .B2(new_n416_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT49), .ZN(new_n783_));
  OR2_X1    g582(.A1(new_n416_), .A2(G71gat), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n783_), .B1(new_n767_), .B2(new_n784_), .ZN(G1334gat));
  INV_X1    g584(.A(KEYINPUT50), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n770_), .A2(new_n706_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n787_), .B2(G78gat), .ZN(new_n788_));
  INV_X1    g587(.A(G78gat), .ZN(new_n789_));
  AOI211_X1 g588(.A(KEYINPUT50), .B(new_n789_), .C1(new_n770_), .C2(new_n706_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n706_), .A2(new_n789_), .ZN(new_n791_));
  OAI22_X1  g590(.A1(new_n788_), .A2(new_n790_), .B1(new_n767_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT110), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n792_), .B(new_n793_), .ZN(G1335gat));
  NAND3_X1  g593(.A1(new_n625_), .A2(new_n530_), .A3(new_n684_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n718_), .B2(new_n728_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n797_));
  OR2_X1    g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n797_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n267_), .A2(new_n251_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(KEYINPUT112), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n798_), .A2(new_n799_), .A3(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n264_), .A2(new_n266_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n803_), .A2(new_n254_), .A3(new_n695_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n468_), .B2(new_n462_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n472_), .A2(new_n724_), .ZN(new_n806_));
  AOI22_X1  g605(.A1(new_n477_), .A2(new_n384_), .B1(new_n389_), .B2(new_n388_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n723_), .A2(new_n807_), .A3(new_n373_), .A4(new_n383_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n457_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n809_));
  OAI211_X1 g608(.A(KEYINPUT107), .B(new_n530_), .C1(new_n805_), .C2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n625_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n713_), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n811_), .A2(new_n765_), .A3(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(G85gat), .B1(new_n813_), .B2(new_n472_), .ZN(new_n814_));
  OR3_X1    g613(.A1(new_n802_), .A2(KEYINPUT113), .A3(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(KEYINPUT113), .B1(new_n802_), .B2(new_n814_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(G1336gat));
  AOI21_X1  g616(.A(G92gat), .B1(new_n813_), .B2(new_n479_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n798_), .A2(new_n799_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n479_), .A2(G92gat), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n818_), .B1(new_n819_), .B2(new_n820_), .ZN(G1337gat));
  NAND2_X1  g620(.A1(new_n461_), .A2(new_n568_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n764_), .A2(new_n766_), .A3(new_n713_), .A4(new_n823_), .ZN(new_n824_));
  XOR2_X1   g623(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n825_));
  AOI211_X1 g624(.A(new_n416_), .B(new_n795_), .C1(new_n718_), .C2(new_n728_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n824_), .B(new_n825_), .C1(new_n826_), .C2(new_n534_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT115), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n534_), .B1(new_n796_), .B2(new_n461_), .ZN(new_n829_));
  NOR4_X1   g628(.A1(new_n811_), .A2(new_n765_), .A3(new_n812_), .A4(new_n822_), .ZN(new_n830_));
  OAI21_X1  g629(.A(KEYINPUT114), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT114), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n824_), .B(new_n832_), .C1(new_n826_), .C2(new_n534_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n828_), .B1(new_n834_), .B2(KEYINPUT51), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT51), .ZN(new_n836_));
  AOI211_X1 g635(.A(KEYINPUT115), .B(new_n836_), .C1(new_n831_), .C2(new_n833_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n827_), .B1(new_n835_), .B2(new_n837_), .ZN(G1338gat));
  NAND3_X1  g637(.A1(new_n813_), .A2(new_n569_), .A3(new_n706_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT52), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n796_), .A2(new_n706_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n840_), .B1(new_n841_), .B2(G106gat), .ZN(new_n842_));
  AOI211_X1 g641(.A(KEYINPUT52), .B(new_n535_), .C1(new_n796_), .C2(new_n706_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n839_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g644(.A1(new_n625_), .A2(new_n529_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n846_), .A2(new_n712_), .A3(new_n664_), .A4(new_n659_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n717_), .A2(KEYINPUT54), .A3(new_n712_), .A4(new_n846_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT56), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT118), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n603_), .A2(new_n598_), .A3(new_n611_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n532_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT55), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(new_n612_), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT117), .B1(new_n612_), .B2(new_n856_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n612_), .A2(KEYINPUT117), .A3(new_n856_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n857_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n853_), .B1(new_n861_), .B2(new_n619_), .ZN(new_n862_));
  OR2_X1    g661(.A1(new_n612_), .A2(new_n856_), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n612_), .A2(KEYINPUT117), .A3(new_n856_), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n863_), .B(new_n855_), .C1(new_n864_), .C2(new_n858_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n865_), .A2(KEYINPUT118), .A3(new_n852_), .A4(new_n617_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n620_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n867_), .B1(new_n525_), .B2(new_n528_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n862_), .A2(new_n866_), .A3(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n511_), .B1(new_n500_), .B2(new_n503_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n508_), .A2(new_n509_), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n870_), .B(new_n527_), .C1(new_n871_), .C2(new_n511_), .ZN(new_n872_));
  AND2_X1   g671(.A1(new_n525_), .A2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n621_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n869_), .A2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(KEYINPUT57), .B1(new_n875_), .B2(new_n662_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877_));
  AOI211_X1 g676(.A(new_n877_), .B(new_n658_), .C1(new_n869_), .C2(new_n874_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n876_), .A2(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n865_), .A2(KEYINPUT56), .A3(new_n617_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(KEYINPUT119), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n865_), .A2(new_n882_), .A3(KEYINPUT56), .A4(new_n617_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n852_), .B1(new_n861_), .B2(new_n619_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n881_), .A2(new_n883_), .A3(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n873_), .A2(new_n620_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NAND4_X1  g686(.A1(new_n885_), .A2(KEYINPUT120), .A3(new_n887_), .A4(KEYINPUT58), .ZN(new_n888_));
  AOI21_X1  g687(.A(KEYINPUT56), .B1(new_n865_), .B2(new_n617_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n889_), .B1(KEYINPUT119), .B2(new_n880_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n886_), .B1(new_n890_), .B2(new_n883_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n888_), .B(new_n665_), .C1(new_n891_), .C2(KEYINPUT58), .ZN(new_n892_));
  AOI21_X1  g691(.A(KEYINPUT120), .B1(new_n891_), .B2(KEYINPUT58), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n879_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n851_), .B1(new_n894_), .B2(new_n684_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n720_), .A2(new_n472_), .A3(new_n695_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(KEYINPUT121), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n895_), .A2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(G113gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n898_), .A2(new_n899_), .A3(new_n529_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(KEYINPUT59), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n902_), .B1(new_n895_), .B2(new_n897_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n530_), .B1(new_n901_), .B2(new_n903_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n900_), .B1(new_n904_), .B2(new_n899_), .ZN(G1340gat));
  INV_X1    g704(.A(KEYINPUT60), .ZN(new_n906_));
  INV_X1    g705(.A(G120gat), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n625_), .A2(new_n906_), .A3(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n908_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n898_), .A2(new_n909_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n624_), .B1(new_n901_), .B2(new_n903_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n911_), .B2(new_n907_), .ZN(G1341gat));
  INV_X1    g711(.A(G127gat), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n898_), .A2(new_n913_), .A3(new_n712_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n684_), .B1(new_n901_), .B2(new_n903_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n915_), .B2(new_n913_), .ZN(G1342gat));
  AOI21_X1  g715(.A(G134gat), .B1(new_n898_), .B2(new_n658_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n901_), .A2(new_n903_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(KEYINPUT122), .B(G134gat), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n717_), .A2(new_n919_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n917_), .B1(new_n918_), .B2(new_n920_), .ZN(G1343gat));
  INV_X1    g720(.A(new_n895_), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n267_), .A2(new_n468_), .A3(new_n479_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(KEYINPUT123), .ZN(new_n924_));
  AND2_X1   g723(.A1(new_n922_), .A2(new_n924_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n529_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(G141gat), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n925_), .A2(new_n211_), .A3(new_n529_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(G1344gat));
  NAND2_X1  g728(.A1(new_n925_), .A2(new_n625_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(G148gat), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n925_), .A2(new_n212_), .A3(new_n625_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1345gat));
  NAND3_X1  g732(.A1(new_n885_), .A2(KEYINPUT58), .A3(new_n887_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT120), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n885_), .A2(new_n887_), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT58), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n937_), .A2(new_n938_), .ZN(new_n939_));
  NAND4_X1  g738(.A1(new_n936_), .A2(new_n939_), .A3(new_n665_), .A4(new_n888_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n712_), .B1(new_n940_), .B2(new_n879_), .ZN(new_n941_));
  OAI211_X1 g740(.A(new_n924_), .B(new_n712_), .C1(new_n941_), .C2(new_n851_), .ZN(new_n942_));
  OR2_X1    g741(.A1(new_n942_), .A2(KEYINPUT124), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(KEYINPUT124), .ZN(new_n944_));
  XOR2_X1   g743(.A(KEYINPUT61), .B(G155gat), .Z(new_n945_));
  AND3_X1   g744(.A1(new_n943_), .A2(new_n944_), .A3(new_n945_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n945_), .B1(new_n943_), .B2(new_n944_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n946_), .A2(new_n947_), .ZN(G1346gat));
  NAND3_X1  g747(.A1(new_n922_), .A2(new_n658_), .A3(new_n924_), .ZN(new_n949_));
  INV_X1    g748(.A(KEYINPUT125), .ZN(new_n950_));
  AND3_X1   g749(.A1(new_n949_), .A2(new_n950_), .A3(new_n223_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n950_), .B1(new_n949_), .B2(new_n223_), .ZN(new_n952_));
  NAND4_X1  g751(.A1(new_n922_), .A2(G162gat), .A3(new_n665_), .A4(new_n924_), .ZN(new_n953_));
  INV_X1    g752(.A(new_n953_), .ZN(new_n954_));
  NOR3_X1   g753(.A1(new_n951_), .A2(new_n952_), .A3(new_n954_), .ZN(G1347gat));
  NOR2_X1   g754(.A1(new_n472_), .A2(new_n695_), .ZN(new_n956_));
  INV_X1    g755(.A(new_n956_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n957_), .A2(new_n416_), .ZN(new_n958_));
  OAI211_X1 g757(.A(new_n707_), .B(new_n958_), .C1(new_n941_), .C2(new_n851_), .ZN(new_n959_));
  OR2_X1    g758(.A1(new_n959_), .A2(new_n530_), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n960_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n961_));
  OAI21_X1  g760(.A(G169gat), .B1(new_n959_), .B2(new_n530_), .ZN(new_n962_));
  INV_X1    g761(.A(KEYINPUT62), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n962_), .A2(new_n963_), .ZN(new_n964_));
  INV_X1    g763(.A(new_n326_), .ZN(new_n965_));
  OAI211_X1 g764(.A(new_n961_), .B(new_n964_), .C1(new_n965_), .C2(new_n960_), .ZN(G1348gat));
  OAI21_X1  g765(.A(KEYINPUT126), .B1(new_n895_), .B2(new_n706_), .ZN(new_n967_));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n968_));
  OAI211_X1 g767(.A(new_n968_), .B(new_n707_), .C1(new_n941_), .C2(new_n851_), .ZN(new_n969_));
  NOR4_X1   g768(.A1(new_n957_), .A2(new_n327_), .A3(new_n416_), .A4(new_n624_), .ZN(new_n970_));
  NAND3_X1  g769(.A1(new_n967_), .A2(new_n969_), .A3(new_n970_), .ZN(new_n971_));
  OAI21_X1  g770(.A(new_n327_), .B1(new_n959_), .B2(new_n624_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n971_), .A2(new_n972_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n973_), .A2(KEYINPUT127), .ZN(new_n974_));
  INV_X1    g773(.A(KEYINPUT127), .ZN(new_n975_));
  NAND3_X1  g774(.A1(new_n971_), .A2(new_n975_), .A3(new_n972_), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n974_), .A2(new_n976_), .ZN(G1349gat));
  AOI211_X1 g776(.A(new_n684_), .B(new_n959_), .C1(new_n305_), .C2(new_n308_), .ZN(new_n978_));
  NAND4_X1  g777(.A1(new_n967_), .A2(new_n712_), .A3(new_n958_), .A4(new_n969_), .ZN(new_n979_));
  AOI21_X1  g778(.A(new_n978_), .B1(new_n302_), .B2(new_n979_), .ZN(G1350gat));
  OAI21_X1  g779(.A(G190gat), .B1(new_n959_), .B2(new_n717_), .ZN(new_n981_));
  NAND2_X1  g780(.A1(new_n658_), .A2(new_n306_), .ZN(new_n982_));
  OAI21_X1  g781(.A(new_n981_), .B1(new_n959_), .B2(new_n982_), .ZN(G1351gat));
  NOR3_X1   g782(.A1(new_n895_), .A2(new_n468_), .A3(new_n957_), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n984_), .A2(new_n529_), .ZN(new_n985_));
  XNOR2_X1  g784(.A(new_n985_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g785(.A1(new_n984_), .A2(new_n625_), .ZN(new_n987_));
  XNOR2_X1  g786(.A(new_n987_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g787(.A1(new_n984_), .A2(new_n712_), .ZN(new_n989_));
  OAI21_X1  g788(.A(new_n989_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n990_));
  XOR2_X1   g789(.A(KEYINPUT63), .B(G211gat), .Z(new_n991_));
  OAI21_X1  g790(.A(new_n990_), .B1(new_n989_), .B2(new_n991_), .ZN(G1354gat));
  NAND3_X1  g791(.A1(new_n984_), .A2(new_n291_), .A3(new_n658_), .ZN(new_n993_));
  NAND2_X1  g792(.A1(new_n984_), .A2(new_n665_), .ZN(new_n994_));
  INV_X1    g793(.A(new_n994_), .ZN(new_n995_));
  OAI21_X1  g794(.A(new_n993_), .B1(new_n995_), .B2(new_n291_), .ZN(G1355gat));
endmodule


