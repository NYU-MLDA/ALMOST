//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 0 0 0 1 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n601_, new_n602_, new_n603_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n810_, new_n811_, new_n812_, new_n814_,
    new_n815_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n824_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT10), .ZN(new_n203_));
  INV_X1    g002(.A(G99gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT64), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n205_), .A2(new_n215_), .A3(new_n206_), .A4(new_n207_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n209_), .A2(new_n214_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G85gat), .ZN(new_n218_));
  INV_X1    g017(.A(G92gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(KEYINPUT9), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT9), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(G85gat), .A3(G92gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT65), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT65), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n222_), .A2(new_n227_), .A3(new_n224_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n217_), .B1(new_n226_), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT66), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT8), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n220_), .A2(new_n231_), .A3(new_n221_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT7), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n233_), .A2(new_n204_), .A3(new_n206_), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  AOI211_X1 g035(.A(new_n230_), .B(new_n232_), .C1(new_n236_), .C2(new_n214_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n214_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n232_), .ZN(new_n239_));
  AOI21_X1  g038(.A(KEYINPUT66), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n237_), .A2(new_n240_), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n211_), .A2(new_n213_), .A3(KEYINPUT67), .ZN(new_n242_));
  AOI21_X1  g041(.A(KEYINPUT67), .B1(new_n211_), .B2(new_n213_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n234_), .A2(new_n235_), .ZN(new_n244_));
  NOR3_X1   g043(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n221_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(G85gat), .A2(G92gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT8), .B1(new_n245_), .B2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n229_), .B1(new_n241_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(G50gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(G43gat), .ZN(new_n253_));
  INV_X1    g052(.A(G43gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(G50gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(G36gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(G29gat), .ZN(new_n258_));
  INV_X1    g057(.A(G29gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(G36gat), .ZN(new_n260_));
  AND3_X1   g059(.A1(new_n258_), .A2(new_n260_), .A3(KEYINPUT72), .ZN(new_n261_));
  AOI21_X1  g060(.A(KEYINPUT72), .B1(new_n258_), .B2(new_n260_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n256_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT72), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n259_), .A2(G36gat), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n257_), .A2(G29gat), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n264_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n258_), .A2(new_n260_), .A3(KEYINPUT72), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n253_), .A2(new_n255_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n267_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n263_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n251_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(KEYINPUT15), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n226_), .A2(new_n228_), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n216_), .A2(new_n214_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n274_), .A2(new_n209_), .A3(new_n275_), .ZN(new_n276_));
  AND2_X1   g075(.A1(new_n211_), .A2(new_n213_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n239_), .B1(new_n277_), .B2(new_n244_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(new_n230_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n238_), .A2(KEYINPUT66), .A3(new_n239_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT67), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n214_), .A2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n211_), .A2(new_n213_), .A3(KEYINPUT67), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n283_), .A2(new_n284_), .A3(new_n236_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n231_), .B1(new_n285_), .B2(new_n248_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n276_), .B1(new_n281_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n273_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G232gat), .A2(G233gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT34), .ZN(new_n290_));
  OAI211_X1 g089(.A(new_n272_), .B(new_n288_), .C1(KEYINPUT35), .C2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(KEYINPUT35), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G190gat), .B(G218gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G134gat), .B(G162gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n296_), .A2(KEYINPUT36), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n296_), .A2(KEYINPUT36), .ZN(new_n298_));
  NOR3_X1   g097(.A1(new_n293_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n293_), .A2(new_n297_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT25), .B(G183gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT26), .B(G190gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT83), .ZN(new_n305_));
  INV_X1    g104(.A(G183gat), .ZN(new_n306_));
  INV_X1    g105(.A(G190gat), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT23), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT23), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n309_), .A2(G183gat), .A3(G190gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n312_), .B1(G169gat), .B2(G176gat), .ZN(new_n313_));
  NOR3_X1   g112(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n305_), .A2(new_n311_), .A3(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(G169gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n310_), .A2(KEYINPUT84), .ZN(new_n319_));
  XOR2_X1   g118(.A(new_n319_), .B(new_n308_), .Z(new_n320_));
  NOR2_X1   g119(.A1(G183gat), .A2(G190gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n318_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n316_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G71gat), .B(G99gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(G43gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n323_), .B(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(G127gat), .B(G134gat), .Z(new_n327_));
  XOR2_X1   g126(.A(G113gat), .B(G120gat), .Z(new_n328_));
  XOR2_X1   g127(.A(new_n327_), .B(new_n328_), .Z(new_n329_));
  XNOR2_X1  g128(.A(new_n326_), .B(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G227gat), .A2(G233gat), .ZN(new_n331_));
  INV_X1    g130(.A(G15gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT30), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT31), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n330_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n330_), .A2(new_n335_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G155gat), .A2(G162gat), .ZN(new_n340_));
  NOR2_X1   g139(.A1(G155gat), .A2(G162gat), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(G141gat), .A2(G148gat), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n343_), .B(KEYINPUT3), .Z(new_n344_));
  NAND2_X1  g143(.A1(G141gat), .A2(G148gat), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n345_), .B(KEYINPUT2), .Z(new_n346_));
  OAI211_X1 g145(.A(new_n340_), .B(new_n342_), .C1(new_n344_), .C2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n341_), .B1(KEYINPUT1), .B2(new_n340_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n348_), .B1(KEYINPUT1), .B2(new_n340_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n343_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(new_n350_), .A3(new_n345_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n347_), .A2(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n352_), .A2(KEYINPUT29), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G22gat), .B(G50gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT28), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n353_), .B(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(G204gat), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n357_), .A2(G197gat), .ZN(new_n358_));
  INV_X1    g157(.A(G197gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n359_), .A2(G204gat), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT21), .B1(new_n358_), .B2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G211gat), .B(G218gat), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT86), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n360_), .B1(new_n363_), .B2(new_n358_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT86), .B1(new_n357_), .B2(G197gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  XOR2_X1   g165(.A(KEYINPUT87), .B(KEYINPUT21), .Z(new_n367_));
  OAI211_X1 g166(.A(new_n361_), .B(new_n362_), .C1(new_n366_), .C2(new_n367_), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n362_), .A2(KEYINPUT88), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n362_), .A2(KEYINPUT88), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n366_), .A2(new_n369_), .A3(KEYINPUT21), .A4(new_n370_), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n352_), .A2(KEYINPUT29), .B1(new_n368_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(G228gat), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n373_), .A2(KEYINPUT85), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n373_), .A2(KEYINPUT85), .ZN(new_n375_));
  OAI21_X1  g174(.A(G233gat), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n372_), .B(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G78gat), .B(G106gat), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n356_), .B1(new_n379_), .B2(KEYINPUT89), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n377_), .B(new_n378_), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n380_), .A2(new_n381_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n329_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(new_n351_), .A3(new_n347_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n352_), .A2(new_n329_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G225gat), .A2(G233gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT97), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  XOR2_X1   g192(.A(G1gat), .B(G29gat), .Z(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT96), .B(G85gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT0), .B(G57gat), .ZN(new_n397_));
  XOR2_X1   g196(.A(new_n396_), .B(new_n397_), .Z(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n387_), .A2(KEYINPUT4), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n388_), .A2(KEYINPUT95), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n393_), .B(new_n399_), .C1(new_n390_), .C2(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(KEYINPUT98), .A2(KEYINPUT33), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n390_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n399_), .B1(new_n389_), .B2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n407_), .B1(new_n402_), .B2(new_n406_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n403_), .A2(new_n404_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n405_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n311_), .B1(G183gat), .B2(G190gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(new_n318_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n315_), .A2(new_n304_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n412_), .B1(new_n320_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n368_), .A2(new_n371_), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT20), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n416_), .B1(new_n323_), .B2(new_n415_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G226gat), .A2(G233gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n417_), .A2(new_n421_), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n422_), .A2(KEYINPUT92), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n414_), .A2(KEYINPUT91), .A3(new_n415_), .ZN(new_n424_));
  AOI21_X1  g223(.A(KEYINPUT91), .B1(new_n414_), .B2(new_n415_), .ZN(new_n425_));
  OAI221_X1 g224(.A(KEYINPUT20), .B1(new_n323_), .B2(new_n415_), .C1(new_n424_), .C2(new_n425_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n426_), .A2(new_n420_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n422_), .A2(KEYINPUT92), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n423_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  XOR2_X1   g228(.A(G8gat), .B(G36gat), .Z(new_n430_));
  XNOR2_X1  g229(.A(G64gat), .B(G92gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  OR3_X1    g233(.A1(new_n429_), .A2(KEYINPUT94), .A3(new_n434_), .ZN(new_n435_));
  OR2_X1    g234(.A1(new_n429_), .A2(new_n434_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n429_), .A2(new_n434_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(KEYINPUT94), .A3(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n410_), .B1(new_n435_), .B2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n417_), .A2(new_n421_), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n426_), .A2(new_n420_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n440_), .B1(new_n441_), .B2(KEYINPUT99), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n442_), .B1(KEYINPUT99), .B2(new_n441_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n434_), .A2(KEYINPUT32), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n393_), .B1(new_n390_), .B2(new_n402_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n398_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n403_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n429_), .A2(new_n444_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n446_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n385_), .B1(new_n439_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT27), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n438_), .A2(new_n435_), .A3(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n449_), .ZN(new_n455_));
  XOR2_X1   g254(.A(new_n434_), .B(KEYINPUT100), .Z(new_n456_));
  NAND2_X1  g255(.A1(new_n443_), .A2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n457_), .A2(KEYINPUT27), .A3(new_n437_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n454_), .A2(new_n384_), .A3(new_n455_), .A4(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n339_), .B1(new_n452_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT101), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n454_), .A2(new_n458_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n462_), .A2(new_n384_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n449_), .A2(new_n338_), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n460_), .A2(new_n461_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n452_), .A2(new_n459_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n338_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT101), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n301_), .B1(new_n465_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G230gat), .A2(G233gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G57gat), .B(G64gat), .ZN(new_n471_));
  OR2_X1    g270(.A1(new_n471_), .A2(KEYINPUT11), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(KEYINPUT11), .ZN(new_n473_));
  XOR2_X1   g272(.A(G71gat), .B(G78gat), .Z(new_n474_));
  NAND3_X1  g273(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n473_), .A2(new_n474_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT68), .B1(new_n287_), .B2(new_n478_), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n276_), .B(new_n477_), .C1(new_n281_), .C2(new_n286_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n470_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n481_), .B1(new_n480_), .B2(new_n479_), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT12), .B1(new_n251_), .B2(new_n477_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT12), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n287_), .A2(new_n484_), .A3(new_n478_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n480_), .A2(new_n470_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT69), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n480_), .A2(KEYINPUT69), .A3(new_n470_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n486_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n482_), .A2(new_n491_), .ZN(new_n492_));
  XOR2_X1   g291(.A(G120gat), .B(G148gat), .Z(new_n493_));
  XNOR2_X1  g292(.A(G176gat), .B(G204gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(KEYINPUT70), .B(KEYINPUT5), .Z(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n492_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n492_), .A2(new_n497_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n502_), .A2(KEYINPUT13), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(KEYINPUT13), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G113gat), .B(G141gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT81), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G169gat), .B(G197gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n507_), .B(new_n508_), .Z(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G229gat), .A2(G233gat), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT77), .ZN(new_n513_));
  NOR3_X1   g312(.A1(new_n261_), .A2(new_n262_), .A3(new_n256_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n269_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n513_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G15gat), .B(G22gat), .ZN(new_n517_));
  INV_X1    g316(.A(G8gat), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  XOR2_X1   g319(.A(G1gat), .B(G8gat), .Z(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n263_), .A2(new_n270_), .A3(KEYINPUT77), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n516_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT78), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT78), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n516_), .A2(new_n526_), .A3(new_n522_), .A4(new_n523_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n522_), .B1(new_n516_), .B2(new_n523_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(KEYINPUT79), .B1(new_n528_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT79), .ZN(new_n532_));
  AOI211_X1 g331(.A(new_n532_), .B(new_n529_), .C1(new_n525_), .C2(new_n527_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n512_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n522_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n273_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n528_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  AOI22_X1  g337(.A1(new_n534_), .A2(KEYINPUT80), .B1(new_n511_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT80), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n540_), .B(new_n512_), .C1(new_n531_), .C2(new_n533_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n510_), .B1(new_n539_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n534_), .A2(KEYINPUT80), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n538_), .A2(new_n511_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n543_), .A2(new_n541_), .A3(new_n544_), .A4(new_n510_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT82), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT82), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n539_), .A2(new_n547_), .A3(new_n541_), .A4(new_n510_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n542_), .B1(new_n546_), .B2(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n505_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G183gat), .B(G211gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT75), .ZN(new_n553_));
  XOR2_X1   g352(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(G127gat), .B(G155gat), .Z(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT17), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n477_), .B(new_n522_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G231gat), .A2(G233gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n558_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n561_), .A2(KEYINPUT17), .A3(new_n557_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n551_), .A2(new_n564_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n469_), .A2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n202_), .B1(new_n566_), .B2(new_n449_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n549_), .B1(new_n465_), .B2(new_n468_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(KEYINPUT73), .A2(KEYINPUT37), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n301_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(KEYINPUT73), .A2(KEYINPUT37), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n572_), .A2(new_n564_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT76), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n505_), .B(KEYINPUT71), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n568_), .A2(new_n577_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n578_), .A2(new_n202_), .A3(new_n449_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n579_), .A2(KEYINPUT102), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(KEYINPUT102), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n567_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT104), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n587_), .B1(new_n582_), .B2(new_n584_), .ZN(new_n588_));
  AOI211_X1 g387(.A(KEYINPUT104), .B(new_n585_), .C1(new_n580_), .C2(new_n581_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n586_), .B1(new_n588_), .B2(new_n589_), .ZN(G1324gat));
  NAND3_X1  g389(.A1(new_n578_), .A2(new_n518_), .A3(new_n462_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n566_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n462_), .ZN(new_n593_));
  OAI21_X1  g392(.A(G8gat), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n594_), .A2(KEYINPUT39), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n594_), .A2(KEYINPUT39), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n591_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n597_), .B(new_n599_), .ZN(G1325gat));
  AOI21_X1  g399(.A(new_n332_), .B1(new_n566_), .B2(new_n339_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT41), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n578_), .A2(new_n332_), .A3(new_n339_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(G1326gat));
  INV_X1    g403(.A(G22gat), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n605_), .B1(new_n566_), .B2(new_n384_), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n606_), .B(KEYINPUT42), .Z(new_n607_));
  NAND3_X1  g406(.A1(new_n578_), .A2(new_n605_), .A3(new_n384_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(G1327gat));
  INV_X1    g408(.A(new_n301_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n564_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n505_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n568_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(G29gat), .B1(new_n614_), .B2(new_n449_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n551_), .A2(new_n611_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT43), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n465_), .A2(new_n468_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n617_), .B1(new_n618_), .B2(new_n572_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n572_), .ZN(new_n620_));
  AOI211_X1 g419(.A(KEYINPUT43), .B(new_n620_), .C1(new_n465_), .C2(new_n468_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n616_), .B1(new_n619_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT44), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT106), .ZN(new_n625_));
  INV_X1    g424(.A(new_n616_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n463_), .A2(new_n464_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n627_), .B1(new_n467_), .B2(KEYINPUT101), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n460_), .A2(new_n461_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n572_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT43), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n618_), .A2(new_n617_), .A3(new_n572_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n626_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n625_), .B1(new_n633_), .B2(KEYINPUT44), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n622_), .A2(KEYINPUT106), .A3(new_n623_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n624_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n455_), .A2(new_n259_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n615_), .B1(new_n636_), .B2(new_n637_), .ZN(G1328gat));
  INV_X1    g437(.A(KEYINPUT107), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n639_), .A2(KEYINPUT46), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n257_), .B1(new_n636_), .B2(new_n462_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n613_), .A2(G36gat), .A3(new_n593_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT45), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n640_), .B1(new_n641_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n640_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n643_), .ZN(new_n646_));
  AOI211_X1 g445(.A(new_n593_), .B(new_n624_), .C1(new_n634_), .C2(new_n635_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n645_), .B(new_n646_), .C1(new_n647_), .C2(new_n257_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n644_), .A2(new_n648_), .ZN(G1329gat));
  NOR2_X1   g448(.A1(new_n338_), .A2(new_n254_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n636_), .A2(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n254_), .B1(new_n613_), .B2(new_n338_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT108), .Z(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT47), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT47), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n651_), .A2(new_n656_), .A3(new_n653_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(G1330gat));
  AND2_X1   g457(.A1(new_n636_), .A2(new_n384_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n384_), .A2(new_n252_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT109), .ZN(new_n661_));
  OAI22_X1  g460(.A1(new_n659_), .A2(new_n252_), .B1(new_n613_), .B2(new_n661_), .ZN(G1331gat));
  NAND4_X1  g461(.A1(new_n469_), .A2(new_n549_), .A3(new_n611_), .A4(new_n576_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G57gat), .B1(new_n663_), .B2(new_n455_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n546_), .A2(new_n548_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n542_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n667_), .B1(new_n465_), .B2(new_n468_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n505_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n574_), .A2(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(G57gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n671_), .A2(new_n672_), .A3(new_n449_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n664_), .A2(new_n673_), .ZN(G1332gat));
  OAI21_X1  g473(.A(G64gat), .B1(new_n663_), .B2(new_n593_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT48), .ZN(new_n676_));
  INV_X1    g475(.A(G64gat), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n671_), .A2(new_n677_), .A3(new_n462_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(G1333gat));
  OAI21_X1  g478(.A(G71gat), .B1(new_n663_), .B2(new_n338_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT49), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n338_), .A2(G71gat), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT110), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n671_), .A2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n681_), .A2(new_n684_), .ZN(G1334gat));
  OAI21_X1  g484(.A(G78gat), .B1(new_n663_), .B2(new_n385_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT50), .ZN(new_n687_));
  INV_X1    g486(.A(G78gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n671_), .A2(new_n688_), .A3(new_n384_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(G1335gat));
  NAND3_X1  g489(.A1(new_n505_), .A2(new_n549_), .A3(new_n564_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT111), .Z(new_n692_));
  OAI21_X1  g491(.A(new_n692_), .B1(new_n619_), .B2(new_n621_), .ZN(new_n693_));
  OAI21_X1  g492(.A(G85gat), .B1(new_n693_), .B2(new_n455_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n668_), .A2(new_n301_), .A3(new_n564_), .A4(new_n576_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n449_), .A2(new_n218_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n694_), .B1(new_n695_), .B2(new_n696_), .ZN(G1336gat));
  OAI21_X1  g496(.A(G92gat), .B1(new_n693_), .B2(new_n593_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n462_), .A2(new_n219_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n698_), .B1(new_n695_), .B2(new_n699_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT112), .Z(G1337gat));
  OAI21_X1  g500(.A(G99gat), .B1(new_n693_), .B2(new_n338_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n339_), .A2(new_n205_), .A3(new_n207_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n695_), .B2(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI211_X1 g504(.A(new_n384_), .B(new_n692_), .C1(new_n619_), .C2(new_n621_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT52), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n706_), .A2(new_n707_), .A3(G106gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n706_), .B2(G106gat), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n384_), .A2(new_n206_), .ZN(new_n710_));
  OAI22_X1  g509(.A1(new_n708_), .A2(new_n709_), .B1(new_n695_), .B2(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT53), .ZN(G1339gat));
  XNOR2_X1  g511(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n713_));
  INV_X1    g512(.A(new_n485_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n484_), .B1(new_n287_), .B2(new_n478_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n480_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n470_), .ZN(new_n717_));
  AOI22_X1  g516(.A1(new_n491_), .A2(new_n713_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n486_), .A2(KEYINPUT55), .A3(new_n489_), .A4(new_n490_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n719_), .A2(KEYINPUT115), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(KEYINPUT115), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n718_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT116), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT116), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n724_), .B(new_n718_), .C1(new_n720_), .C2(new_n721_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n723_), .A2(new_n497_), .A3(new_n725_), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n726_), .A2(KEYINPUT56), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n509_), .B1(new_n537_), .B2(new_n511_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n531_), .A2(new_n533_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n728_), .B1(new_n730_), .B2(new_n511_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n546_), .B2(new_n548_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n732_), .A2(new_n499_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n726_), .A2(KEYINPUT56), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n727_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT58), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n727_), .A2(new_n733_), .A3(KEYINPUT58), .A4(new_n734_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n737_), .A2(new_n572_), .A3(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n732_), .A2(new_n501_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n667_), .A2(KEYINPUT113), .A3(new_n499_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT113), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n743_), .B1(new_n549_), .B2(new_n498_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n725_), .A2(new_n497_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n486_), .A2(new_n490_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT115), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n746_), .A2(new_n747_), .A3(KEYINPUT55), .A4(new_n489_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n719_), .A2(KEYINPUT115), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n724_), .B1(new_n750_), .B2(new_n718_), .ZN(new_n751_));
  OAI21_X1  g550(.A(KEYINPUT117), .B1(new_n745_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT56), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT56), .ZN(new_n754_));
  OAI211_X1 g553(.A(KEYINPUT117), .B(new_n754_), .C1(new_n745_), .C2(new_n751_), .ZN(new_n755_));
  AOI22_X1  g554(.A1(new_n742_), .A2(new_n744_), .B1(new_n753_), .B2(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n741_), .B1(new_n756_), .B2(KEYINPUT118), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n742_), .A2(new_n744_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n753_), .A2(new_n755_), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n758_), .A2(KEYINPUT118), .A3(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n610_), .B1(new_n757_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT57), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n740_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n741_), .ZN(new_n764_));
  AOI21_X1  g563(.A(KEYINPUT113), .B1(new_n667_), .B2(new_n499_), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n549_), .A2(new_n743_), .A3(new_n498_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n754_), .B1(new_n726_), .B2(KEYINPUT117), .ZN(new_n767_));
  INV_X1    g566(.A(new_n755_), .ZN(new_n768_));
  OAI22_X1  g567(.A1(new_n765_), .A2(new_n766_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT118), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n764_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n758_), .A2(KEYINPUT118), .A3(new_n759_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n301_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT57), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n611_), .B1(new_n763_), .B2(new_n774_), .ZN(new_n775_));
  NOR4_X1   g574(.A1(new_n572_), .A2(new_n505_), .A3(new_n667_), .A4(new_n564_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT54), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n775_), .A2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n463_), .A2(new_n339_), .A3(new_n449_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(G113gat), .B1(new_n780_), .B2(new_n667_), .ZN(new_n781_));
  OAI21_X1  g580(.A(KEYINPUT59), .B1(new_n778_), .B2(new_n779_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT119), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n769_), .A2(new_n770_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n784_), .A2(new_n772_), .A3(new_n741_), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT57), .B1(new_n785_), .B2(new_n610_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n783_), .B1(new_n786_), .B2(new_n740_), .ZN(new_n787_));
  OAI211_X1 g586(.A(KEYINPUT119), .B(new_n739_), .C1(new_n773_), .C2(KEYINPUT57), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n774_), .A3(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n777_), .B1(new_n789_), .B2(new_n564_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n779_), .A2(KEYINPUT59), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n782_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(G113gat), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n667_), .B2(KEYINPUT120), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n796_), .B1(KEYINPUT120), .B2(new_n795_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n781_), .B1(new_n794_), .B2(new_n797_), .ZN(G1340gat));
  OAI211_X1 g597(.A(new_n782_), .B(new_n576_), .C1(new_n790_), .C2(new_n792_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(KEYINPUT121), .B(G120gat), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n800_), .B1(new_n669_), .B2(KEYINPUT60), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n780_), .B(new_n803_), .C1(KEYINPUT60), .C2(new_n800_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT122), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n802_), .A2(KEYINPUT122), .A3(new_n804_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(G1341gat));
  OAI21_X1  g608(.A(G127gat), .B1(new_n793_), .B2(new_n564_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n780_), .ZN(new_n811_));
  OR2_X1    g610(.A1(new_n564_), .A2(G127gat), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n810_), .B1(new_n811_), .B2(new_n812_), .ZN(G1342gat));
  OAI21_X1  g612(.A(G134gat), .B1(new_n793_), .B2(new_n620_), .ZN(new_n814_));
  OR2_X1    g613(.A1(new_n610_), .A2(G134gat), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n814_), .B1(new_n811_), .B2(new_n815_), .ZN(G1343gat));
  OR2_X1    g615(.A1(new_n775_), .A2(new_n777_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n384_), .A2(new_n338_), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n462_), .A2(new_n455_), .A3(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n667_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n576_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(G148gat), .ZN(G1345gat));
  OR3_X1    g624(.A1(new_n820_), .A2(KEYINPUT123), .A3(new_n564_), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT123), .B1(new_n820_), .B2(new_n564_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(KEYINPUT61), .B(G155gat), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n828_), .B(new_n829_), .ZN(G1346gat));
  OAI21_X1  g629(.A(G162gat), .B1(new_n820_), .B2(new_n620_), .ZN(new_n831_));
  OR2_X1    g630(.A1(new_n610_), .A2(G162gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n820_), .B2(new_n832_), .ZN(G1347gat));
  INV_X1    g632(.A(KEYINPUT125), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n462_), .A2(new_n464_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n835_), .A2(new_n384_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n834_), .B1(new_n790_), .B2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n761_), .A2(new_n762_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n739_), .B1(new_n773_), .B2(KEYINPUT57), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n839_), .B1(new_n840_), .B2(new_n783_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n611_), .B1(new_n841_), .B2(new_n788_), .ZN(new_n842_));
  OAI211_X1 g641(.A(KEYINPUT125), .B(new_n836_), .C1(new_n842_), .C2(new_n777_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n838_), .A2(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n845_));
  AND2_X1   g644(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n844_), .B(new_n667_), .C1(new_n845_), .C2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT124), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n774_), .B1(new_n763_), .B2(KEYINPUT119), .ZN(new_n849_));
  INV_X1    g648(.A(new_n788_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n564_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n777_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n853_), .A2(new_n667_), .A3(new_n836_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT62), .ZN(new_n855_));
  AND4_X1   g654(.A1(new_n848_), .A2(new_n854_), .A3(new_n855_), .A4(G169gat), .ZN(new_n856_));
  INV_X1    g655(.A(G169gat), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n857_), .B1(KEYINPUT124), .B2(KEYINPUT62), .ZN(new_n858_));
  AOI22_X1  g657(.A1(new_n854_), .A2(new_n858_), .B1(new_n848_), .B2(new_n855_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n847_), .B1(new_n856_), .B2(new_n859_), .ZN(G1348gat));
  AOI21_X1  g659(.A(G176gat), .B1(new_n844_), .B2(new_n505_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n778_), .A2(new_n384_), .ZN(new_n862_));
  INV_X1    g661(.A(G176gat), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n575_), .A2(new_n863_), .A3(new_n835_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n861_), .B1(new_n862_), .B2(new_n864_), .ZN(G1349gat));
  NOR2_X1   g664(.A1(new_n835_), .A2(new_n564_), .ZN(new_n866_));
  AOI21_X1  g665(.A(G183gat), .B1(new_n862_), .B2(new_n866_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n564_), .A2(new_n302_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n844_), .B2(new_n868_), .ZN(G1350gat));
  NAND3_X1  g668(.A1(new_n844_), .A2(new_n303_), .A3(new_n301_), .ZN(new_n870_));
  AOI21_X1  g669(.A(KEYINPUT125), .B1(new_n853_), .B2(new_n836_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n790_), .A2(new_n834_), .A3(new_n837_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n572_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(KEYINPUT126), .B1(new_n873_), .B2(G190gat), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n620_), .B1(new_n838_), .B2(new_n843_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT126), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n875_), .A2(new_n876_), .A3(new_n307_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n870_), .B1(new_n874_), .B2(new_n877_), .ZN(G1351gat));
  XOR2_X1   g677(.A(KEYINPUT127), .B(G197gat), .Z(new_n879_));
  NOR2_X1   g678(.A1(KEYINPUT127), .A2(G197gat), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n593_), .A2(new_n449_), .A3(new_n818_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n817_), .A2(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n549_), .ZN(new_n883_));
  MUX2_X1   g682(.A(new_n879_), .B(new_n880_), .S(new_n883_), .Z(G1352gat));
  NOR2_X1   g683(.A1(new_n882_), .A2(new_n575_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(new_n357_), .ZN(G1353gat));
  NAND3_X1  g685(.A1(new_n817_), .A2(new_n611_), .A3(new_n881_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n888_));
  AND2_X1   g687(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n887_), .A2(new_n888_), .A3(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n890_), .B1(new_n887_), .B2(new_n888_), .ZN(G1354gat));
  OAI21_X1  g690(.A(G218gat), .B1(new_n882_), .B2(new_n620_), .ZN(new_n892_));
  OR2_X1    g691(.A1(new_n610_), .A2(G218gat), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n882_), .B2(new_n893_), .ZN(G1355gat));
endmodule


