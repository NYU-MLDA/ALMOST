//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 0 1 0 0 0 1 0 1 1 1 1 1 1 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 1 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n854_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n863_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G232gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT34), .ZN(new_n204_));
  AND2_X1   g003(.A1(new_n204_), .A2(KEYINPUT35), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(KEYINPUT35), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(G29gat), .B(G36gat), .Z(new_n209_));
  XOR2_X1   g008(.A(G43gat), .B(G50gat), .Z(new_n210_));
  XOR2_X1   g009(.A(new_n209_), .B(new_n210_), .Z(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT15), .ZN(new_n212_));
  XOR2_X1   g011(.A(G85gat), .B(G92gat), .Z(new_n213_));
  NOR2_X1   g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT7), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G99gat), .A2(G106gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT6), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n213_), .B1(new_n216_), .B2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT8), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT10), .B(G99gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(KEYINPUT64), .ZN(new_n223_));
  INV_X1    g022(.A(G106gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n219_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n213_), .A2(KEYINPUT9), .ZN(new_n227_));
  INV_X1    g026(.A(G85gat), .ZN(new_n228_));
  INV_X1    g027(.A(G92gat), .ZN(new_n229_));
  OR3_X1    g028(.A1(new_n228_), .A2(new_n229_), .A3(KEYINPUT9), .ZN(new_n230_));
  AND3_X1   g029(.A1(new_n226_), .A2(new_n227_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n225_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n221_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n212_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n221_), .A2(new_n211_), .A3(new_n232_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n208_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT15), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n211_), .B(new_n237_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n220_), .A2(KEYINPUT8), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n220_), .A2(KEYINPUT8), .ZN(new_n240_));
  AOI22_X1  g039(.A1(new_n239_), .A2(new_n240_), .B1(new_n225_), .B2(new_n231_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n235_), .B(new_n205_), .C1(new_n238_), .C2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT67), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n234_), .A2(new_n244_), .A3(new_n205_), .A4(new_n235_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n236_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G190gat), .B(G218gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G134gat), .B(G162gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n249_), .A2(KEYINPUT36), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n246_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n246_), .A2(KEYINPUT68), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n249_), .B(KEYINPUT36), .Z(new_n254_));
  OAI21_X1  g053(.A(new_n254_), .B1(new_n246_), .B2(KEYINPUT68), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n202_), .B(new_n251_), .C1(new_n253_), .C2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n254_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n251_), .B1(new_n246_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT37), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n256_), .A2(new_n259_), .A3(KEYINPUT69), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n246_), .A2(KEYINPUT68), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n262_), .A2(new_n263_), .A3(new_n202_), .A4(new_n251_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n260_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n265_), .B1(new_n260_), .B2(new_n264_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G230gat), .A2(G233gat), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G57gat), .B(G64gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT11), .ZN(new_n272_));
  XOR2_X1   g071(.A(G71gat), .B(G78gat), .Z(new_n273_));
  OR2_X1    g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n271_), .A2(KEYINPUT11), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n272_), .A2(new_n273_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n274_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n233_), .A2(new_n278_), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n279_), .A2(KEYINPUT12), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n241_), .A2(new_n277_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(new_n281_), .A3(KEYINPUT12), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n270_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n269_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G176gat), .B(G204gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT66), .ZN(new_n287_));
  XOR2_X1   g086(.A(KEYINPUT65), .B(KEYINPUT5), .Z(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G120gat), .B(G148gat), .ZN(new_n290_));
  XOR2_X1   g089(.A(new_n289_), .B(new_n290_), .Z(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n285_), .A2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n291_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT13), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n293_), .A2(KEYINPUT13), .A3(new_n294_), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  AND2_X1   g098(.A1(G231gat), .A2(G233gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n277_), .B(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G15gat), .B(G22gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT71), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT14), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n306_), .B1(G1gat), .B2(G8gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT72), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n305_), .A2(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(G1gat), .B(G8gat), .Z(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n303_), .B(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G127gat), .B(G155gat), .Z(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT16), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G183gat), .B(G211gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT17), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n317_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n312_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n320_), .A2(KEYINPUT74), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n320_), .B(KEYINPUT74), .C1(new_n318_), .C2(new_n312_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n268_), .A2(new_n299_), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(G8gat), .B(G36gat), .Z(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G64gat), .B(G92gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G226gat), .A2(G233gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT19), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT93), .B(KEYINPUT20), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G183gat), .A2(G190gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT23), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT23), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n337_), .A2(G183gat), .A3(G190gat), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT24), .ZN(new_n339_));
  NOR2_X1   g138(.A1(G169gat), .A2(G176gat), .ZN(new_n340_));
  AOI22_X1  g139(.A1(new_n336_), .A2(new_n338_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(G169gat), .ZN(new_n342_));
  INV_X1    g141(.A(G176gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G169gat), .A2(G176gat), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n344_), .A2(KEYINPUT24), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(G190gat), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT77), .B1(new_n347_), .B2(KEYINPUT26), .ZN(new_n348_));
  INV_X1    g147(.A(G183gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT25), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT25), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(G183gat), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n348_), .A2(new_n350_), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT26), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(G190gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n347_), .A2(KEYINPUT26), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT77), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n341_), .B(new_n346_), .C1(new_n353_), .C2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n335_), .A2(new_n337_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n359_), .B(new_n360_), .C1(G183gat), .C2(G190gat), .ZN(new_n361_));
  OAI21_X1  g160(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n362_));
  OR3_X1    g161(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n361_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n358_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT78), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n358_), .A2(new_n367_), .A3(new_n364_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G211gat), .B(G218gat), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT21), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(G197gat), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT83), .B1(new_n373_), .B2(G204gat), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT83), .ZN(new_n375_));
  INV_X1    g174(.A(G204gat), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(new_n376_), .A3(G197gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n373_), .A2(G204gat), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n374_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n372_), .A2(new_n379_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n374_), .A2(new_n377_), .A3(new_n371_), .A4(new_n378_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G197gat), .B(G204gat), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n370_), .B1(new_n383_), .B2(new_n371_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT84), .ZN(new_n385_));
  NOR3_X1   g184(.A1(new_n382_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(G218gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(G211gat), .ZN(new_n388_));
  INV_X1    g187(.A(G211gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(G218gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n376_), .A2(G197gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n378_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n391_), .B1(KEYINPUT21), .B2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(KEYINPUT84), .B1(new_n394_), .B2(new_n381_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n380_), .B1(new_n386_), .B2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n334_), .B1(new_n369_), .B2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n385_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n394_), .A2(KEYINPUT84), .A3(new_n381_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT22), .B(G169gat), .ZN(new_n401_));
  AND2_X1   g200(.A1(new_n401_), .A2(KEYINPUT88), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n401_), .A2(KEYINPUT88), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n343_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n361_), .A2(new_n345_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n355_), .A2(new_n356_), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n350_), .A2(new_n352_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n409_), .A2(new_n346_), .A3(new_n341_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n400_), .A2(new_n406_), .A3(new_n380_), .A4(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n333_), .B1(new_n397_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n336_), .A2(new_n338_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n340_), .A2(new_n339_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n346_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  AND4_X1   g214(.A1(new_n355_), .A2(new_n356_), .A3(new_n350_), .A4(new_n352_), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT87), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT87), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n409_), .A2(new_n341_), .A3(new_n418_), .A4(new_n346_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n406_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n396_), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n398_), .A2(new_n399_), .B1(new_n379_), .B2(new_n372_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n423_), .A2(new_n366_), .A3(new_n368_), .ZN(new_n424_));
  AND4_X1   g223(.A1(KEYINPUT20), .A2(new_n422_), .A3(new_n424_), .A4(new_n333_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT94), .B1(new_n412_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n334_), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n358_), .A2(new_n367_), .A3(new_n364_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n367_), .B1(new_n358_), .B2(new_n364_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n411_), .B(new_n427_), .C1(new_n430_), .C2(new_n423_), .ZN(new_n431_));
  AOI21_X1  g230(.A(KEYINPUT94), .B1(new_n431_), .B2(new_n332_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n330_), .B1(new_n426_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT20), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n435_), .B1(new_n421_), .B2(new_n396_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n424_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(new_n332_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n332_), .A2(new_n435_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n440_), .B1(new_n369_), .B2(new_n396_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n423_), .A2(new_n406_), .A3(new_n420_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n438_), .A2(new_n330_), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT27), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT95), .B1(new_n434_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n330_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT94), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n431_), .A2(new_n332_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n436_), .A2(new_n333_), .A3(new_n424_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n448_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n447_), .B1(new_n451_), .B2(new_n432_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT95), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT27), .ZN(new_n454_));
  AOI22_X1  g253(.A1(new_n437_), .A2(new_n332_), .B1(new_n442_), .B2(new_n441_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n454_), .B1(new_n455_), .B2(new_n330_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n452_), .A2(new_n453_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n446_), .A2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT86), .B(G106gat), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT29), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT82), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  OAI211_X1 g262(.A(KEYINPUT82), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G141gat), .A2(G148gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT80), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT80), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(G141gat), .A3(G148gat), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT2), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n467_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  NOR3_X1   g270(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n472_));
  AND3_X1   g271(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n465_), .A2(new_n471_), .A3(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT81), .B1(G155gat), .B2(G162gat), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NOR3_X1   g276(.A1(KEYINPUT81), .A2(G155gat), .A3(G162gat), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(G155gat), .ZN(new_n480_));
  INV_X1    g279(.A(G162gat), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n479_), .A2(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT1), .B1(new_n480_), .B2(new_n481_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT1), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n485_), .A2(G155gat), .A3(G162gat), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n484_), .B(new_n486_), .C1(new_n477_), .C2(new_n478_), .ZN(new_n487_));
  OR2_X1    g286(.A1(G141gat), .A2(G148gat), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n467_), .A2(new_n469_), .A3(new_n488_), .ZN(new_n489_));
  AOI22_X1  g288(.A1(new_n475_), .A2(new_n483_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n396_), .B1(new_n460_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(G78gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G22gat), .B(G50gat), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT28), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n490_), .A2(new_n495_), .A3(new_n460_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n495_), .B1(new_n490_), .B2(new_n460_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n494_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G228gat), .A2(G233gat), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT85), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n499_), .B1(new_n396_), .B2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n475_), .A2(new_n483_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n487_), .A2(new_n489_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT28), .B1(new_n504_), .B2(KEYINPUT29), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n490_), .A2(new_n495_), .A3(new_n460_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n494_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n498_), .A2(new_n501_), .A3(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n501_), .B1(new_n498_), .B2(new_n508_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n493_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n501_), .ZN(new_n512_));
  NOR3_X1   g311(.A1(new_n496_), .A2(new_n497_), .A3(new_n494_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n507_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n512_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n491_), .B(G78gat), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n498_), .A2(new_n501_), .A3(new_n508_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n515_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n459_), .B1(new_n511_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n511_), .A2(new_n518_), .A3(new_n459_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n441_), .A2(new_n442_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n333_), .B1(new_n436_), .B2(new_n424_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n447_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n525_), .A2(new_n444_), .A3(KEYINPUT90), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT90), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n455_), .A2(new_n527_), .A3(new_n330_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n526_), .A2(new_n454_), .A3(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n458_), .A2(new_n522_), .A3(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(G127gat), .B(G134gat), .Z(new_n531_));
  XOR2_X1   g330(.A(G113gat), .B(G120gat), .Z(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n533_), .B(KEYINPUT31), .Z(new_n534_));
  XNOR2_X1  g333(.A(G71gat), .B(G99gat), .ZN(new_n535_));
  INV_X1    g334(.A(G43gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n369_), .B(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G227gat), .A2(G233gat), .ZN(new_n539_));
  INV_X1    g338(.A(G15gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT30), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n538_), .B(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n534_), .B1(new_n543_), .B2(KEYINPUT79), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n544_), .B1(KEYINPUT79), .B2(new_n543_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n543_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT79), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n546_), .A2(new_n547_), .A3(new_n534_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n545_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G225gat), .A2(G233gat), .ZN(new_n550_));
  INV_X1    g349(.A(new_n533_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n504_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n490_), .A2(new_n533_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n552_), .A2(KEYINPUT4), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT4), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n504_), .A2(new_n555_), .A3(new_n551_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n550_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G1gat), .B(G29gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G57gat), .B(G85gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT91), .B(KEYINPUT0), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n550_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n564_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n565_));
  OR3_X1    g364(.A1(new_n557_), .A2(new_n563_), .A3(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n563_), .B1(new_n557_), .B2(new_n565_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NOR3_X1   g367(.A1(new_n530_), .A2(new_n549_), .A3(new_n568_), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n452_), .A2(new_n453_), .A3(new_n456_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n453_), .B1(new_n452_), .B2(new_n456_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n529_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n568_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n520_), .A2(new_n573_), .A3(new_n521_), .ZN(new_n574_));
  OAI21_X1  g373(.A(KEYINPUT96), .B1(new_n572_), .B2(new_n574_), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n511_), .A2(new_n459_), .A3(new_n518_), .ZN(new_n576_));
  NOR3_X1   g375(.A1(new_n576_), .A2(new_n519_), .A3(new_n568_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT96), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n458_), .A2(new_n577_), .A3(new_n578_), .A4(new_n529_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n526_), .A2(new_n528_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n552_), .A2(new_n564_), .A3(new_n553_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n562_), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n582_), .A2(KEYINPUT92), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(KEYINPUT92), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n554_), .A2(new_n550_), .A3(new_n556_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n583_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT33), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n567_), .A2(new_n587_), .ZN(new_n588_));
  OAI211_X1 g387(.A(KEYINPUT33), .B(new_n563_), .C1(new_n557_), .C2(new_n565_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n586_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n580_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n330_), .A2(KEYINPUT32), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n455_), .A2(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n451_), .A2(new_n432_), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n568_), .B(new_n593_), .C1(new_n594_), .C2(new_n592_), .ZN(new_n595_));
  AOI22_X1  g394(.A1(new_n591_), .A2(new_n595_), .B1(new_n521_), .B2(new_n520_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n575_), .A2(new_n579_), .A3(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n569_), .B1(new_n598_), .B2(new_n549_), .ZN(new_n599_));
  XOR2_X1   g398(.A(G113gat), .B(G141gat), .Z(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT75), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G169gat), .B(G197gat), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n601_), .B(new_n602_), .Z(new_n603_));
  INV_X1    g402(.A(new_n211_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n311_), .B(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(G229gat), .A2(G233gat), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n212_), .A2(new_n311_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n311_), .A2(new_n604_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n609_), .A2(new_n610_), .A3(new_n606_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n603_), .B1(new_n608_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT76), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n608_), .A2(new_n611_), .A3(new_n603_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n613_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n614_), .B1(new_n613_), .B2(new_n615_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n599_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n325_), .A2(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n568_), .A2(KEYINPUT97), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n568_), .A2(KEYINPUT97), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n621_), .A2(G1gat), .A3(new_n625_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT98), .Z(new_n627_));
  INV_X1    g426(.A(KEYINPUT38), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n628_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n262_), .A2(new_n251_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n599_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n299_), .A2(new_n618_), .A3(new_n323_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT99), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(G1gat), .B1(new_n636_), .B2(new_n573_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n629_), .A2(new_n630_), .A3(new_n637_), .ZN(G1324gat));
  INV_X1    g437(.A(new_n572_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n636_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT100), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(KEYINPUT100), .B1(new_n636_), .B2(new_n639_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n642_), .A2(G8gat), .A3(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT39), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT101), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT102), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n647_), .B1(new_n644_), .B2(KEYINPUT39), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT101), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n644_), .A2(new_n649_), .A3(KEYINPUT39), .ZN(new_n650_));
  INV_X1    g449(.A(G8gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT39), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n652_), .A2(KEYINPUT102), .A3(new_n653_), .A4(new_n643_), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n646_), .A2(new_n648_), .A3(new_n650_), .A4(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n621_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n656_), .A2(new_n651_), .A3(new_n572_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT40), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n655_), .A2(KEYINPUT40), .A3(new_n657_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(G1325gat));
  OAI21_X1  g461(.A(G15gat), .B1(new_n636_), .B2(new_n549_), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT41), .Z(new_n664_));
  INV_X1    g463(.A(new_n549_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n656_), .A2(new_n540_), .A3(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(G1326gat));
  OAI21_X1  g466(.A(G22gat), .B1(new_n636_), .B2(new_n522_), .ZN(new_n668_));
  XOR2_X1   g467(.A(new_n668_), .B(KEYINPUT42), .Z(new_n669_));
  NOR3_X1   g468(.A1(new_n621_), .A2(G22gat), .A3(new_n522_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT103), .ZN(G1327gat));
  NOR2_X1   g471(.A1(new_n323_), .A2(new_n631_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n673_), .A2(new_n299_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n620_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(G29gat), .B1(new_n676_), .B2(new_n568_), .ZN(new_n677_));
  OAI21_X1  g476(.A(KEYINPUT43), .B1(new_n599_), .B2(new_n268_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n260_), .A2(new_n264_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT70), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n260_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n458_), .A2(new_n577_), .A3(new_n529_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n596_), .B1(new_n684_), .B2(KEYINPUT96), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n665_), .B1(new_n685_), .B2(new_n579_), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n679_), .B(new_n683_), .C1(new_n686_), .C2(new_n569_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n678_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n323_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(new_n299_), .A3(new_n618_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(KEYINPUT44), .B1(new_n688_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693_));
  AOI211_X1 g492(.A(new_n693_), .B(new_n690_), .C1(new_n678_), .C2(new_n687_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n692_), .A2(new_n694_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n624_), .A2(G29gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n677_), .B1(new_n695_), .B2(new_n696_), .ZN(G1328gat));
  NOR3_X1   g496(.A1(new_n675_), .A2(G36gat), .A3(new_n639_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n698_), .B(new_n699_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n692_), .A2(new_n694_), .A3(new_n639_), .ZN(new_n701_));
  INV_X1    g500(.A(G36gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n700_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT46), .Z(G1329gat));
  OAI21_X1  g503(.A(new_n536_), .B1(new_n675_), .B2(new_n549_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT106), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n549_), .A2(new_n536_), .ZN(new_n707_));
  AOI21_X1  g506(.A(KEYINPUT105), .B1(new_n695_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT105), .ZN(new_n709_));
  INV_X1    g508(.A(new_n707_), .ZN(new_n710_));
  NOR4_X1   g509(.A1(new_n692_), .A2(new_n694_), .A3(new_n709_), .A4(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n706_), .B1(new_n708_), .B2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT108), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT108), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n714_), .B(new_n706_), .C1(new_n708_), .C2(new_n711_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n713_), .A2(new_n715_), .A3(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n713_), .B2(new_n715_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1330gat));
  INV_X1    g518(.A(new_n522_), .ZN(new_n720_));
  AOI21_X1  g519(.A(G50gat), .B1(new_n676_), .B2(new_n720_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n720_), .A2(G50gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n695_), .B2(new_n722_), .ZN(G1331gat));
  NOR2_X1   g522(.A1(new_n299_), .A2(new_n618_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n599_), .A2(new_n725_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n683_), .A2(new_n689_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT109), .ZN(new_n729_));
  AOI21_X1  g528(.A(G57gat), .B1(new_n729_), .B2(new_n624_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT110), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n730_), .A2(new_n731_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n725_), .A2(new_n689_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n633_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n736_), .A2(G57gat), .A3(new_n568_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT111), .Z(new_n738_));
  NOR3_X1   g537(.A1(new_n732_), .A2(new_n733_), .A3(new_n738_), .ZN(G1332gat));
  OAI21_X1  g538(.A(G64gat), .B1(new_n735_), .B2(new_n639_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT48), .ZN(new_n741_));
  INV_X1    g540(.A(G64gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n729_), .A2(new_n742_), .A3(new_n572_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1333gat));
  OAI21_X1  g543(.A(G71gat), .B1(new_n735_), .B2(new_n549_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT49), .ZN(new_n746_));
  INV_X1    g545(.A(G71gat), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n729_), .A2(new_n747_), .A3(new_n665_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(G1334gat));
  OAI21_X1  g548(.A(G78gat), .B1(new_n735_), .B2(new_n522_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT112), .Z(new_n751_));
  OR2_X1    g550(.A1(new_n751_), .A2(KEYINPUT50), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(KEYINPUT50), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n729_), .A2(new_n492_), .A3(new_n720_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n752_), .A2(new_n753_), .A3(new_n754_), .ZN(G1335gat));
  INV_X1    g554(.A(new_n688_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n725_), .A2(new_n323_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n756_), .A2(new_n573_), .A3(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n726_), .A2(new_n673_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n624_), .A2(new_n228_), .ZN(new_n761_));
  OAI22_X1  g560(.A1(new_n759_), .A2(new_n228_), .B1(new_n760_), .B2(new_n761_), .ZN(G1336gat));
  OAI21_X1  g561(.A(new_n229_), .B1(new_n760_), .B2(new_n639_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT113), .Z(new_n764_));
  NOR2_X1   g563(.A1(new_n756_), .A2(new_n758_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n639_), .A2(new_n229_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n764_), .B1(new_n765_), .B2(new_n766_), .ZN(G1337gat));
  NOR3_X1   g566(.A1(new_n756_), .A2(new_n549_), .A3(new_n758_), .ZN(new_n768_));
  INV_X1    g567(.A(G99gat), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n665_), .A2(new_n223_), .ZN(new_n770_));
  OAI22_X1  g569(.A1(new_n768_), .A2(new_n769_), .B1(new_n760_), .B2(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT51), .ZN(G1338gat));
  NOR3_X1   g571(.A1(new_n756_), .A2(new_n522_), .A3(new_n758_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n774_));
  OR3_X1    g573(.A1(new_n773_), .A2(new_n774_), .A3(new_n224_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n773_), .B2(new_n224_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(KEYINPUT52), .A3(new_n776_), .ZN(new_n777_));
  OR2_X1    g576(.A1(new_n776_), .A2(KEYINPUT52), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n726_), .A2(new_n224_), .A3(new_n720_), .A4(new_n673_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n777_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g580(.A(KEYINPUT57), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n603_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n609_), .A2(new_n610_), .A3(new_n607_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n615_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n786_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n293_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT56), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n283_), .A2(KEYINPUT55), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n283_), .A2(KEYINPUT55), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n280_), .A2(new_n270_), .A3(new_n282_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT116), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n280_), .A2(new_n794_), .A3(new_n270_), .A4(new_n282_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n790_), .A2(new_n791_), .A3(new_n793_), .A4(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n789_), .B1(new_n796_), .B2(new_n291_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT117), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n788_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n796_), .A2(new_n291_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT56), .B1(new_n800_), .B2(new_n798_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n787_), .B1(new_n799_), .B2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n782_), .B1(new_n803_), .B2(new_n632_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n787_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n800_), .A2(new_n798_), .A3(KEYINPUT56), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(new_n618_), .A3(new_n293_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n805_), .B1(new_n807_), .B2(new_n801_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n808_), .A2(KEYINPUT57), .A3(new_n631_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT58), .ZN(new_n810_));
  INV_X1    g609(.A(new_n797_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n786_), .B1(new_n285_), .B2(new_n292_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n800_), .A2(KEYINPUT56), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n810_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n814_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n816_), .A2(KEYINPUT58), .A3(new_n811_), .A4(new_n812_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n815_), .A2(new_n683_), .A3(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n804_), .A2(new_n809_), .A3(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n689_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT120), .ZN(new_n821_));
  XNOR2_X1  g620(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n324_), .B2(new_n618_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n727_), .A2(new_n619_), .A3(new_n299_), .A4(new_n822_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT120), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n819_), .A2(new_n827_), .A3(new_n689_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n821_), .A2(new_n826_), .A3(new_n828_), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n530_), .A2(new_n549_), .A3(new_n625_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(KEYINPUT118), .ZN(new_n831_));
  XOR2_X1   g630(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n832_));
  AND3_X1   g631(.A1(new_n829_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n820_), .A2(new_n826_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n831_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n835_), .A2(KEYINPUT59), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n833_), .A2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(G113gat), .B1(new_n837_), .B2(new_n619_), .ZN(new_n838_));
  OR3_X1    g637(.A1(new_n835_), .A2(G113gat), .A3(new_n619_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(G1340gat));
  OAI21_X1  g639(.A(G120gat), .B1(new_n837_), .B2(new_n299_), .ZN(new_n841_));
  INV_X1    g640(.A(G120gat), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(new_n299_), .B2(KEYINPUT60), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n843_), .B1(KEYINPUT60), .B2(new_n842_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n841_), .B1(new_n835_), .B2(new_n844_), .ZN(G1341gat));
  INV_X1    g644(.A(new_n835_), .ZN(new_n846_));
  AOI21_X1  g645(.A(G127gat), .B1(new_n846_), .B2(new_n323_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(KEYINPUT121), .ZN(new_n848_));
  INV_X1    g647(.A(new_n837_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n323_), .A2(G127gat), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n848_), .B1(new_n849_), .B2(new_n850_), .ZN(G1342gat));
  AOI21_X1  g650(.A(G134gat), .B1(new_n846_), .B2(new_n632_), .ZN(new_n852_));
  XOR2_X1   g651(.A(KEYINPUT122), .B(G134gat), .Z(new_n853_));
  NOR2_X1   g652(.A1(new_n268_), .A2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n852_), .B1(new_n849_), .B2(new_n854_), .ZN(G1343gat));
  AOI21_X1  g654(.A(new_n665_), .B1(new_n820_), .B2(new_n826_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n625_), .A2(new_n572_), .A3(new_n522_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n618_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g660(.A(new_n299_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n859_), .A2(new_n862_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G148gat), .ZN(G1345gat));
  OR3_X1    g663(.A1(new_n858_), .A2(KEYINPUT123), .A3(new_n689_), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT123), .B1(new_n858_), .B2(new_n689_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT61), .B(G155gat), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(G1346gat));
  OAI21_X1  g668(.A(G162gat), .B1(new_n858_), .B2(new_n268_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n632_), .A2(new_n481_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n858_), .B2(new_n871_), .ZN(G1347gat));
  INV_X1    g671(.A(new_n828_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n827_), .B1(new_n819_), .B2(new_n689_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n824_), .A2(new_n825_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n873_), .A2(new_n874_), .A3(new_n875_), .ZN(new_n876_));
  NOR4_X1   g675(.A1(new_n639_), .A2(new_n549_), .A3(new_n720_), .A4(new_n624_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(KEYINPUT124), .B1(new_n876_), .B2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT124), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n829_), .A2(new_n880_), .A3(new_n877_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n618_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(KEYINPUT125), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n882_), .A2(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n829_), .A2(new_n618_), .A3(new_n877_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT62), .ZN(new_n887_));
  AND3_X1   g686(.A1(new_n886_), .A2(new_n887_), .A3(G169gat), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n886_), .B2(G169gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n885_), .B1(new_n888_), .B2(new_n889_), .ZN(G1348gat));
  AOI21_X1  g689(.A(new_n878_), .B1(new_n820_), .B2(new_n826_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n891_), .A2(G176gat), .A3(new_n862_), .ZN(new_n892_));
  XOR2_X1   g691(.A(new_n892_), .B(KEYINPUT126), .Z(new_n893_));
  NAND2_X1  g692(.A1(new_n882_), .A2(new_n862_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n893_), .B1(new_n894_), .B2(new_n343_), .ZN(G1349gat));
  AOI21_X1  g694(.A(G183gat), .B1(new_n891_), .B2(new_n323_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n689_), .A2(new_n408_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n896_), .B1(new_n882_), .B2(new_n897_), .ZN(G1350gat));
  NAND3_X1  g697(.A1(new_n882_), .A2(new_n407_), .A3(new_n632_), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n829_), .A2(new_n880_), .A3(new_n877_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n880_), .B1(new_n829_), .B2(new_n877_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n683_), .B1(new_n900_), .B2(new_n901_), .ZN(new_n902_));
  AND3_X1   g701(.A1(new_n902_), .A2(KEYINPUT127), .A3(G190gat), .ZN(new_n903_));
  AOI21_X1  g702(.A(KEYINPUT127), .B1(new_n902_), .B2(G190gat), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n899_), .B1(new_n903_), .B2(new_n904_), .ZN(G1351gat));
  NOR2_X1   g704(.A1(new_n639_), .A2(new_n574_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n856_), .A2(new_n906_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(new_n619_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(new_n373_), .ZN(G1352gat));
  NOR2_X1   g708(.A1(new_n907_), .A2(new_n299_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(new_n376_), .ZN(G1353gat));
  NAND3_X1  g710(.A1(new_n856_), .A2(new_n323_), .A3(new_n906_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n913_));
  AND2_X1   g712(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n912_), .A2(new_n913_), .A3(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n915_), .B1(new_n912_), .B2(new_n913_), .ZN(G1354gat));
  OAI21_X1  g715(.A(G218gat), .B1(new_n907_), .B2(new_n268_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n632_), .A2(new_n387_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n907_), .B2(new_n918_), .ZN(G1355gat));
endmodule


