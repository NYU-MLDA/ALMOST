//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 1 1 1 0 0 0 1 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n915_, new_n917_, new_n918_, new_n920_,
    new_n921_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_, new_n938_, new_n939_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n954_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_;
  XOR2_X1   g000(.A(G190gat), .B(G218gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT36), .ZN(new_n205_));
  AND3_X1   g004(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n206_));
  AOI21_X1  g005(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT10), .B(G99gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n208_), .B1(G106gat), .B2(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G92gat), .Z(new_n211_));
  INV_X1    g010(.A(KEYINPUT9), .ZN(new_n212_));
  AND2_X1   g011(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n212_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G85gat), .ZN(new_n216_));
  INV_X1    g015(.A(G92gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  OAI22_X1  g017(.A1(new_n211_), .A2(new_n215_), .B1(new_n212_), .B2(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G85gat), .A2(G92gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n210_), .B1(new_n219_), .B2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NOR3_X1   g023(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT68), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT7), .ZN(new_n227_));
  INV_X1    g026(.A(G99gat), .ZN(new_n228_));
  INV_X1    g027(.A(G106gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT68), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n230_), .A2(new_n231_), .A3(new_n223_), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT67), .B1(new_n206_), .B2(new_n207_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G99gat), .A2(G106gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT6), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n237_));
  NAND3_X1  g036(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  AOI22_X1  g038(.A1(new_n226_), .A2(new_n232_), .B1(new_n233_), .B2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G85gat), .B(G92gat), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT8), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n230_), .A2(new_n236_), .A3(new_n238_), .A4(new_n223_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n208_), .A2(KEYINPUT66), .A3(new_n230_), .A4(new_n223_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n241_), .A2(KEYINPUT8), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n222_), .B1(new_n242_), .B2(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(G43gat), .B(G50gat), .Z(new_n250_));
  INV_X1    g049(.A(G36gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(G29gat), .ZN(new_n252_));
  INV_X1    g051(.A(G29gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(G36gat), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n252_), .A2(new_n254_), .A3(KEYINPUT77), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT77), .B1(new_n252_), .B2(new_n254_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n250_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT77), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n253_), .A2(G36gat), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n251_), .A2(G29gat), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n258_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n252_), .A2(new_n254_), .A3(KEYINPUT77), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G43gat), .B(G50gat), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n261_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n257_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT35), .ZN(new_n266_));
  XOR2_X1   g065(.A(KEYINPUT75), .B(KEYINPUT34), .Z(new_n267_));
  NAND2_X1  g066(.A1(G232gat), .A2(G233gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  AOI22_X1  g068(.A1(new_n249_), .A2(new_n265_), .B1(new_n266_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT8), .ZN(new_n272_));
  AND3_X1   g071(.A1(new_n230_), .A2(new_n231_), .A3(new_n223_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n231_), .B1(new_n230_), .B2(new_n223_), .ZN(new_n274_));
  NOR3_X1   g073(.A1(new_n206_), .A2(new_n207_), .A3(KEYINPUT67), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n237_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n276_));
  OAI22_X1  g075(.A1(new_n273_), .A2(new_n274_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n241_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n272_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n271_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n242_), .A2(KEYINPUT70), .A3(new_n248_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n222_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NOR3_X1   g082(.A1(new_n255_), .A2(new_n256_), .A3(new_n250_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n263_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n285_));
  NOR3_X1   g084(.A1(new_n284_), .A2(new_n285_), .A3(KEYINPUT15), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT15), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n287_), .B1(new_n257_), .B2(new_n264_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n270_), .B1(new_n283_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT76), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n269_), .A2(new_n266_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT76), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n293_), .B(new_n270_), .C1(new_n283_), .C2(new_n289_), .ZN(new_n294_));
  AND3_X1   g093(.A1(new_n291_), .A2(new_n292_), .A3(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n292_), .B1(new_n291_), .B2(new_n294_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n205_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT80), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  OAI211_X1 g098(.A(KEYINPUT80), .B(new_n205_), .C1(new_n295_), .C2(new_n296_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n292_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n222_), .ZN(new_n302_));
  NOR3_X1   g101(.A1(new_n279_), .A2(new_n271_), .A3(new_n280_), .ZN(new_n303_));
  AOI21_X1  g102(.A(KEYINPUT70), .B1(new_n242_), .B2(new_n248_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n302_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n289_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n293_), .B1(new_n307_), .B2(new_n270_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n294_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n301_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n291_), .A2(new_n292_), .A3(new_n294_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT36), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n204_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT78), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n310_), .A2(new_n311_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT79), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n310_), .A2(KEYINPUT79), .A3(new_n311_), .A4(new_n314_), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n299_), .A2(new_n300_), .A3(new_n317_), .A4(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT37), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT37), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n297_), .A2(new_n321_), .A3(new_n315_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G15gat), .B(G22gat), .ZN(new_n324_));
  INV_X1    g123(.A(G1gat), .ZN(new_n325_));
  INV_X1    g124(.A(G8gat), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT14), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n324_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G1gat), .B(G8gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G231gat), .A2(G233gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(G71gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT69), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT69), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(G71gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(G78gat), .ZN(new_n338_));
  INV_X1    g137(.A(G78gat), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n334_), .A2(new_n336_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(G64gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(G57gat), .ZN(new_n342_));
  INV_X1    g141(.A(G57gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(G64gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n342_), .A2(new_n344_), .A3(KEYINPUT11), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(KEYINPUT11), .B1(new_n342_), .B2(new_n344_), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n338_), .B(new_n340_), .C1(new_n346_), .C2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n340_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n339_), .B1(new_n334_), .B2(new_n336_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n345_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n348_), .A2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n332_), .B(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G127gat), .B(G155gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT16), .ZN(new_n355_));
  XOR2_X1   g154(.A(G183gat), .B(G211gat), .Z(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n353_), .B1(KEYINPUT17), .B2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n358_), .A2(KEYINPUT81), .A3(KEYINPUT17), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n323_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT82), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT73), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT72), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n348_), .A2(new_n351_), .ZN(new_n366_));
  AOI211_X1 g165(.A(new_n222_), .B(new_n366_), .C1(new_n242_), .C2(new_n248_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G230gat), .A2(G233gat), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n365_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n302_), .B(new_n352_), .C1(new_n279_), .C2(new_n280_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n371_), .A2(KEYINPUT72), .A3(new_n368_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  XOR2_X1   g172(.A(KEYINPUT71), .B(KEYINPUT12), .Z(new_n374_));
  OAI21_X1  g173(.A(new_n374_), .B1(new_n249_), .B2(new_n352_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n366_), .A2(KEYINPUT12), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n375_), .B1(new_n283_), .B2(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n364_), .B1(new_n373_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n376_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n302_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n366_), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n305_), .A2(new_n379_), .B1(new_n381_), .B2(new_n374_), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n371_), .A2(KEYINPUT72), .A3(new_n368_), .ZN(new_n383_));
  AOI21_X1  g182(.A(KEYINPUT72), .B1(new_n371_), .B2(new_n368_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n382_), .A2(new_n385_), .A3(KEYINPUT73), .ZN(new_n386_));
  INV_X1    g185(.A(new_n381_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n369_), .B1(new_n387_), .B2(new_n367_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n378_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G120gat), .B(G148gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT5), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G176gat), .B(G204gat), .ZN(new_n392_));
  XOR2_X1   g191(.A(new_n391_), .B(new_n392_), .Z(new_n393_));
  NAND2_X1  g192(.A1(new_n389_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n393_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n378_), .A2(new_n386_), .A3(new_n388_), .A4(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(KEYINPUT74), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT74), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n389_), .A2(new_n398_), .A3(new_n393_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT13), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT13), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n397_), .A2(new_n402_), .A3(new_n399_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n329_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n328_), .B(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT83), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n257_), .A2(new_n408_), .A3(new_n264_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n408_), .B1(new_n257_), .B2(new_n264_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n407_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT83), .B1(new_n284_), .B2(new_n285_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n257_), .A2(new_n264_), .A3(new_n408_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n412_), .A2(new_n330_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n411_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G229gat), .A2(G233gat), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n416_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n330_), .B1(new_n286_), .B2(new_n288_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n418_), .B1(new_n419_), .B2(new_n411_), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n417_), .A2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G113gat), .B(G141gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G169gat), .B(G197gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n421_), .B(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n405_), .A2(new_n426_), .ZN(new_n427_));
  XOR2_X1   g226(.A(G211gat), .B(G218gat), .Z(new_n428_));
  INV_X1    g227(.A(KEYINPUT21), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  XOR2_X1   g229(.A(G197gat), .B(G204gat), .Z(new_n431_));
  XNOR2_X1  g230(.A(G211gat), .B(G218gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT21), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n430_), .A2(new_n431_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n431_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n435_), .A2(KEYINPUT21), .A3(new_n432_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G141gat), .A2(G148gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT84), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT84), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n440_), .A2(G141gat), .A3(G148gat), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT2), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n439_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT87), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT86), .B1(new_n445_), .B2(KEYINPUT3), .ZN(new_n446_));
  NOR2_X1   g245(.A1(G141gat), .A2(G148gat), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT86), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n450_), .B1(G141gat), .B2(G148gat), .ZN(new_n451_));
  AOI21_X1  g250(.A(KEYINPUT3), .B1(new_n451_), .B2(new_n445_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n443_), .B(new_n444_), .C1(new_n449_), .C2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(G155gat), .A2(G162gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT85), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G155gat), .A2(G162gat), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  XOR2_X1   g256(.A(new_n456_), .B(KEYINPUT1), .Z(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n455_), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n448_), .A2(new_n439_), .A3(new_n441_), .ZN(new_n460_));
  AOI22_X1  g259(.A1(new_n453_), .A2(new_n457_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT29), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n437_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(G228gat), .A3(G233gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G228gat), .A2(G233gat), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n465_), .B(new_n437_), .C1(new_n461_), .C2(new_n462_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT88), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n464_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G78gat), .B(G106gat), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n464_), .A2(new_n466_), .A3(new_n467_), .A4(new_n469_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n467_), .B1(new_n464_), .B2(new_n466_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT28), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n475_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n461_), .A2(new_n475_), .A3(new_n462_), .ZN(new_n478_));
  XOR2_X1   g277(.A(G22gat), .B(G50gat), .Z(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n477_), .A2(new_n478_), .A3(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n478_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n479_), .B1(new_n482_), .B2(new_n476_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n474_), .B1(new_n481_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n473_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G127gat), .B(G134gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G113gat), .B(G120gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G183gat), .A2(G190gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT23), .ZN(new_n491_));
  OR2_X1    g290(.A1(G183gat), .A2(G190gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G169gat), .A2(G176gat), .ZN(new_n495_));
  XOR2_X1   g294(.A(KEYINPUT22), .B(G169gat), .Z(new_n496_));
  OAI21_X1  g295(.A(new_n495_), .B1(new_n496_), .B2(G176gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT25), .B(G183gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT26), .B(G190gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(new_n491_), .ZN(new_n501_));
  INV_X1    g300(.A(G169gat), .ZN(new_n502_));
  INV_X1    g301(.A(G176gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n504_), .A2(KEYINPUT24), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(KEYINPUT24), .A3(new_n495_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  OAI22_X1  g306(.A1(new_n494_), .A2(new_n497_), .B1(new_n501_), .B2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT30), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  OR2_X1    g309(.A1(new_n501_), .A2(new_n507_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n493_), .B(new_n495_), .C1(G176gat), .C2(new_n496_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(KEYINPUT30), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G71gat), .B(G99gat), .ZN(new_n515_));
  INV_X1    g314(.A(G43gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G227gat), .A2(G233gat), .ZN(new_n518_));
  INV_X1    g317(.A(G15gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n517_), .B(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n514_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n521_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n523_), .A2(new_n510_), .A3(new_n513_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT31), .ZN(new_n525_));
  AND3_X1   g324(.A1(new_n522_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n525_), .B1(new_n522_), .B2(new_n524_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n489_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n522_), .A2(new_n524_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT31), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n522_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n488_), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n528_), .A2(new_n532_), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n483_), .A2(new_n481_), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n471_), .B(new_n472_), .C1(new_n534_), .C2(new_n474_), .ZN(new_n535_));
  AND3_X1   g334(.A1(new_n485_), .A2(new_n533_), .A3(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n533_), .B1(new_n485_), .B2(new_n535_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT27), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G8gat), .B(G36gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G64gat), .B(G92gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(KEYINPUT92), .B(KEYINPUT18), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT99), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G226gat), .A2(G233gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT19), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n491_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n499_), .B(KEYINPUT89), .Z(new_n549_));
  INV_X1    g348(.A(new_n498_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n548_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n437_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n496_), .A2(KEYINPUT90), .ZN(new_n553_));
  XNOR2_X1  g352(.A(KEYINPUT22), .B(G169gat), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT90), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n553_), .A2(new_n503_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT91), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n491_), .A2(new_n558_), .A3(new_n492_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n558_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n557_), .B(new_n495_), .C1(new_n559_), .C2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n551_), .A2(new_n552_), .A3(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT20), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n563_), .A2(KEYINPUT97), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n563_), .A2(KEYINPUT97), .B1(new_n508_), .B2(new_n437_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n547_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n552_), .B1(new_n551_), .B2(new_n561_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT20), .B1(new_n508_), .B2(new_n437_), .ZN(new_n568_));
  NOR3_X1   g367(.A1(new_n567_), .A2(new_n546_), .A3(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n544_), .B1(new_n566_), .B2(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n546_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n546_), .B1(new_n508_), .B2(new_n437_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n562_), .A2(new_n572_), .A3(KEYINPUT20), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n571_), .A2(new_n543_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT100), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n538_), .B1(new_n570_), .B2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n571_), .A2(new_n573_), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n578_), .B(new_n543_), .Z(new_n579_));
  NOR2_X1   g378(.A1(new_n579_), .A2(KEYINPUT27), .ZN(new_n580_));
  OAI22_X1  g379(.A1(new_n536_), .A2(new_n537_), .B1(new_n577_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT98), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n453_), .A2(new_n457_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT94), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n459_), .A2(new_n460_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n583_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n586_), .A2(KEYINPUT93), .A3(new_n488_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT93), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n583_), .A2(new_n588_), .A3(new_n585_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(new_n489_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n588_), .B1(new_n461_), .B2(new_n584_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n587_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G225gat), .A2(G233gat), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n592_), .A2(KEYINPUT4), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT95), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n592_), .A2(KEYINPUT95), .A3(KEYINPUT4), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  OR3_X1    g399(.A1(new_n461_), .A2(KEYINPUT4), .A3(new_n488_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n593_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n595_), .B1(new_n600_), .B2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G1gat), .B(G29gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT0), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(new_n343_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(G85gat), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n582_), .B1(new_n605_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n609_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n603_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n612_));
  OAI211_X1 g411(.A(KEYINPUT98), .B(new_n611_), .C1(new_n612_), .C2(new_n595_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n599_), .ZN(new_n614_));
  AOI21_X1  g413(.A(KEYINPUT95), .B1(new_n592_), .B2(KEYINPUT4), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n604_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n616_), .A2(new_n594_), .A3(new_n609_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n610_), .A2(new_n613_), .A3(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n581_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(KEYINPUT96), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(KEYINPUT33), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT33), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n617_), .A2(KEYINPUT96), .A3(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n600_), .A2(new_n593_), .A3(new_n601_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n609_), .B1(new_n602_), .B2(new_n592_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n579_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n621_), .A2(new_n623_), .A3(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n566_), .A2(new_n569_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n543_), .A2(KEYINPUT32), .ZN(new_n629_));
  MUX2_X1   g428(.A(new_n628_), .B(new_n578_), .S(new_n629_), .Z(new_n630_));
  NAND2_X1  g429(.A1(new_n613_), .A2(new_n617_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n616_), .A2(new_n594_), .ZN(new_n632_));
  AOI21_X1  g431(.A(KEYINPUT98), .B1(new_n632_), .B2(new_n611_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n630_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n627_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n485_), .A2(new_n535_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n533_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n619_), .B1(new_n635_), .B2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n427_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n363_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n643_), .A2(new_n325_), .A3(new_n618_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT38), .ZN(new_n645_));
  INV_X1    g444(.A(new_n361_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n427_), .A2(new_n646_), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n297_), .A2(KEYINPUT101), .A3(new_n315_), .ZN(new_n648_));
  AOI21_X1  g447(.A(KEYINPUT101), .B1(new_n297_), .B2(new_n315_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n640_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n647_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n618_), .ZN(new_n654_));
  OAI21_X1  g453(.A(G1gat), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n645_), .A2(new_n655_), .ZN(G1324gat));
  OR2_X1    g455(.A1(new_n577_), .A2(new_n580_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G8gat), .B1(new_n653_), .B2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT39), .ZN(new_n659_));
  INV_X1    g458(.A(new_n657_), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n363_), .A2(new_n326_), .A3(new_n660_), .A4(new_n641_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT102), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n659_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT40), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n663_), .B(new_n664_), .ZN(G1325gat));
  INV_X1    g464(.A(new_n653_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n519_), .B1(new_n666_), .B2(new_n638_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n668_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n643_), .A2(new_n519_), .A3(new_n638_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n669_), .A2(new_n670_), .A3(new_n671_), .ZN(G1326gat));
  OAI21_X1  g471(.A(G22gat), .B1(new_n653_), .B2(new_n636_), .ZN(new_n673_));
  XOR2_X1   g472(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n636_), .A2(G22gat), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n642_), .B2(new_n676_), .ZN(G1327gat));
  NOR2_X1   g476(.A1(new_n650_), .A2(new_n361_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n641_), .A2(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(G29gat), .B1(new_n679_), .B2(new_n618_), .ZN(new_n680_));
  OAI21_X1  g479(.A(KEYINPUT43), .B1(new_n640_), .B2(new_n323_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n322_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n319_), .B2(KEYINPUT37), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT43), .ZN(new_n684_));
  INV_X1    g483(.A(new_n639_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n685_), .B1(new_n627_), .B2(new_n634_), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n683_), .B(new_n684_), .C1(new_n686_), .C2(new_n619_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n681_), .A2(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n427_), .A2(new_n361_), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT44), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n690_), .A2(new_n253_), .A3(new_n654_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n688_), .A2(new_n689_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n680_), .B1(new_n691_), .B2(new_n695_), .ZN(G1328gat));
  NAND3_X1  g495(.A1(new_n679_), .A2(new_n251_), .A3(new_n660_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT45), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n694_), .A2(new_n657_), .A3(new_n690_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n698_), .B1(new_n699_), .B2(new_n251_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  OAI221_X1 g501(.A(new_n698_), .B1(KEYINPUT104), .B2(KEYINPUT46), .C1(new_n251_), .C2(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1329gat));
  AOI21_X1  g503(.A(G43gat), .B1(new_n679_), .B2(new_n638_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n694_), .A2(new_n690_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n533_), .A2(new_n516_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n705_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g508(.A(G50gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n679_), .A2(new_n710_), .A3(new_n637_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n706_), .A2(new_n712_), .A3(new_n637_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(G50gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n712_), .B1(new_n706_), .B2(new_n637_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n711_), .B1(new_n714_), .B2(new_n715_), .ZN(G1331gat));
  NOR3_X1   g515(.A1(new_n640_), .A2(new_n405_), .A3(new_n426_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n363_), .A2(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n718_), .A2(new_n343_), .A3(new_n618_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n405_), .A2(new_n426_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n652_), .A2(new_n720_), .A3(new_n361_), .ZN(new_n721_));
  OAI21_X1  g520(.A(G57gat), .B1(new_n721_), .B2(new_n654_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n719_), .A2(new_n722_), .ZN(G1332gat));
  OAI21_X1  g522(.A(G64gat), .B1(new_n721_), .B2(new_n657_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT48), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n718_), .A2(new_n341_), .A3(new_n660_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1333gat));
  OAI21_X1  g526(.A(G71gat), .B1(new_n721_), .B2(new_n533_), .ZN(new_n728_));
  XOR2_X1   g527(.A(KEYINPUT106), .B(KEYINPUT49), .Z(new_n729_));
  XNOR2_X1  g528(.A(new_n728_), .B(new_n729_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n533_), .A2(G71gat), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT107), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n718_), .A2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n730_), .A2(new_n733_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT108), .Z(G1334gat));
  NAND3_X1  g534(.A1(new_n718_), .A2(new_n339_), .A3(new_n637_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n721_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n339_), .B1(new_n737_), .B2(new_n637_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT50), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n738_), .A2(new_n739_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n736_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT109), .ZN(G1335gat));
  NAND2_X1  g542(.A1(new_n688_), .A2(KEYINPUT110), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n681_), .A2(new_n745_), .A3(new_n687_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n426_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n404_), .A2(new_n747_), .A3(new_n646_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n744_), .A2(new_n746_), .A3(new_n749_), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n750_), .B(new_n618_), .C1(new_n214_), .C2(new_n213_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n717_), .A2(new_n678_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n216_), .B1(new_n753_), .B2(new_n654_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n751_), .A2(new_n754_), .ZN(G1336gat));
  AOI21_X1  g554(.A(G92gat), .B1(new_n752_), .B2(new_n660_), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT111), .Z(new_n757_));
  NOR2_X1   g556(.A1(new_n657_), .A2(new_n211_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n750_), .B2(new_n758_), .ZN(G1337gat));
  NAND4_X1  g558(.A1(new_n744_), .A2(new_n638_), .A3(new_n746_), .A4(new_n749_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(G99gat), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n533_), .A2(new_n209_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n752_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT113), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n766_), .A2(KEYINPUT112), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT113), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n761_), .A2(new_n768_), .A3(new_n763_), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n765_), .A2(new_n767_), .A3(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n767_), .B1(new_n765_), .B2(new_n769_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n770_), .A2(new_n771_), .ZN(G1338gat));
  AND2_X1   g571(.A1(new_n681_), .A2(new_n687_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n404_), .A2(new_n637_), .A3(new_n747_), .A4(new_n646_), .ZN(new_n774_));
  OAI21_X1  g573(.A(KEYINPUT114), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n681_), .B2(new_n687_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n229_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n775_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n775_), .A2(new_n778_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT52), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n775_), .A2(new_n778_), .A3(KEYINPUT115), .A4(new_n779_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n782_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n752_), .A2(new_n229_), .A3(new_n637_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT53), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n786_), .A2(new_n790_), .A3(new_n787_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(G1339gat));
  INV_X1    g591(.A(KEYINPUT120), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT117), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n418_), .B1(new_n411_), .B2(new_n414_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n794_), .B1(new_n795_), .B2(new_n425_), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n409_), .A2(new_n410_), .A3(new_n407_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n330_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n416_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n799_), .A2(KEYINPUT117), .A3(new_n424_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n419_), .A2(new_n418_), .A3(new_n411_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT118), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n796_), .A2(new_n800_), .A3(new_n802_), .A4(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n425_), .B1(new_n417_), .B2(new_n420_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n425_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n801_), .B1(new_n807_), .B2(KEYINPUT117), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n803_), .B1(new_n808_), .B2(new_n796_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n806_), .A2(new_n809_), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n810_), .A2(KEYINPUT119), .A3(new_n396_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT119), .B1(new_n810_), .B2(new_n396_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n371_), .B(new_n375_), .C1(new_n283_), .C2(new_n376_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n369_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT116), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n814_), .A2(new_n817_), .A3(new_n369_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n378_), .A2(new_n386_), .A3(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n382_), .A2(new_n385_), .A3(KEYINPUT55), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n819_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT56), .B1(new_n823_), .B2(new_n393_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT56), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n373_), .A2(new_n377_), .A3(new_n820_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n826_), .B1(new_n816_), .B2(new_n818_), .ZN(new_n827_));
  AOI211_X1 g626(.A(new_n825_), .B(new_n395_), .C1(new_n827_), .C2(new_n821_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n813_), .B(KEYINPUT58), .C1(new_n824_), .C2(new_n828_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n829_), .A2(new_n683_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT58), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n828_), .A2(new_n824_), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n811_), .A2(new_n812_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n831_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n396_), .A2(new_n426_), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n378_), .A2(new_n386_), .A3(new_n820_), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n814_), .A2(new_n817_), .A3(new_n369_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n817_), .B1(new_n814_), .B2(new_n369_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n822_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n393_), .B1(new_n837_), .B2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n825_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n823_), .A2(KEYINPUT56), .A3(new_n393_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n836_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n397_), .A2(new_n399_), .A3(new_n810_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n650_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n830_), .A2(new_n834_), .B1(new_n835_), .B2(new_n846_), .ZN(new_n847_));
  OAI211_X1 g646(.A(KEYINPUT57), .B(new_n650_), .C1(new_n844_), .C2(new_n845_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n361_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n401_), .A2(new_n747_), .A3(new_n403_), .ZN(new_n850_));
  NOR4_X1   g649(.A1(new_n850_), .A2(new_n683_), .A3(KEYINPUT54), .A4(new_n646_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n646_), .B1(new_n320_), .B2(new_n322_), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n401_), .A2(new_n747_), .A3(new_n403_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n852_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n851_), .A2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n793_), .B1(new_n849_), .B2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n846_), .A2(new_n835_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n834_), .A2(new_n683_), .A3(new_n829_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n858_), .A2(new_n859_), .A3(new_n848_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n646_), .ZN(new_n861_));
  OAI21_X1  g660(.A(KEYINPUT54), .B1(new_n362_), .B2(new_n850_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n853_), .A2(new_n854_), .A3(new_n852_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n861_), .A2(KEYINPUT120), .A3(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n660_), .A2(new_n654_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n537_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n857_), .A2(new_n865_), .A3(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(KEYINPUT59), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n856_), .B1(new_n861_), .B2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n860_), .A2(KEYINPUT121), .A3(new_n646_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n867_), .A2(KEYINPUT59), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n871_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n876_), .ZN(new_n878_));
  AOI211_X1 g677(.A(KEYINPUT122), .B(new_n878_), .C1(new_n873_), .C2(new_n874_), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n870_), .B(new_n426_), .C1(new_n877_), .C2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(G113gat), .ZN(new_n881_));
  OR3_X1    g680(.A1(new_n869_), .A2(G113gat), .A3(new_n747_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(G1340gat));
  OAI211_X1 g682(.A(new_n870_), .B(new_n404_), .C1(new_n877_), .C2(new_n879_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(G120gat), .ZN(new_n885_));
  INV_X1    g684(.A(new_n869_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT60), .ZN(new_n887_));
  INV_X1    g686(.A(G120gat), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n404_), .A2(new_n887_), .A3(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n889_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n886_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n885_), .A2(new_n891_), .ZN(G1341gat));
  AOI21_X1  g691(.A(G127gat), .B1(new_n886_), .B2(new_n361_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n877_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n879_), .ZN(new_n895_));
  AOI22_X1  g694(.A1(new_n894_), .A2(new_n895_), .B1(KEYINPUT59), .B2(new_n869_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT123), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n361_), .A2(new_n897_), .A3(G127gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n898_), .B1(new_n897_), .B2(G127gat), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n893_), .B1(new_n896_), .B2(new_n899_), .ZN(G1342gat));
  INV_X1    g699(.A(G134gat), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n323_), .A2(new_n901_), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n870_), .B(new_n902_), .C1(new_n877_), .C2(new_n879_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n901_), .B1(new_n869_), .B2(new_n650_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(KEYINPUT124), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT124), .ZN(new_n906_));
  OAI211_X1 g705(.A(new_n906_), .B(new_n901_), .C1(new_n869_), .C2(new_n650_), .ZN(new_n907_));
  AND3_X1   g706(.A1(new_n903_), .A2(new_n905_), .A3(new_n907_), .ZN(G1343gat));
  AND3_X1   g707(.A1(new_n861_), .A2(KEYINPUT120), .A3(new_n864_), .ZN(new_n909_));
  AOI21_X1  g708(.A(KEYINPUT120), .B1(new_n861_), .B2(new_n864_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n536_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n909_), .A2(new_n910_), .A3(new_n911_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n912_), .A2(new_n426_), .A3(new_n866_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g713(.A1(new_n912_), .A2(new_n404_), .A3(new_n866_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g715(.A1(new_n912_), .A2(new_n361_), .A3(new_n866_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(KEYINPUT61), .B(G155gat), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n917_), .B(new_n918_), .ZN(G1346gat));
  NAND2_X1  g718(.A1(new_n912_), .A2(new_n866_), .ZN(new_n920_));
  OAI21_X1  g719(.A(G162gat), .B1(new_n920_), .B2(new_n323_), .ZN(new_n921_));
  OR2_X1    g720(.A1(new_n650_), .A2(G162gat), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n920_), .B2(new_n922_), .ZN(G1347gat));
  INV_X1    g722(.A(KEYINPUT62), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n657_), .A2(new_n618_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n925_), .A2(new_n638_), .A3(new_n636_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n926_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(new_n426_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n924_), .B1(new_n929_), .B2(new_n502_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n928_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n929_), .A2(new_n553_), .A3(new_n556_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n930_), .A2(new_n931_), .A3(new_n932_), .ZN(G1348gat));
  AOI21_X1  g732(.A(G176gat), .B1(new_n927_), .B2(new_n404_), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n909_), .A2(new_n910_), .A3(new_n926_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n405_), .A2(new_n503_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n934_), .B1(new_n935_), .B2(new_n936_), .ZN(G1349gat));
  AOI21_X1  g736(.A(G183gat), .B1(new_n935_), .B2(new_n361_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n646_), .A2(new_n498_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n938_), .B1(new_n927_), .B2(new_n939_), .ZN(G1350gat));
  INV_X1    g739(.A(new_n549_), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n927_), .A2(new_n941_), .A3(new_n651_), .ZN(new_n942_));
  AND2_X1   g741(.A1(new_n927_), .A2(new_n683_), .ZN(new_n943_));
  INV_X1    g742(.A(G190gat), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n942_), .B1(new_n943_), .B2(new_n944_), .ZN(G1351gat));
  INV_X1    g744(.A(KEYINPUT125), .ZN(new_n946_));
  INV_X1    g745(.A(G197gat), .ZN(new_n947_));
  NAND4_X1  g746(.A1(new_n857_), .A2(new_n536_), .A3(new_n865_), .A4(new_n925_), .ZN(new_n948_));
  OAI211_X1 g747(.A(new_n946_), .B(new_n947_), .C1(new_n948_), .C2(new_n747_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n912_), .A2(new_n426_), .A3(new_n925_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n949_), .B1(new_n950_), .B2(new_n947_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n946_), .B1(new_n950_), .B2(new_n947_), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n951_), .A2(new_n952_), .ZN(G1352gat));
  NOR2_X1   g752(.A1(new_n948_), .A2(new_n405_), .ZN(new_n954_));
  XOR2_X1   g753(.A(new_n954_), .B(G204gat), .Z(G1353gat));
  NAND2_X1  g754(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n361_), .A2(new_n956_), .ZN(new_n957_));
  XOR2_X1   g756(.A(new_n957_), .B(KEYINPUT126), .Z(new_n958_));
  NOR2_X1   g757(.A1(new_n948_), .A2(new_n958_), .ZN(new_n959_));
  NOR2_X1   g758(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n959_), .B(new_n960_), .ZN(G1354gat));
  OAI21_X1  g760(.A(G218gat), .B1(new_n948_), .B2(new_n323_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n650_), .A2(G218gat), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n912_), .A2(new_n925_), .A3(new_n963_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n962_), .A2(new_n964_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n965_), .A2(KEYINPUT127), .ZN(new_n966_));
  INV_X1    g765(.A(KEYINPUT127), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n962_), .A2(new_n964_), .A3(new_n967_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n966_), .A2(new_n968_), .ZN(G1355gat));
endmodule


