//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n781_, new_n782_, new_n783_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n940_, new_n941_, new_n943_, new_n944_, new_n945_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n953_, new_n954_,
    new_n956_, new_n957_, new_n958_, new_n960_, new_n961_, new_n962_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_, new_n986_, new_n988_, new_n989_,
    new_n990_, new_n992_, new_n993_, new_n994_, new_n996_, new_n997_,
    new_n998_, new_n999_, new_n1001_, new_n1002_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1010_, new_n1011_, new_n1012_;
  AND2_X1   g000(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n202_));
  NOR2_X1   g001(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n203_));
  OAI22_X1  g002(.A1(new_n202_), .A2(new_n203_), .B1(G99gat), .B2(G106gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT6), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(G99gat), .A3(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n204_), .A2(new_n209_), .A3(new_n212_), .ZN(new_n213_));
  XOR2_X1   g012(.A(new_n213_), .B(KEYINPUT66), .Z(new_n214_));
  XNOR2_X1  g013(.A(G85gat), .B(G92gat), .ZN(new_n215_));
  XOR2_X1   g014(.A(new_n215_), .B(KEYINPUT67), .Z(new_n216_));
  INV_X1    g015(.A(KEYINPUT8), .ZN(new_n217_));
  AND2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT7), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n210_), .B1(new_n222_), .B2(new_n211_), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n210_), .A2(new_n211_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT69), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT69), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n204_), .A2(new_n226_), .A3(new_n212_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n206_), .A2(new_n208_), .A3(KEYINPUT68), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT68), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n209_), .A2(new_n229_), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n225_), .A2(new_n227_), .A3(new_n228_), .A4(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n231_), .A2(KEYINPUT70), .A3(new_n216_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT8), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT70), .B1(new_n231_), .B2(new_n216_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n219_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT9), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n215_), .A2(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(KEYINPUT10), .B(G99gat), .Z(new_n238_));
  INV_X1    g037(.A(G106gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n236_), .A2(G85gat), .A3(G92gat), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n237_), .A2(new_n240_), .A3(new_n209_), .A4(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n235_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G57gat), .B(G64gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT11), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G71gat), .B(G78gat), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n245_), .A2(new_n247_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n244_), .A2(KEYINPUT11), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n249_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n243_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT71), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n235_), .A2(new_n252_), .A3(new_n242_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n254_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G230gat), .A2(G233gat), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n258_), .B(KEYINPUT64), .Z(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n243_), .A2(KEYINPUT71), .A3(new_n253_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n257_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(G120gat), .B(G148gat), .Z(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT5), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G176gat), .B(G204gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT72), .ZN(new_n267_));
  INV_X1    g066(.A(new_n242_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n231_), .A2(new_n216_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT70), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n271_), .A2(KEYINPUT8), .A3(new_n232_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n268_), .B1(new_n272_), .B2(new_n219_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n260_), .B1(new_n273_), .B2(new_n252_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT12), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n275_), .B1(new_n243_), .B2(new_n253_), .ZN(new_n276_));
  AOI211_X1 g075(.A(KEYINPUT12), .B(new_n252_), .C1(new_n235_), .C2(new_n242_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n274_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n262_), .A2(new_n267_), .A3(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n267_), .B1(new_n262_), .B2(new_n278_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT13), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT14), .ZN(new_n283_));
  INV_X1    g082(.A(G8gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT75), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT75), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(G8gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n283_), .B1(new_n288_), .B2(G1gat), .ZN(new_n289_));
  XOR2_X1   g088(.A(G15gat), .B(G22gat), .Z(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT76), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT77), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT75), .B(G8gat), .ZN(new_n293_));
  INV_X1    g092(.A(G1gat), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT14), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT76), .ZN(new_n296_));
  INV_X1    g095(.A(new_n290_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n295_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  AND3_X1   g097(.A1(new_n291_), .A2(new_n292_), .A3(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n292_), .B1(new_n291_), .B2(new_n298_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G1gat), .B(G8gat), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NOR3_X1   g101(.A1(new_n299_), .A2(new_n300_), .A3(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n291_), .A2(new_n298_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT77), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n291_), .A2(new_n292_), .A3(new_n298_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n301_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n303_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(G231gat), .ZN(new_n309_));
  INV_X1    g108(.A(G233gat), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n308_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n302_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n305_), .A2(new_n301_), .A3(new_n306_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(G231gat), .A3(G233gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n311_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n252_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n311_), .A2(new_n253_), .A3(new_n315_), .ZN(new_n318_));
  XOR2_X1   g117(.A(G127gat), .B(G155gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT16), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G183gat), .B(G211gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT17), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n317_), .A2(new_n318_), .A3(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT78), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n317_), .A2(new_n318_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n322_), .B(KEYINPUT17), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n326_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G29gat), .B(G36gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G43gat), .B(G50gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n235_), .A2(new_n333_), .A3(new_n242_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G232gat), .A2(G233gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT34), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT35), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n333_), .B(KEYINPUT15), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n334_), .B(new_n339_), .C1(new_n273_), .C2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n342_), .A2(KEYINPUT73), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT73), .ZN(new_n344_));
  AOI22_X1  g143(.A1(new_n243_), .A2(new_n340_), .B1(new_n338_), .B2(new_n337_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n344_), .B1(new_n345_), .B2(new_n334_), .ZN(new_n346_));
  OAI22_X1  g145(.A1(new_n343_), .A2(new_n346_), .B1(new_n338_), .B2(new_n337_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n342_), .A2(KEYINPUT73), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n345_), .A2(new_n344_), .A3(new_n334_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n337_), .A2(new_n338_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n348_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT74), .B1(new_n347_), .B2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G190gat), .B(G218gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G134gat), .B(G162gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT36), .B1(new_n352_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT74), .ZN(new_n357_));
  INV_X1    g156(.A(new_n351_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n350_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n357_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT36), .ZN(new_n361_));
  INV_X1    g160(.A(new_n355_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n360_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n362_), .B1(new_n347_), .B2(new_n351_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n356_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT37), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n347_), .A2(new_n351_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n355_), .B1(new_n369_), .B2(new_n357_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n364_), .B1(new_n370_), .B2(new_n361_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n371_), .A2(KEYINPUT37), .A3(new_n356_), .ZN(new_n372_));
  AOI211_X1 g171(.A(new_n282_), .B(new_n330_), .C1(new_n368_), .C2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT80), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n374_), .B1(new_n314_), .B2(new_n341_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n312_), .A2(new_n313_), .A3(KEYINPUT80), .A4(new_n340_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G229gat), .A2(G233gat), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n379_), .B1(new_n314_), .B2(new_n333_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n377_), .A2(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n333_), .B1(new_n303_), .B2(new_n307_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT79), .ZN(new_n383_));
  INV_X1    g182(.A(new_n333_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n312_), .A2(new_n313_), .A3(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n382_), .A2(new_n383_), .A3(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n308_), .A2(KEYINPUT79), .A3(new_n384_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n386_), .A2(new_n379_), .A3(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(G113gat), .B(G141gat), .Z(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT81), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G169gat), .B(G197gat), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n390_), .B(new_n391_), .Z(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n381_), .A2(new_n388_), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n393_), .B1(new_n381_), .B2(new_n388_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT108), .ZN(new_n398_));
  XOR2_X1   g197(.A(G197gat), .B(G204gat), .Z(new_n399_));
  NAND3_X1  g198(.A1(new_n399_), .A2(KEYINPUT98), .A3(KEYINPUT21), .ZN(new_n400_));
  XOR2_X1   g199(.A(G211gat), .B(G218gat), .Z(new_n401_));
  OAI22_X1  g200(.A1(new_n400_), .A2(new_n401_), .B1(KEYINPUT21), .B2(new_n399_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n400_), .A2(new_n401_), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G155gat), .A2(G162gat), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(G155gat), .A2(G162gat), .ZN(new_n407_));
  OR2_X1    g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  OR2_X1    g207(.A1(new_n408_), .A2(KEYINPUT96), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(KEYINPUT96), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT94), .ZN(new_n411_));
  NOR2_X1   g210(.A1(G141gat), .A2(G148gat), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n411_), .B1(new_n413_), .B2(KEYINPUT3), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G141gat), .A2(G148gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT2), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT3), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n412_), .A2(KEYINPUT94), .A3(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n413_), .A2(KEYINPUT3), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n414_), .A2(new_n417_), .A3(new_n419_), .A4(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT95), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n409_), .B(new_n410_), .C1(new_n421_), .C2(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n416_), .A2(new_n412_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n405_), .B1(new_n407_), .B2(KEYINPUT1), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT1), .ZN(new_n428_));
  AOI22_X1  g227(.A1(new_n427_), .A2(KEYINPUT92), .B1(new_n428_), .B2(new_n406_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT92), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n430_), .B(new_n405_), .C1(new_n407_), .C2(KEYINPUT1), .ZN(new_n431_));
  AOI211_X1 g230(.A(KEYINPUT93), .B(new_n426_), .C1(new_n429_), .C2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT93), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n427_), .A2(KEYINPUT92), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n406_), .A2(new_n428_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n434_), .A2(new_n431_), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n433_), .B1(new_n436_), .B2(new_n425_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n424_), .B1(new_n432_), .B2(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n404_), .B1(new_n438_), .B2(KEYINPUT29), .ZN(new_n439_));
  INV_X1    g238(.A(G228gat), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n440_), .A2(new_n310_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n439_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  AOI211_X1 g243(.A(new_n441_), .B(new_n404_), .C1(new_n438_), .C2(KEYINPUT29), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G78gat), .B(G106gat), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n444_), .A2(new_n446_), .A3(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n447_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n443_), .A2(new_n445_), .ZN(new_n452_));
  AOI21_X1  g251(.A(KEYINPUT99), .B1(new_n452_), .B2(new_n448_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G22gat), .B(G50gat), .ZN(new_n454_));
  OR3_X1    g253(.A1(new_n438_), .A2(KEYINPUT29), .A3(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n454_), .B1(new_n438_), .B2(KEYINPUT29), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  XOR2_X1   g256(.A(KEYINPUT97), .B(KEYINPUT28), .Z(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n455_), .A2(new_n458_), .A3(new_n456_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n451_), .B1(new_n453_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n461_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n458_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n466_), .A2(KEYINPUT99), .A3(new_n449_), .A4(new_n450_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n463_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT27), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G8gat), .B(G36gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT18), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G64gat), .B(G92gat), .ZN(new_n473_));
  XOR2_X1   g272(.A(new_n472_), .B(new_n473_), .Z(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G226gat), .A2(G233gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT19), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT88), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT85), .ZN(new_n479_));
  INV_X1    g278(.A(G169gat), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT22), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(G176gat), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT22), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n483_), .A2(KEYINPUT85), .A3(G169gat), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n481_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G169gat), .A2(G176gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT84), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT84), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(G169gat), .A3(G176gat), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n485_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT86), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT86), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n485_), .A2(new_n490_), .A3(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(G183gat), .A2(G190gat), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G183gat), .A2(G190gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT23), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT23), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n499_), .A2(G183gat), .A3(G190gat), .ZN(new_n500_));
  AOI21_X1  g299(.A(KEYINPUT87), .B1(new_n498_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT87), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n502_), .B1(new_n497_), .B2(KEYINPUT23), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n496_), .B1(new_n501_), .B2(new_n503_), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n492_), .A2(new_n494_), .A3(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n507_), .A2(new_n487_), .A3(new_n489_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n498_), .A2(new_n500_), .ZN(new_n509_));
  NOR3_X1   g308(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n508_), .A2(new_n509_), .A3(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(KEYINPUT26), .B(G190gat), .Z(new_n513_));
  INV_X1    g312(.A(KEYINPUT82), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT83), .ZN(new_n516_));
  XNOR2_X1  g315(.A(KEYINPUT25), .B(G183gat), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT26), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT82), .B1(new_n518_), .B2(G190gat), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n515_), .A2(new_n516_), .A3(new_n517_), .A4(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT26), .B(G190gat), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n517_), .B(new_n519_), .C1(new_n521_), .C2(KEYINPUT82), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT83), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n512_), .B1(new_n520_), .B2(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n478_), .B1(new_n505_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n512_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n522_), .A2(KEYINPUT83), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n522_), .A2(KEYINPUT83), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n526_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n492_), .A2(new_n494_), .A3(new_n504_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(KEYINPUT88), .A3(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n404_), .B1(new_n525_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n509_), .A2(new_n496_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT22), .B(G169gat), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(new_n482_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n533_), .A2(new_n490_), .A3(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n404_), .A2(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n510_), .B1(new_n507_), .B2(new_n486_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n521_), .A2(new_n517_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n501_), .A2(new_n503_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT20), .B1(new_n537_), .B2(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n477_), .B1(new_n532_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT106), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT106), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n546_), .B(new_n477_), .C1(new_n532_), .C2(new_n543_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT20), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT100), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n549_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NOR3_X1   g350(.A1(new_n540_), .A2(new_n541_), .A3(new_n549_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n536_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n404_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n548_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n525_), .A2(new_n404_), .A3(new_n531_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n477_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n545_), .A2(new_n547_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT101), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n477_), .A2(new_n548_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n561_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n560_), .B1(new_n532_), .B2(new_n562_), .ZN(new_n563_));
  NOR3_X1   g362(.A1(new_n505_), .A2(new_n524_), .A3(new_n478_), .ZN(new_n564_));
  AOI21_X1  g363(.A(KEYINPUT88), .B1(new_n529_), .B2(new_n530_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n554_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n561_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n536_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n542_), .A2(KEYINPUT100), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n568_), .B1(new_n569_), .B2(new_n550_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n567_), .B1(new_n570_), .B2(new_n404_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n566_), .A2(KEYINPUT101), .A3(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n563_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n555_), .A2(new_n556_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(new_n477_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n573_), .A2(new_n575_), .A3(new_n474_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT107), .ZN(new_n577_));
  AOI22_X1  g376(.A1(new_n475_), .A2(new_n559_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n573_), .A2(KEYINPUT107), .A3(new_n575_), .A4(new_n474_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n470_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n573_), .A2(new_n575_), .A3(new_n474_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n474_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n581_), .A2(new_n582_), .A3(KEYINPUT27), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n469_), .B1(new_n580_), .B2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G127gat), .B(G134gat), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n585_), .A2(KEYINPUT91), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(KEYINPUT91), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G113gat), .B(G120gat), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n586_), .A2(new_n587_), .A3(new_n589_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT31), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G227gat), .A2(G233gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(G15gat), .ZN(new_n597_));
  INV_X1    g396(.A(G71gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(G99gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT89), .B(G43gat), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n600_), .A2(new_n601_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT90), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n525_), .A2(KEYINPUT30), .A3(new_n531_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(KEYINPUT30), .B1(new_n525_), .B2(new_n531_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n605_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT30), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n610_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n611_), .A2(KEYINPUT90), .A3(new_n606_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n604_), .B1(new_n609_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n604_), .ZN(new_n614_));
  AOI21_X1  g413(.A(KEYINPUT90), .B1(new_n611_), .B2(new_n606_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n595_), .B1(new_n613_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n612_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n614_), .B1(new_n618_), .B2(new_n615_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n609_), .A2(new_n604_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(new_n620_), .A3(new_n594_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n617_), .A2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G1gat), .B(G29gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(G85gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT0), .B(G57gat), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n624_), .B(new_n625_), .Z(new_n626_));
  NAND2_X1  g425(.A1(G225gat), .A2(G233gat), .ZN(new_n627_));
  AOI21_X1  g426(.A(KEYINPUT4), .B1(new_n438_), .B2(new_n593_), .ZN(new_n628_));
  OAI21_X1  g427(.A(KEYINPUT103), .B1(new_n438_), .B2(new_n593_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n432_), .A2(new_n437_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT103), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n591_), .A2(new_n592_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n630_), .A2(new_n631_), .A3(new_n632_), .A4(new_n424_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT102), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n438_), .A2(new_n634_), .A3(new_n593_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n634_), .B1(new_n438_), .B2(new_n593_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n629_), .B(new_n633_), .C1(new_n635_), .C2(new_n636_), .ZN(new_n637_));
  AOI211_X1 g436(.A(new_n627_), .B(new_n628_), .C1(new_n637_), .C2(KEYINPUT4), .ZN(new_n638_));
  INV_X1    g437(.A(new_n627_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n633_), .A2(new_n629_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n636_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n438_), .A2(new_n634_), .A3(new_n593_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n639_), .B1(new_n640_), .B2(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n626_), .B1(new_n638_), .B2(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n628_), .B1(new_n637_), .B2(KEYINPUT4), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n644_), .B1(new_n646_), .B2(new_n639_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n626_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n622_), .A2(new_n645_), .A3(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n398_), .B1(new_n584_), .B2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n559_), .A2(new_n475_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n576_), .A2(new_n577_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n652_), .A2(new_n653_), .A3(new_n579_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT27), .ZN(new_n655_));
  INV_X1    g454(.A(new_n583_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n468_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n650_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n657_), .A2(KEYINPUT108), .A3(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n651_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n622_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n646_), .A2(new_n639_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n648_), .B1(new_n637_), .B2(new_n627_), .ZN(new_n663_));
  OAI21_X1  g462(.A(KEYINPUT104), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT4), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n665_), .B1(new_n640_), .B2(new_n643_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n627_), .B1(new_n666_), .B2(new_n628_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT104), .ZN(new_n668_));
  INV_X1    g467(.A(new_n663_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n667_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n664_), .A2(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n581_), .A2(new_n582_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT33), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n646_), .A2(new_n639_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n644_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n673_), .B1(new_n676_), .B2(new_n626_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n647_), .A2(KEYINPUT33), .A3(new_n648_), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n671_), .B(new_n672_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n474_), .A2(KEYINPUT32), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n573_), .A2(new_n575_), .A3(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n680_), .ZN(new_n684_));
  AOI22_X1  g483(.A1(new_n559_), .A2(new_n684_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n676_), .A2(new_n626_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n647_), .A2(new_n648_), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n683_), .B(new_n685_), .C1(new_n686_), .C2(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n468_), .B1(new_n679_), .B2(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n468_), .A2(new_n645_), .A3(new_n649_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n690_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n661_), .B1(new_n689_), .B2(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n397_), .B1(new_n660_), .B2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n373_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT109), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n686_), .A2(new_n687_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n373_), .A2(KEYINPUT109), .A3(new_n693_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n696_), .A2(new_n294_), .A3(new_n698_), .A4(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT38), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n366_), .B1(new_n660_), .B2(new_n692_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n282_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n397_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n706_), .A2(new_n330_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n703_), .A2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(G1gat), .B1(new_n708_), .B2(new_n697_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n700_), .A2(new_n701_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n702_), .A2(new_n709_), .A3(new_n710_), .ZN(G1324gat));
  AOI21_X1  g510(.A(new_n583_), .B1(new_n654_), .B2(KEYINPUT27), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n696_), .A2(new_n712_), .A3(new_n293_), .A4(new_n699_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n703_), .A2(new_n712_), .A3(new_n707_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT110), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n715_), .A2(KEYINPUT39), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n284_), .B1(new_n715_), .B2(KEYINPUT39), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n714_), .A2(new_n716_), .A3(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n716_), .B1(new_n714_), .B2(new_n717_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n713_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  XOR2_X1   g519(.A(new_n720_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g520(.A(G15gat), .B1(new_n708_), .B2(new_n661_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT41), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n694_), .A2(G15gat), .A3(new_n661_), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1326gat));
  OAI21_X1  g524(.A(G22gat), .B1(new_n708_), .B2(new_n469_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT42), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n469_), .A2(G22gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n727_), .B1(new_n694_), .B2(new_n728_), .ZN(G1327gat));
  INV_X1    g528(.A(KEYINPUT111), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT37), .B1(new_n371_), .B2(new_n356_), .ZN(new_n731_));
  AND4_X1   g530(.A1(KEYINPUT37), .A2(new_n356_), .A3(new_n363_), .A4(new_n365_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n730_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n677_), .A2(new_n678_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n662_), .A2(KEYINPUT104), .A3(new_n663_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n668_), .B1(new_n667_), .B2(new_n669_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n672_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n688_), .B1(new_n734_), .B2(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n691_), .B1(new_n738_), .B2(new_n469_), .ZN(new_n739_));
  AOI21_X1  g538(.A(KEYINPUT108), .B1(new_n657_), .B2(new_n658_), .ZN(new_n740_));
  NOR4_X1   g539(.A1(new_n712_), .A2(new_n650_), .A3(new_n398_), .A4(new_n468_), .ZN(new_n741_));
  OAI22_X1  g540(.A1(new_n739_), .A2(new_n622_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n368_), .A2(new_n372_), .A3(KEYINPUT111), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n733_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT43), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT43), .B1(new_n660_), .B2(new_n692_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n731_), .A2(new_n732_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n745_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n330_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n706_), .A2(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n749_), .A2(KEYINPUT44), .A3(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n753_));
  AOI22_X1  g552(.A1(new_n744_), .A2(KEYINPUT43), .B1(new_n747_), .B2(new_n746_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n751_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n753_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n752_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(new_n698_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(G29gat), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n366_), .A2(new_n330_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n760_), .A2(new_n282_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n693_), .A2(new_n761_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n697_), .A2(G29gat), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT112), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n759_), .B1(new_n762_), .B2(new_n764_), .ZN(G1328gat));
  NAND3_X1  g564(.A1(new_n752_), .A2(new_n756_), .A3(new_n712_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(G36gat), .ZN(new_n767_));
  INV_X1    g566(.A(new_n712_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n762_), .A2(G36gat), .A3(new_n768_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT45), .Z(new_n770_));
  NAND2_X1  g569(.A1(new_n767_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT46), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n767_), .A2(KEYINPUT46), .A3(new_n770_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(G1329gat));
  NAND4_X1  g574(.A1(new_n752_), .A2(new_n756_), .A3(G43gat), .A4(new_n622_), .ZN(new_n776_));
  INV_X1    g575(.A(G43gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n777_), .B1(new_n762_), .B2(new_n661_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g579(.A(G50gat), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n469_), .A2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n693_), .A2(new_n468_), .A3(new_n761_), .ZN(new_n783_));
  AOI22_X1  g582(.A1(new_n757_), .A2(new_n782_), .B1(new_n781_), .B2(new_n783_), .ZN(G1331gat));
  NOR3_X1   g583(.A1(new_n704_), .A2(new_n705_), .A3(new_n330_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n703_), .A2(G57gat), .A3(new_n698_), .A4(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n330_), .B1(new_n368_), .B2(new_n372_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n282_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n742_), .A2(new_n397_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n787_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n705_), .B1(new_n660_), .B2(new_n692_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n792_), .A2(KEYINPUT113), .A3(new_n282_), .A4(new_n788_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n791_), .A2(new_n698_), .A3(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n795_));
  INV_X1    g594(.A(G57gat), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n794_), .A2(new_n795_), .A3(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n795_), .B1(new_n794_), .B2(new_n796_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n786_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT115), .ZN(G1332gat));
  AND2_X1   g599(.A1(new_n791_), .A2(new_n793_), .ZN(new_n801_));
  INV_X1    g600(.A(G64gat), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(new_n802_), .A3(new_n712_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n703_), .A2(new_n712_), .A3(new_n785_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(G64gat), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n805_), .A2(KEYINPUT48), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(KEYINPUT48), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n803_), .B1(new_n806_), .B2(new_n807_), .ZN(G1333gat));
  NAND3_X1  g607(.A1(new_n801_), .A2(new_n598_), .A3(new_n622_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n703_), .A2(new_n622_), .A3(new_n785_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(G71gat), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n811_), .A2(KEYINPUT49), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n811_), .A2(KEYINPUT49), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n809_), .B1(new_n812_), .B2(new_n813_), .ZN(G1334gat));
  INV_X1    g613(.A(G78gat), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n801_), .A2(new_n815_), .A3(new_n468_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n703_), .A2(new_n468_), .A3(new_n785_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(G78gat), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n818_), .A2(KEYINPUT50), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(KEYINPUT50), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n816_), .B1(new_n819_), .B2(new_n820_), .ZN(G1335gat));
  NAND3_X1  g620(.A1(new_n282_), .A2(new_n330_), .A3(new_n397_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT116), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n754_), .B2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n749_), .A2(KEYINPUT116), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(G85gat), .B1(new_n826_), .B2(new_n697_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n760_), .A2(new_n704_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n792_), .A2(new_n828_), .ZN(new_n829_));
  OR2_X1    g628(.A1(new_n697_), .A2(G85gat), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n827_), .B1(new_n829_), .B2(new_n830_), .ZN(G1336gat));
  OAI21_X1  g630(.A(G92gat), .B1(new_n826_), .B2(new_n768_), .ZN(new_n832_));
  OR2_X1    g631(.A1(new_n768_), .A2(G92gat), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n832_), .B1(new_n829_), .B2(new_n833_), .ZN(G1337gat));
  NAND3_X1  g633(.A1(new_n824_), .A2(new_n825_), .A3(new_n622_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(G99gat), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n792_), .A2(new_n622_), .A3(new_n238_), .A4(new_n828_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT51), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT51), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n836_), .A2(new_n840_), .A3(new_n837_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n841_), .ZN(G1338gat));
  NAND4_X1  g641(.A1(new_n792_), .A2(new_n239_), .A3(new_n468_), .A4(new_n828_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n822_), .A2(new_n469_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n749_), .A2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n844_), .B1(new_n846_), .B2(G106gat), .ZN(new_n847_));
  INV_X1    g646(.A(new_n845_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n844_), .B(G106gat), .C1(new_n754_), .C2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n843_), .B1(new_n847_), .B2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(KEYINPUT53), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n853_), .B(new_n843_), .C1(new_n847_), .C2(new_n850_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n854_), .ZN(G1339gat));
  NOR2_X1   g654(.A1(new_n697_), .A2(new_n661_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n657_), .A2(new_n856_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n788_), .A2(new_n704_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n860_), .B2(new_n705_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n788_), .A2(new_n397_), .A3(new_n704_), .A4(new_n858_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT118), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT118), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n373_), .A2(new_n864_), .A3(new_n397_), .A4(new_n858_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n861_), .A2(new_n863_), .A3(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT58), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n256_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n260_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT55), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n278_), .A2(new_n870_), .ZN(new_n871_));
  OAI211_X1 g670(.A(KEYINPUT55), .B(new_n274_), .C1(new_n276_), .C2(new_n277_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n869_), .A2(new_n871_), .A3(new_n872_), .ZN(new_n873_));
  AND3_X1   g672(.A1(new_n873_), .A2(KEYINPUT56), .A3(new_n266_), .ZN(new_n874_));
  AOI21_X1  g673(.A(KEYINPUT56), .B1(new_n873_), .B2(new_n266_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n874_), .A2(new_n875_), .A3(KEYINPUT121), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n873_), .A2(new_n266_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT56), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n877_), .A2(KEYINPUT121), .A3(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n378_), .B1(new_n314_), .B2(new_n333_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n377_), .A2(new_n880_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n386_), .A2(new_n378_), .A3(new_n387_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n881_), .A2(new_n882_), .A3(new_n392_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n394_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n262_), .A2(new_n278_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n266_), .B2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n879_), .A2(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n867_), .B1(new_n876_), .B2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n877_), .A2(new_n878_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n873_), .A2(KEYINPUT56), .A3(new_n266_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n890_), .A2(new_n891_), .A3(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n886_), .B1(new_n875_), .B2(KEYINPUT121), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n893_), .A2(new_n894_), .A3(KEYINPUT58), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n889_), .A2(new_n368_), .A3(new_n372_), .A4(new_n895_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n897_));
  OAI22_X1  g696(.A1(new_n395_), .A2(new_n396_), .B1(new_n885_), .B2(new_n266_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n898_), .B1(new_n890_), .B2(new_n892_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n884_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT119), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n884_), .B(KEYINPUT119), .C1(new_n279_), .C2(new_n280_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n899_), .A2(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n897_), .B1(new_n905_), .B2(new_n366_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n896_), .A2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n366_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n908_), .B1(new_n899_), .B2(new_n904_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT57), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n330_), .B1(new_n907_), .B2(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n857_), .B1(new_n866_), .B2(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(G113gat), .B1(new_n913_), .B2(new_n705_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n913_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT123), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n907_), .A2(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n911_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n896_), .A2(new_n906_), .A3(KEYINPUT123), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n917_), .A2(new_n918_), .A3(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n330_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(new_n866_), .ZN(new_n922_));
  XOR2_X1   g721(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n923_));
  NOR2_X1   g722(.A1(new_n857_), .A2(new_n923_), .ZN(new_n924_));
  AOI22_X1  g723(.A1(new_n915_), .A2(KEYINPUT59), .B1(new_n922_), .B2(new_n924_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n705_), .A2(G113gat), .ZN(new_n926_));
  XOR2_X1   g725(.A(new_n926_), .B(KEYINPUT124), .Z(new_n927_));
  AOI21_X1  g726(.A(new_n914_), .B1(new_n925_), .B2(new_n927_), .ZN(G1340gat));
  AND3_X1   g727(.A1(new_n861_), .A2(new_n863_), .A3(new_n865_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n911_), .B1(new_n907_), .B2(new_n916_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n750_), .B1(new_n930_), .B2(new_n919_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n924_), .B1(new_n929_), .B2(new_n931_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT59), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n932_), .B1(new_n933_), .B2(new_n913_), .ZN(new_n934_));
  OAI21_X1  g733(.A(G120gat), .B1(new_n934_), .B2(new_n704_), .ZN(new_n935_));
  INV_X1    g734(.A(G120gat), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n936_), .B1(new_n704_), .B2(KEYINPUT60), .ZN(new_n937_));
  OAI211_X1 g736(.A(new_n913_), .B(new_n937_), .C1(KEYINPUT60), .C2(new_n936_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n935_), .A2(new_n938_), .ZN(G1341gat));
  OAI21_X1  g738(.A(G127gat), .B1(new_n934_), .B2(new_n330_), .ZN(new_n940_));
  OR3_X1    g739(.A1(new_n915_), .A2(G127gat), .A3(new_n330_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(G1342gat));
  NAND2_X1  g741(.A1(new_n368_), .A2(new_n372_), .ZN(new_n943_));
  OAI21_X1  g742(.A(G134gat), .B1(new_n934_), .B2(new_n943_), .ZN(new_n944_));
  OR3_X1    g743(.A1(new_n915_), .A2(G134gat), .A3(new_n908_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(G1343gat));
  NAND2_X1  g745(.A1(new_n866_), .A2(new_n912_), .ZN(new_n947_));
  NOR4_X1   g746(.A1(new_n712_), .A2(new_n697_), .A3(new_n469_), .A4(new_n622_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n947_), .A2(new_n948_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n949_), .A2(new_n397_), .ZN(new_n950_));
  INV_X1    g749(.A(G141gat), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n950_), .B(new_n951_), .ZN(G1344gat));
  NOR2_X1   g751(.A1(new_n949_), .A2(new_n704_), .ZN(new_n953_));
  INV_X1    g752(.A(G148gat), .ZN(new_n954_));
  XNOR2_X1  g753(.A(new_n953_), .B(new_n954_), .ZN(G1345gat));
  NOR2_X1   g754(.A1(new_n949_), .A2(new_n330_), .ZN(new_n956_));
  XNOR2_X1  g755(.A(KEYINPUT61), .B(G155gat), .ZN(new_n957_));
  INV_X1    g756(.A(new_n957_), .ZN(new_n958_));
  XNOR2_X1  g757(.A(new_n956_), .B(new_n958_), .ZN(G1346gat));
  AND2_X1   g758(.A1(new_n947_), .A2(new_n948_), .ZN(new_n960_));
  AOI21_X1  g759(.A(G162gat), .B1(new_n960_), .B2(new_n366_), .ZN(new_n961_));
  AND3_X1   g760(.A1(new_n733_), .A2(G162gat), .A3(new_n743_), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n961_), .B1(new_n960_), .B2(new_n962_), .ZN(G1347gat));
  NOR2_X1   g762(.A1(new_n768_), .A2(new_n650_), .ZN(new_n964_));
  INV_X1    g763(.A(new_n964_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n965_), .A2(new_n468_), .ZN(new_n966_));
  OAI211_X1 g765(.A(new_n705_), .B(new_n966_), .C1(new_n929_), .C2(new_n931_), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n480_), .B1(KEYINPUT125), .B2(KEYINPUT62), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n967_), .A2(new_n968_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n969_), .A2(new_n970_), .ZN(new_n971_));
  OAI211_X1 g770(.A(new_n967_), .B(new_n968_), .C1(KEYINPUT125), .C2(KEYINPUT62), .ZN(new_n972_));
  INV_X1    g771(.A(new_n966_), .ZN(new_n973_));
  AOI21_X1  g772(.A(new_n973_), .B1(new_n921_), .B2(new_n866_), .ZN(new_n974_));
  NAND3_X1  g773(.A1(new_n974_), .A2(new_n534_), .A3(new_n705_), .ZN(new_n975_));
  NAND3_X1  g774(.A1(new_n971_), .A2(new_n972_), .A3(new_n975_), .ZN(G1348gat));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n977_));
  AOI21_X1  g776(.A(G176gat), .B1(new_n974_), .B2(new_n282_), .ZN(new_n978_));
  AOI21_X1  g777(.A(new_n468_), .B1(new_n866_), .B2(new_n912_), .ZN(new_n979_));
  NOR3_X1   g778(.A1(new_n965_), .A2(new_n704_), .A3(new_n482_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n979_), .A2(new_n980_), .ZN(new_n981_));
  INV_X1    g780(.A(new_n981_), .ZN(new_n982_));
  OAI21_X1  g781(.A(new_n977_), .B1(new_n978_), .B2(new_n982_), .ZN(new_n983_));
  OAI211_X1 g782(.A(new_n282_), .B(new_n966_), .C1(new_n929_), .C2(new_n931_), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n984_), .A2(new_n482_), .ZN(new_n985_));
  NAND3_X1  g784(.A1(new_n985_), .A2(KEYINPUT126), .A3(new_n981_), .ZN(new_n986_));
  NAND2_X1  g785(.A1(new_n983_), .A2(new_n986_), .ZN(G1349gat));
  NAND3_X1  g786(.A1(new_n979_), .A2(new_n750_), .A3(new_n964_), .ZN(new_n988_));
  INV_X1    g787(.A(G183gat), .ZN(new_n989_));
  NOR2_X1   g788(.A1(new_n330_), .A2(new_n517_), .ZN(new_n990_));
  AOI22_X1  g789(.A1(new_n988_), .A2(new_n989_), .B1(new_n974_), .B2(new_n990_), .ZN(G1350gat));
  NAND2_X1  g790(.A1(new_n974_), .A2(new_n747_), .ZN(new_n992_));
  NAND2_X1  g791(.A1(new_n992_), .A2(G190gat), .ZN(new_n993_));
  NAND3_X1  g792(.A1(new_n974_), .A2(new_n521_), .A3(new_n366_), .ZN(new_n994_));
  NAND2_X1  g793(.A1(new_n993_), .A2(new_n994_), .ZN(G1351gat));
  NOR3_X1   g794(.A1(new_n768_), .A2(new_n690_), .A3(new_n622_), .ZN(new_n996_));
  NAND2_X1  g795(.A1(new_n947_), .A2(new_n996_), .ZN(new_n997_));
  NOR2_X1   g796(.A1(new_n997_), .A2(new_n397_), .ZN(new_n998_));
  INV_X1    g797(.A(G197gat), .ZN(new_n999_));
  XNOR2_X1  g798(.A(new_n998_), .B(new_n999_), .ZN(G1352gat));
  NOR2_X1   g799(.A1(new_n997_), .A2(new_n704_), .ZN(new_n1001_));
  INV_X1    g800(.A(G204gat), .ZN(new_n1002_));
  XNOR2_X1  g801(.A(new_n1001_), .B(new_n1002_), .ZN(G1353gat));
  OR2_X1    g802(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1004_));
  AND2_X1   g803(.A1(new_n947_), .A2(new_n996_), .ZN(new_n1005_));
  AOI21_X1  g804(.A(new_n1004_), .B1(new_n1005_), .B2(new_n750_), .ZN(new_n1006_));
  NOR2_X1   g805(.A1(new_n997_), .A2(new_n330_), .ZN(new_n1007_));
  XOR2_X1   g806(.A(KEYINPUT63), .B(G211gat), .Z(new_n1008_));
  AOI21_X1  g807(.A(new_n1006_), .B1(new_n1007_), .B2(new_n1008_), .ZN(G1354gat));
  INV_X1    g808(.A(G218gat), .ZN(new_n1010_));
  NAND3_X1  g809(.A1(new_n1005_), .A2(new_n1010_), .A3(new_n366_), .ZN(new_n1011_));
  OAI21_X1  g810(.A(G218gat), .B1(new_n997_), .B2(new_n943_), .ZN(new_n1012_));
  NAND2_X1  g811(.A1(new_n1011_), .A2(new_n1012_), .ZN(G1355gat));
endmodule


