//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 0 1 0 1 0 1 0 0 0 0 0 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 0 0 0 1 1 1 1 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n872_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n904_, new_n905_, new_n907_,
    new_n908_, new_n910_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT23), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND3_X1  g003(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n205_));
  OAI211_X1 g004(.A(new_n204_), .B(new_n205_), .C1(G183gat), .C2(G190gat), .ZN(new_n206_));
  INV_X1    g005(.A(G176gat), .ZN(new_n207_));
  AND2_X1   g006(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n207_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n206_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  AND2_X1   g011(.A1(new_n204_), .A2(new_n205_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT78), .ZN(new_n214_));
  INV_X1    g013(.A(G169gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n215_), .A3(new_n207_), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT78), .B1(G169gat), .B2(G176gat), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n216_), .A2(KEYINPUT24), .A3(new_n217_), .A4(new_n211_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n217_), .ZN(new_n219_));
  NOR3_X1   g018(.A1(KEYINPUT78), .A2(G169gat), .A3(G176gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n213_), .B(new_n218_), .C1(new_n221_), .C2(KEYINPUT24), .ZN(new_n222_));
  INV_X1    g021(.A(G190gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT26), .B1(new_n223_), .B2(KEYINPUT77), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT77), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT26), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(G190gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n224_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(G183gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(KEYINPUT76), .A3(KEYINPUT25), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(KEYINPUT25), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT25), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(G183gat), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT76), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n231_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n228_), .B1(new_n230_), .B2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n212_), .B1(new_n222_), .B2(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(G197gat), .B(G204gat), .Z(new_n238_));
  XNOR2_X1  g037(.A(G211gat), .B(G218gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT88), .ZN(new_n240_));
  INV_X1    g039(.A(G197gat), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n240_), .B1(new_n241_), .B2(G204gat), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n238_), .A2(KEYINPUT21), .A3(new_n239_), .A4(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G197gat), .B(G204gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(KEYINPUT21), .ZN(new_n245_));
  AND2_X1   g044(.A1(G211gat), .A2(G218gat), .ZN(new_n246_));
  NOR2_X1   g045(.A1(G211gat), .A2(G218gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n244_), .B1(new_n245_), .B2(new_n248_), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n239_), .A2(KEYINPUT21), .ZN(new_n250_));
  AND3_X1   g049(.A1(new_n243_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n237_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT95), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G226gat), .A2(G233gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT19), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n216_), .A2(new_n217_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT91), .B(KEYINPUT24), .ZN(new_n259_));
  INV_X1    g058(.A(new_n211_), .ZN(new_n260_));
  OR3_X1    g059(.A1(new_n258_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n259_), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n231_), .A2(new_n233_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT26), .B(G190gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n261_), .A2(new_n262_), .A3(new_n213_), .A4(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n260_), .A2(KEYINPUT92), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT92), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n211_), .A2(new_n268_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n206_), .A2(new_n267_), .A3(new_n210_), .A4(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT93), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n270_), .A2(new_n271_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n266_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n274_), .A2(new_n251_), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n254_), .A2(KEYINPUT20), .A3(new_n257_), .A4(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT20), .B1(new_n237_), .B2(new_n251_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT90), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(new_n251_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT90), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n280_), .B(KEYINPUT20), .C1(new_n237_), .C2(new_n251_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n278_), .A2(new_n279_), .A3(new_n281_), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n282_), .A2(KEYINPUT94), .A3(new_n256_), .ZN(new_n283_));
  AOI21_X1  g082(.A(KEYINPUT94), .B1(new_n282_), .B2(new_n256_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n276_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(G8gat), .B(G36gat), .Z(new_n286_));
  XNOR2_X1  g085(.A(G64gat), .B(G92gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n288_), .B(new_n289_), .Z(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n285_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT97), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n290_), .B(new_n276_), .C1(new_n283_), .C2(new_n284_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n292_), .A2(new_n293_), .A3(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT27), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n283_), .A2(new_n284_), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n297_), .A2(KEYINPUT97), .A3(new_n290_), .A4(new_n276_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n295_), .A2(new_n296_), .A3(new_n298_), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n294_), .A2(KEYINPUT100), .ZN(new_n300_));
  INV_X1    g099(.A(new_n251_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(new_n266_), .A3(new_n270_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n254_), .A2(KEYINPUT20), .A3(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n256_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n304_), .B1(new_n256_), .B2(new_n282_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n296_), .B1(new_n305_), .B2(new_n291_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n294_), .A2(KEYINPUT100), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n300_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT83), .B(G113gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(G120gat), .ZN(new_n310_));
  XOR2_X1   g109(.A(G127gat), .B(G134gat), .Z(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  OR2_X1    g111(.A1(G141gat), .A2(G148gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G141gat), .A2(G148gat), .ZN(new_n314_));
  NOR2_X1   g113(.A1(G155gat), .A2(G162gat), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT85), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n317_), .B1(KEYINPUT1), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(KEYINPUT1), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT86), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n313_), .B(new_n314_), .C1(new_n319_), .C2(new_n321_), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n313_), .A2(KEYINPUT3), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n313_), .A2(KEYINPUT3), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT2), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n314_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n323_), .A2(new_n324_), .A3(new_n326_), .A4(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n328_), .A2(new_n318_), .A3(new_n317_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n312_), .A2(new_n322_), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n322_), .A2(new_n329_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n311_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n310_), .B(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n330_), .A2(new_n334_), .A3(KEYINPUT4), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G225gat), .A2(G233gat), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT4), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n331_), .A2(new_n333_), .A3(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n335_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT98), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n330_), .A2(new_n334_), .A3(new_n341_), .A4(new_n336_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n330_), .A2(new_n334_), .A3(new_n336_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT98), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n340_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT0), .B(G57gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(G85gat), .ZN(new_n347_));
  XOR2_X1   g146(.A(G1gat), .B(G29gat), .Z(new_n348_));
  XOR2_X1   g147(.A(new_n347_), .B(new_n348_), .Z(new_n349_));
  NAND2_X1  g148(.A1(new_n345_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n349_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n340_), .A2(new_n344_), .A3(new_n351_), .A4(new_n342_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n301_), .B1(new_n331_), .B2(KEYINPUT29), .ZN(new_n355_));
  INV_X1    g154(.A(G233gat), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT87), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n357_), .A2(G228gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(G228gat), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n356_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT28), .ZN(new_n361_));
  XOR2_X1   g160(.A(G22gat), .B(G50gat), .Z(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n355_), .B(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n331_), .A2(KEYINPUT29), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G78gat), .B(G106gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT89), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n365_), .B(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n364_), .B(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n299_), .A2(new_n308_), .A3(new_n354_), .A4(new_n370_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n290_), .A2(KEYINPUT32), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n285_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n305_), .A2(new_n372_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(new_n353_), .A3(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT33), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n352_), .A2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n330_), .A2(new_n334_), .A3(new_n337_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n335_), .A2(new_n339_), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n349_), .B(new_n379_), .C1(new_n380_), .C2(new_n337_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n378_), .A2(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n382_), .B1(new_n295_), .B2(new_n298_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n352_), .A2(new_n377_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT99), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n376_), .B1(new_n383_), .B2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n371_), .B1(new_n386_), .B2(new_n370_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G227gat), .A2(G233gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT80), .ZN(new_n389_));
  INV_X1    g188(.A(G71gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(G99gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G15gat), .B(G43gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT81), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n392_), .B(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n237_), .A2(KEYINPUT79), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT79), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n397_), .B(new_n212_), .C1(new_n222_), .C2(new_n236_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT30), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT82), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n396_), .A2(KEYINPUT30), .A3(new_n398_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n401_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT84), .ZN(new_n405_));
  AND3_X1   g204(.A1(new_n395_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n405_), .B1(new_n395_), .B2(new_n404_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n333_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n395_), .A2(new_n404_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT84), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n395_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(new_n312_), .A3(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n402_), .B1(new_n401_), .B2(new_n403_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT31), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n408_), .A2(new_n412_), .A3(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n414_), .B1(new_n408_), .B2(new_n412_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n299_), .A2(new_n308_), .ZN(new_n419_));
  NOR3_X1   g218(.A1(new_n415_), .A2(new_n416_), .A3(new_n353_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n419_), .A2(KEYINPUT101), .A3(new_n369_), .A4(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT101), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n417_), .A2(new_n354_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n299_), .A2(new_n369_), .A3(new_n308_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n422_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  AOI22_X1  g224(.A1(new_n387_), .A2(new_n418_), .B1(new_n421_), .B2(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(G85gat), .A2(G92gat), .ZN(new_n427_));
  AND2_X1   g226(.A1(G85gat), .A2(G92gat), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n427_), .B1(new_n428_), .B2(KEYINPUT9), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT65), .ZN(new_n430_));
  INV_X1    g229(.A(G92gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(G85gat), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT66), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT9), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n434_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n435_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n429_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT67), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT67), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n441_), .B(new_n429_), .C1(new_n437_), .C2(new_n438_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G99gat), .A2(G106gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT6), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT10), .B(G99gat), .ZN(new_n446_));
  OR3_X1    g245(.A1(new_n446_), .A2(KEYINPUT64), .A3(G106gat), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT64), .B1(new_n446_), .B2(G106gat), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n445_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n440_), .A2(new_n442_), .A3(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n451_));
  OR3_X1    g250(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n444_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n428_), .A2(new_n427_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT8), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT8), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n453_), .A2(new_n457_), .A3(new_n454_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n450_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G57gat), .B(G64gat), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n461_), .A2(KEYINPUT11), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(KEYINPUT11), .ZN(new_n463_));
  XOR2_X1   g262(.A(G71gat), .B(G78gat), .Z(new_n464_));
  NAND3_X1  g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  OR2_X1    g264(.A1(new_n463_), .A2(new_n464_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n460_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT12), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n450_), .A2(new_n459_), .A3(new_n467_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G230gat), .A2(G233gat), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n460_), .A2(KEYINPUT12), .A3(new_n468_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n471_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n469_), .A2(new_n472_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n473_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n476_), .A2(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(G120gat), .B(G148gat), .Z(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(G204gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT5), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(new_n207_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT68), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n480_), .A2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n476_), .A2(new_n479_), .A3(new_n484_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT13), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n486_), .A2(KEYINPUT13), .A3(new_n487_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(G15gat), .B(G22gat), .Z(new_n494_));
  NAND2_X1  g293(.A1(G1gat), .A2(G8gat), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n494_), .B1(KEYINPUT14), .B2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT72), .ZN(new_n497_));
  XOR2_X1   g296(.A(G1gat), .B(G8gat), .Z(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT72), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n496_), .B(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n498_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n499_), .A2(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(KEYINPUT69), .B(G29gat), .Z(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(G36gat), .ZN(new_n506_));
  XOR2_X1   g305(.A(G43gat), .B(G50gat), .Z(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT69), .B(G29gat), .ZN(new_n508_));
  INV_X1    g307(.A(G36gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n506_), .A2(new_n507_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n507_), .B1(new_n506_), .B2(new_n510_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n504_), .A2(new_n514_), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n499_), .B(new_n503_), .C1(new_n512_), .C2(new_n513_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G229gat), .A2(G233gat), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT15), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n521_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n506_), .A2(new_n510_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n507_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n525_), .A2(KEYINPUT15), .A3(new_n511_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n522_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n504_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n529_), .A2(new_n518_), .A3(new_n516_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n520_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G113gat), .B(G141gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(new_n215_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(new_n241_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n531_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n534_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n520_), .A2(new_n530_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n535_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n493_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n426_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G190gat), .B(G218gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(G134gat), .ZN(new_n544_));
  INV_X1    g343(.A(G162gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n460_), .A2(new_n514_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n527_), .B1(new_n459_), .B2(new_n450_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G232gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT34), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n460_), .A2(new_n528_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT70), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n550_), .A2(KEYINPUT35), .A3(new_n552_), .A4(new_n555_), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n552_), .A2(KEYINPUT35), .ZN(new_n557_));
  OAI211_X1 g356(.A(KEYINPUT35), .B(new_n552_), .C1(new_n549_), .C2(KEYINPUT70), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n553_), .B1(new_n514_), .B2(new_n460_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n556_), .A2(new_n557_), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT71), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n547_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT36), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n563_), .A2(new_n564_), .B1(new_n561_), .B2(new_n547_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n561_), .A2(new_n562_), .ZN(new_n566_));
  OAI21_X1  g365(.A(KEYINPUT36), .B1(new_n566_), .B2(new_n547_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n565_), .A2(new_n567_), .A3(KEYINPUT37), .ZN(new_n568_));
  AOI21_X1  g367(.A(KEYINPUT37), .B1(new_n565_), .B2(new_n567_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(G231gat), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n571_), .A2(new_n356_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n499_), .A2(new_n503_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n467_), .B(KEYINPUT73), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n573_), .B1(new_n499_), .B2(new_n503_), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n575_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n576_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n504_), .A2(new_n572_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n579_), .B1(new_n580_), .B2(new_n574_), .ZN(new_n581_));
  XOR2_X1   g380(.A(G127gat), .B(G155gat), .Z(new_n582_));
  XNOR2_X1  g381(.A(G183gat), .B(G211gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT17), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n586_), .A2(new_n587_), .ZN(new_n589_));
  NOR4_X1   g388(.A1(new_n578_), .A2(new_n581_), .A3(new_n588_), .A4(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n588_), .B1(new_n578_), .B2(new_n581_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n591_), .A2(KEYINPUT75), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(KEYINPUT75), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n590_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n570_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n542_), .A2(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n597_), .B(KEYINPUT102), .Z(new_n598_));
  INV_X1    g397(.A(G1gat), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n598_), .A2(new_n599_), .A3(new_n353_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT38), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n563_), .A2(new_n564_), .ZN(new_n602_));
  AOI211_X1 g401(.A(KEYINPUT36), .B(new_n547_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n561_), .A2(new_n547_), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n602_), .A2(new_n603_), .A3(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT103), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(new_n595_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n542_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT104), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(G1gat), .B1(new_n610_), .B2(new_n354_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT105), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n601_), .A2(new_n612_), .ZN(G1324gat));
  INV_X1    g412(.A(KEYINPUT39), .ZN(new_n614_));
  OAI21_X1  g413(.A(G8gat), .B1(new_n608_), .B2(new_n419_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT106), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n615_), .A2(KEYINPUT106), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n614_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n618_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(KEYINPUT39), .A3(new_n616_), .ZN(new_n621_));
  INV_X1    g420(.A(G8gat), .ZN(new_n622_));
  INV_X1    g421(.A(new_n419_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n598_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n619_), .A2(new_n621_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT40), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n619_), .A2(new_n621_), .A3(new_n624_), .A4(KEYINPUT40), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(G1325gat));
  OAI21_X1  g428(.A(G15gat), .B1(new_n610_), .B2(new_n418_), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n630_), .B(KEYINPUT41), .Z(new_n631_));
  INV_X1    g430(.A(G15gat), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n598_), .A2(new_n632_), .A3(new_n417_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(G1326gat));
  NOR2_X1   g433(.A1(new_n369_), .A2(G22gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT108), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n598_), .A2(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(G22gat), .B1(new_n610_), .B2(new_n369_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT107), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT107), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n640_), .B(G22gat), .C1(new_n610_), .C2(new_n369_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n639_), .A2(KEYINPUT42), .A3(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(KEYINPUT42), .B1(new_n639_), .B2(new_n641_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n637_), .B1(new_n642_), .B2(new_n643_), .ZN(G1327gat));
  NOR2_X1   g443(.A1(new_n605_), .A2(new_n594_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n542_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(G29gat), .B1(new_n647_), .B2(new_n353_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n565_), .A2(new_n567_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT37), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n565_), .A2(new_n567_), .A3(KEYINPUT37), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  OAI21_X1  g452(.A(KEYINPUT43), .B1(new_n426_), .B2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n421_), .A2(new_n425_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n295_), .A2(new_n298_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n382_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n656_), .A2(new_n657_), .A3(new_n385_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n370_), .B1(new_n658_), .B2(new_n375_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n371_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n418_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n655_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT43), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n662_), .A2(new_n663_), .A3(new_n570_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n654_), .A2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(new_n540_), .A3(new_n595_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n665_), .A2(KEYINPUT44), .A3(new_n540_), .A4(new_n595_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n670_), .A2(new_n353_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n648_), .B1(new_n671_), .B2(G29gat), .ZN(G1328gat));
  NAND3_X1  g471(.A1(new_n668_), .A2(new_n623_), .A3(new_n669_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(G36gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n647_), .A2(new_n509_), .A3(new_n623_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT45), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT46), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n677_), .B(new_n678_), .ZN(G1329gat));
  INV_X1    g478(.A(KEYINPUT47), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n668_), .A2(G43gat), .A3(new_n417_), .A4(new_n669_), .ZN(new_n681_));
  INV_X1    g480(.A(G43gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n682_), .B1(new_n646_), .B2(new_n418_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT109), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  OAI211_X1 g484(.A(KEYINPUT109), .B(new_n682_), .C1(new_n646_), .C2(new_n418_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT110), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n681_), .A2(new_n687_), .A3(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n681_), .B2(new_n687_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n680_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n681_), .A2(new_n687_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT110), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n681_), .A2(new_n687_), .A3(new_n688_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(KEYINPUT47), .A3(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n691_), .A2(new_n695_), .ZN(G1330gat));
  AOI21_X1  g495(.A(G50gat), .B1(new_n647_), .B2(new_n370_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n370_), .A2(G50gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n670_), .B2(new_n698_), .ZN(G1331gat));
  NOR2_X1   g498(.A1(new_n426_), .A2(new_n538_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT111), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n701_), .A2(new_n492_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n702_), .A2(new_n596_), .ZN(new_n703_));
  AOI21_X1  g502(.A(G57gat), .B1(new_n703_), .B2(new_n353_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n700_), .A2(new_n493_), .A3(new_n607_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n705_), .A2(new_n354_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n704_), .B1(G57gat), .B2(new_n706_), .ZN(G1332gat));
  INV_X1    g506(.A(G64gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n703_), .A2(new_n708_), .A3(new_n623_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G64gat), .B1(new_n705_), .B2(new_n419_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT48), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n711_), .ZN(G1333gat));
  NAND3_X1  g511(.A1(new_n703_), .A2(new_n390_), .A3(new_n417_), .ZN(new_n713_));
  OAI21_X1  g512(.A(G71gat), .B1(new_n705_), .B2(new_n418_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT49), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1334gat));
  INV_X1    g515(.A(G78gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n703_), .A2(new_n717_), .A3(new_n370_), .ZN(new_n718_));
  OAI21_X1  g517(.A(G78gat), .B1(new_n705_), .B2(new_n369_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT50), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1335gat));
  NAND2_X1  g520(.A1(new_n702_), .A2(new_n645_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(G85gat), .B1(new_n723_), .B2(new_n353_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n492_), .A2(new_n538_), .A3(new_n594_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n665_), .A2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT112), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n727_), .A2(new_n354_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n724_), .B1(G85gat), .B2(new_n728_), .ZN(G1336gat));
  AOI21_X1  g528(.A(G92gat), .B1(new_n723_), .B2(new_n623_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n432_), .A2(new_n433_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n727_), .A2(new_n419_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n730_), .B1(new_n731_), .B2(new_n732_), .ZN(G1337gat));
  OR2_X1    g532(.A1(new_n418_), .A2(new_n446_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n726_), .A2(new_n417_), .ZN(new_n735_));
  INV_X1    g534(.A(G99gat), .ZN(new_n736_));
  OAI22_X1  g535(.A1(new_n722_), .A2(new_n734_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT51), .ZN(G1338gat));
  AOI21_X1  g537(.A(new_n663_), .B1(new_n662_), .B2(new_n570_), .ZN(new_n739_));
  AOI211_X1 g538(.A(KEYINPUT43), .B(new_n653_), .C1(new_n655_), .C2(new_n661_), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n370_), .B(new_n725_), .C1(new_n739_), .C2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT113), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT113), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n665_), .A2(new_n743_), .A3(new_n370_), .A4(new_n725_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n742_), .A2(G106gat), .A3(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT52), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT52), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n742_), .A2(new_n747_), .A3(new_n744_), .A4(G106gat), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n369_), .A2(G106gat), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n702_), .A2(new_n645_), .A3(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT53), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT53), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n749_), .A2(new_n754_), .A3(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1339gat));
  INV_X1    g555(.A(G113gat), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n419_), .A2(new_n369_), .A3(new_n417_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n758_), .A2(new_n354_), .ZN(new_n759_));
  AOI21_X1  g558(.A(KEYINPUT59), .B1(new_n759_), .B2(KEYINPUT120), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n760_), .B1(KEYINPUT120), .B2(new_n759_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n538_), .A2(new_n487_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n471_), .A2(new_n474_), .A3(KEYINPUT55), .A4(new_n475_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT116), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(KEYINPUT12), .B1(new_n460_), .B2(new_n468_), .ZN(new_n766_));
  AOI211_X1 g565(.A(new_n470_), .B(new_n467_), .C1(new_n450_), .C2(new_n459_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n768_), .A2(KEYINPUT116), .A3(KEYINPUT55), .A4(new_n474_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n765_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n472_), .A2(new_n473_), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n766_), .A2(new_n767_), .A3(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n472_), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n766_), .A2(new_n767_), .A3(new_n773_), .ZN(new_n774_));
  OAI22_X1  g573(.A1(KEYINPUT55), .A2(new_n772_), .B1(new_n774_), .B2(new_n473_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n485_), .B1(new_n770_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT56), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT55), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n476_), .A2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n471_), .A2(new_n472_), .A3(new_n475_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n478_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n765_), .A2(new_n780_), .A3(new_n769_), .A4(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n783_), .A2(KEYINPUT56), .A3(new_n485_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n762_), .B1(new_n778_), .B2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n517_), .A2(new_n518_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n529_), .A2(new_n519_), .A3(new_n516_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n786_), .A2(new_n534_), .A3(new_n787_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n788_), .A2(new_n537_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n488_), .A2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n605_), .B1(new_n785_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT117), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  XOR2_X1   g592(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n794_));
  OAI211_X1 g593(.A(new_n605_), .B(KEYINPUT117), .C1(new_n785_), .C2(new_n790_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n793_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n783_), .A2(KEYINPUT56), .A3(new_n485_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT56), .B1(new_n783_), .B2(new_n485_), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n487_), .B(new_n789_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT58), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n778_), .A2(new_n784_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n802_), .A2(KEYINPUT58), .A3(new_n487_), .A4(new_n789_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n570_), .A2(new_n801_), .A3(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n796_), .A2(KEYINPUT121), .A3(new_n804_), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n605_), .B(KEYINPUT57), .C1(new_n785_), .C2(new_n790_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT121), .B1(new_n796_), .B2(new_n804_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n595_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n492_), .A2(new_n810_), .A3(new_n539_), .A4(new_n594_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n594_), .A2(new_n490_), .A3(new_n539_), .A4(new_n491_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT114), .ZN(new_n813_));
  AOI22_X1  g612(.A1(new_n651_), .A2(new_n652_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT115), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n811_), .A2(new_n813_), .ZN(new_n818_));
  OAI21_X1  g617(.A(KEYINPUT54), .B1(new_n818_), .B2(new_n570_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT115), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n814_), .A2(new_n820_), .A3(new_n815_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n817_), .A2(new_n819_), .A3(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n761_), .B1(new_n809_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT59), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT119), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n801_), .A2(new_n803_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(new_n653_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n570_), .A2(KEYINPUT119), .A3(new_n801_), .A4(new_n803_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n796_), .A2(new_n827_), .A3(new_n806_), .A4(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n595_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n822_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n824_), .B1(new_n831_), .B2(new_n759_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n823_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n757_), .B1(new_n833_), .B2(new_n538_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n831_), .A2(new_n759_), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n835_), .A2(G113gat), .A3(new_n539_), .ZN(new_n836_));
  OAI21_X1  g635(.A(KEYINPUT122), .B1(new_n834_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT122), .ZN(new_n838_));
  INV_X1    g637(.A(new_n836_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n823_), .A2(new_n832_), .A3(new_n539_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n838_), .B(new_n839_), .C1(new_n840_), .C2(new_n757_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n837_), .A2(new_n841_), .ZN(G1340gat));
  INV_X1    g641(.A(G120gat), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n843_), .B1(new_n833_), .B2(new_n493_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n835_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT60), .ZN(new_n846_));
  AOI21_X1  g645(.A(G120gat), .B1(new_n493_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n845_), .B(new_n848_), .C1(KEYINPUT60), .C2(new_n843_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(KEYINPUT123), .B1(new_n844_), .B2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT123), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n823_), .A2(new_n832_), .A3(new_n492_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n852_), .B(new_n849_), .C1(new_n853_), .C2(new_n843_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n851_), .A2(new_n854_), .ZN(G1341gat));
  AND3_X1   g654(.A1(new_n833_), .A2(G127gat), .A3(new_n594_), .ZN(new_n856_));
  AOI21_X1  g655(.A(G127gat), .B1(new_n845_), .B2(new_n594_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(G1342gat));
  AOI21_X1  g657(.A(G134gat), .B1(new_n845_), .B2(new_n606_), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n833_), .A2(G134gat), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n859_), .B1(new_n860_), .B2(new_n570_), .ZN(G1343gat));
  NOR4_X1   g660(.A1(new_n818_), .A2(new_n570_), .A3(KEYINPUT115), .A4(KEYINPUT54), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n820_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  AOI22_X1  g663(.A1(new_n864_), .A2(new_n819_), .B1(new_n829_), .B2(new_n595_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n865_), .A2(new_n369_), .A3(new_n417_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n866_), .A2(new_n353_), .A3(new_n419_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(new_n539_), .ZN(new_n868_));
  XOR2_X1   g667(.A(KEYINPUT124), .B(G141gat), .Z(new_n869_));
  XNOR2_X1  g668(.A(new_n868_), .B(new_n869_), .ZN(G1344gat));
  NOR2_X1   g669(.A1(new_n867_), .A2(new_n492_), .ZN(new_n871_));
  INV_X1    g670(.A(G148gat), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n871_), .B(new_n872_), .ZN(G1345gat));
  NOR2_X1   g672(.A1(new_n867_), .A2(new_n595_), .ZN(new_n874_));
  XOR2_X1   g673(.A(KEYINPUT61), .B(G155gat), .Z(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1346gat));
  NOR3_X1   g675(.A1(new_n867_), .A2(new_n545_), .A3(new_n653_), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n866_), .A2(new_n353_), .A3(new_n419_), .A4(new_n606_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(new_n545_), .B2(new_n878_), .ZN(G1347gat));
  AOI21_X1  g678(.A(new_n370_), .B1(new_n809_), .B2(new_n822_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n419_), .A2(new_n353_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n417_), .ZN(new_n882_));
  XOR2_X1   g681(.A(new_n882_), .B(KEYINPUT125), .Z(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n880_), .A2(new_n538_), .A3(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(G169gat), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT62), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n880_), .A2(new_n884_), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n889_), .B(new_n538_), .C1(new_n209_), .C2(new_n208_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n885_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n888_), .A2(new_n890_), .A3(new_n891_), .ZN(G1348gat));
  AOI21_X1  g691(.A(G176gat), .B1(new_n889_), .B2(new_n493_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n865_), .A2(new_n370_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n883_), .A2(new_n207_), .A3(new_n492_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n894_), .B2(new_n895_), .ZN(G1349gat));
  INV_X1    g695(.A(KEYINPUT126), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n883_), .A2(new_n263_), .A3(new_n595_), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n880_), .A2(new_n897_), .A3(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n897_), .B1(new_n880_), .B2(new_n898_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n883_), .A2(new_n595_), .ZN(new_n901_));
  AOI21_X1  g700(.A(G183gat), .B1(new_n894_), .B2(new_n901_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n899_), .A2(new_n900_), .A3(new_n902_), .ZN(G1350gat));
  NAND3_X1  g702(.A1(new_n889_), .A2(new_n264_), .A3(new_n606_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n889_), .A2(new_n570_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n905_), .B2(new_n223_), .ZN(G1351gat));
  NAND2_X1  g705(.A1(new_n866_), .A2(new_n881_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(new_n539_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(new_n241_), .ZN(G1352gat));
  NAND3_X1  g708(.A1(new_n866_), .A2(new_n493_), .A3(new_n881_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(G204gat), .ZN(G1353gat));
  XNOR2_X1  g710(.A(KEYINPUT63), .B(G211gat), .ZN(new_n912_));
  OR2_X1    g711(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n866_), .A2(new_n594_), .A3(new_n881_), .ZN(new_n914_));
  MUX2_X1   g713(.A(new_n912_), .B(new_n913_), .S(new_n914_), .Z(G1354gat));
  NAND3_X1  g714(.A1(new_n866_), .A2(new_n606_), .A3(new_n881_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(KEYINPUT127), .ZN(new_n917_));
  INV_X1    g716(.A(G218gat), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT127), .ZN(new_n919_));
  NAND4_X1  g718(.A1(new_n866_), .A2(new_n919_), .A3(new_n606_), .A4(new_n881_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n917_), .A2(new_n918_), .A3(new_n920_), .ZN(new_n921_));
  NAND4_X1  g720(.A1(new_n866_), .A2(G218gat), .A3(new_n570_), .A4(new_n881_), .ZN(new_n922_));
  AND2_X1   g721(.A1(new_n921_), .A2(new_n922_), .ZN(G1355gat));
endmodule


