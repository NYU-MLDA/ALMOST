//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1 0 0 1 1 0 0 1 1 1 1 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n922_, new_n923_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_;
  INV_X1    g000(.A(G197gat), .ZN(new_n202_));
  INV_X1    g001(.A(G204gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G197gat), .A2(G204gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n204_), .A2(KEYINPUT21), .A3(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT83), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  OR2_X1    g007(.A1(KEYINPUT84), .A2(KEYINPUT21), .ZN(new_n209_));
  NAND2_X1  g008(.A1(KEYINPUT84), .A2(KEYINPUT21), .ZN(new_n210_));
  INV_X1    g009(.A(new_n205_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G197gat), .A2(G204gat), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n209_), .B(new_n210_), .C1(new_n211_), .C2(new_n212_), .ZN(new_n213_));
  NAND4_X1  g012(.A1(new_n204_), .A2(KEYINPUT83), .A3(KEYINPUT21), .A4(new_n205_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G211gat), .B(G218gat), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n208_), .A2(new_n213_), .A3(new_n214_), .A4(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT85), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  XOR2_X1   g017(.A(G211gat), .B(G218gat), .Z(new_n219_));
  NAND2_X1  g018(.A1(new_n204_), .A2(new_n205_), .ZN(new_n220_));
  XOR2_X1   g019(.A(KEYINPUT84), .B(KEYINPUT21), .Z(new_n221_));
  AOI21_X1  g020(.A(new_n219_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n222_), .A2(KEYINPUT85), .A3(new_n214_), .A4(new_n208_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n218_), .A2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n206_), .A2(new_n215_), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n225_), .A2(KEYINPUT86), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(KEYINPUT86), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n224_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(G228gat), .ZN(new_n230_));
  INV_X1    g029(.A(G233gat), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT29), .ZN(new_n232_));
  OR2_X1    g031(.A1(G155gat), .A2(G162gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G155gat), .A2(G162gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(G141gat), .A2(G148gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT3), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G141gat), .A2(G148gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT2), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n235_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT82), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n233_), .B1(KEYINPUT1), .B2(new_n234_), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n234_), .A2(KEYINPUT81), .A3(KEYINPUT1), .ZN(new_n243_));
  AOI21_X1  g042(.A(KEYINPUT81), .B1(new_n234_), .B2(KEYINPUT1), .ZN(new_n244_));
  NOR3_X1   g043(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n236_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(new_n238_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n241_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n234_), .A2(KEYINPUT1), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT81), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n234_), .A2(KEYINPUT1), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n234_), .A2(KEYINPUT81), .A3(KEYINPUT1), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n251_), .A2(new_n252_), .A3(new_n253_), .A4(new_n233_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n247_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n254_), .A2(KEYINPUT82), .A3(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n240_), .B1(new_n248_), .B2(new_n256_), .ZN(new_n257_));
  OAI221_X1 g056(.A(new_n229_), .B1(new_n230_), .B2(new_n231_), .C1(new_n232_), .C2(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT87), .B1(new_n257_), .B2(new_n232_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n240_), .ZN(new_n260_));
  AND3_X1   g059(.A1(new_n254_), .A2(KEYINPUT82), .A3(new_n255_), .ZN(new_n261_));
  AOI21_X1  g060(.A(KEYINPUT82), .B1(new_n254_), .B2(new_n255_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n260_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT87), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(new_n264_), .A3(KEYINPUT29), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n259_), .A2(new_n229_), .A3(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n230_), .A2(new_n231_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n266_), .A2(KEYINPUT88), .A3(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(KEYINPUT88), .B1(new_n266_), .B2(new_n267_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n258_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(G78gat), .B(G106gat), .Z(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n257_), .A2(new_n232_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT28), .ZN(new_n274_));
  XOR2_X1   g073(.A(G22gat), .B(G50gat), .Z(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n271_), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n277_), .B(new_n258_), .C1(new_n268_), .C2(new_n269_), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n272_), .A2(new_n276_), .A3(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n276_), .B1(new_n272_), .B2(new_n278_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT27), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G183gat), .A2(G190gat), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT23), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(G183gat), .ZN(new_n289_));
  INV_X1    g088(.A(G190gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n288_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT22), .B(G169gat), .ZN(new_n295_));
  INV_X1    g094(.A(G176gat), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n294_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n292_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT26), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n300_), .A2(G190gat), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n290_), .A2(KEYINPUT26), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT89), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT25), .B(G183gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n290_), .A2(KEYINPUT26), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n300_), .A2(G190gat), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT89), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n303_), .A2(new_n304_), .A3(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT90), .B(KEYINPUT24), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT76), .ZN(new_n311_));
  INV_X1    g110(.A(G169gat), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n311_), .A2(new_n312_), .A3(new_n296_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT76), .B1(G169gat), .B2(G176gat), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n310_), .A2(new_n313_), .A3(new_n314_), .A4(new_n293_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n309_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n314_), .ZN(new_n317_));
  AND2_X1   g116(.A1(KEYINPUT90), .A2(KEYINPUT24), .ZN(new_n318_));
  NOR2_X1   g117(.A1(KEYINPUT90), .A2(KEYINPUT24), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n317_), .A2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(KEYINPUT91), .B1(new_n321_), .B2(new_n288_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n316_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(KEYINPUT91), .A3(new_n288_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n299_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  AOI22_X1  g124(.A1(new_n218_), .A2(new_n223_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT92), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT91), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n310_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n328_), .B1(new_n329_), .B2(new_n287_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n330_), .A2(new_n324_), .A3(new_n309_), .A4(new_n315_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(new_n298_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT92), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n229_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT20), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n295_), .A2(new_n296_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n293_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT77), .ZN(new_n338_));
  AOI22_X1  g137(.A1(new_n337_), .A2(new_n338_), .B1(new_n288_), .B2(new_n291_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n297_), .A2(KEYINPUT77), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n304_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n313_), .A2(KEYINPUT24), .A3(new_n314_), .A4(new_n293_), .ZN(new_n342_));
  AND3_X1   g141(.A1(new_n341_), .A2(new_n342_), .A3(new_n288_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT24), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n317_), .A2(new_n344_), .ZN(new_n345_));
  AOI22_X1  g144(.A1(new_n339_), .A2(new_n340_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n335_), .B1(new_n326_), .B2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n327_), .A2(new_n334_), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G226gat), .A2(G233gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT19), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n335_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT93), .ZN(new_n353_));
  INV_X1    g152(.A(new_n350_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n339_), .A2(new_n340_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n343_), .A2(new_n345_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n229_), .A2(new_n357_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n352_), .A2(new_n353_), .A3(new_n354_), .A4(new_n358_), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n224_), .A2(new_n331_), .A3(new_n228_), .A4(new_n298_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n358_), .A2(KEYINPUT20), .A3(new_n354_), .A4(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT93), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n351_), .A2(new_n359_), .A3(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G8gat), .B(G36gat), .Z(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT18), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G64gat), .B(G92gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n363_), .A2(new_n368_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n351_), .A2(new_n367_), .A3(new_n362_), .A4(new_n359_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n333_), .B1(new_n229_), .B2(new_n332_), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT20), .B1(new_n229_), .B2(new_n357_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n374_), .A2(KEYINPUT98), .A3(new_n354_), .A4(new_n334_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT98), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n376_), .B1(new_n348_), .B2(new_n350_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT97), .ZN(new_n379_));
  AOI211_X1 g178(.A(new_n379_), .B(new_n354_), .C1(new_n352_), .C2(new_n358_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n358_), .A2(KEYINPUT20), .A3(new_n360_), .ZN(new_n381_));
  AOI21_X1  g180(.A(KEYINPUT97), .B1(new_n381_), .B2(new_n350_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n368_), .B1(new_n378_), .B2(new_n383_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n370_), .A2(KEYINPUT27), .ZN(new_n385_));
  AOI22_X1  g184(.A1(new_n282_), .A2(new_n371_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n281_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G227gat), .A2(G233gat), .ZN(new_n388_));
  INV_X1    g187(.A(G15gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n357_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT31), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G113gat), .B(G120gat), .ZN(new_n393_));
  INV_X1    g192(.A(G134gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(G127gat), .ZN(new_n395_));
  INV_X1    g194(.A(G127gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(G134gat), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n395_), .A2(new_n397_), .A3(KEYINPUT79), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(KEYINPUT79), .B1(new_n395_), .B2(new_n397_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n393_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n395_), .A2(new_n397_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT79), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n393_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n404_), .A2(new_n398_), .A3(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n401_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT80), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n401_), .A2(KEYINPUT80), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G71gat), .B(G99gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(G43gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT78), .B(KEYINPUT30), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n411_), .B(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n392_), .B(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n407_), .B(new_n260_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n419_));
  OAI211_X1 g218(.A(KEYINPUT4), .B(new_n419_), .C1(new_n411_), .C2(new_n257_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT4), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n263_), .A2(new_n421_), .A3(new_n410_), .A4(new_n409_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G225gat), .A2(G233gat), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n420_), .A2(new_n422_), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT94), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n419_), .B1(new_n411_), .B2(new_n257_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  AOI22_X1  g227(.A1(new_n425_), .A2(new_n426_), .B1(new_n428_), .B2(new_n423_), .ZN(new_n429_));
  XOR2_X1   g228(.A(G1gat), .B(G29gat), .Z(new_n430_));
  XNOR2_X1  g229(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G57gat), .B(G85gat), .ZN(new_n433_));
  XOR2_X1   g232(.A(new_n432_), .B(new_n433_), .Z(new_n434_));
  NAND4_X1  g233(.A1(new_n420_), .A2(new_n422_), .A3(KEYINPUT94), .A4(new_n424_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n429_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n434_), .B1(new_n429_), .B2(new_n435_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n418_), .A2(new_n439_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n387_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT99), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n384_), .A2(new_n385_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n370_), .ZN(new_n444_));
  AOI22_X1  g243(.A1(new_n348_), .A2(new_n350_), .B1(new_n361_), .B2(KEYINPUT93), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n367_), .B1(new_n445_), .B2(new_n359_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n282_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n443_), .A2(new_n447_), .A3(new_n439_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n442_), .B1(new_n281_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n276_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n269_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n266_), .A2(KEYINPUT88), .A3(new_n267_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n277_), .B1(new_n453_), .B2(new_n258_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n278_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n450_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n272_), .A2(new_n276_), .A3(new_n278_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n458_), .A2(new_n386_), .A3(KEYINPUT99), .A4(new_n439_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n367_), .A2(KEYINPUT32), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n460_), .B(KEYINPUT96), .Z(new_n461_));
  OAI22_X1  g260(.A1(new_n437_), .A2(new_n438_), .B1(new_n363_), .B2(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n378_), .A2(new_n383_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n463_), .A2(new_n460_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT33), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n436_), .A2(new_n465_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n429_), .A2(KEYINPUT33), .A3(new_n434_), .A4(new_n435_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n420_), .A2(new_n423_), .A3(new_n422_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n434_), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n469_), .B(new_n470_), .C1(new_n427_), .C2(new_n423_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n369_), .A2(new_n370_), .A3(new_n471_), .ZN(new_n472_));
  OAI22_X1  g271(.A1(new_n462_), .A2(new_n464_), .B1(new_n468_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(new_n281_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n449_), .A2(new_n459_), .A3(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n441_), .B1(new_n475_), .B2(new_n417_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  OR2_X1    g276(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n478_));
  INV_X1    g277(.A(G106gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  AND3_X1   g280(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n482_));
  AOI21_X1  g281(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(G85gat), .ZN(new_n485_));
  INV_X1    g284(.A(G92gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G85gat), .A2(G92gat), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(KEYINPUT9), .A3(new_n488_), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n488_), .A2(KEYINPUT9), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n481_), .A2(new_n484_), .A3(new_n489_), .A4(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT7), .ZN(new_n492_));
  INV_X1    g291(.A(G99gat), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n492_), .A2(new_n493_), .A3(new_n479_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G99gat), .A2(G106gat), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT6), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n494_), .A2(new_n497_), .A3(new_n498_), .A4(new_n499_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n487_), .A2(new_n488_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT8), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n502_), .A2(KEYINPUT64), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n500_), .A2(new_n501_), .A3(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n504_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n491_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT65), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT65), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n509_), .B(new_n491_), .C1(new_n505_), .C2(new_n506_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G57gat), .B(G64gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G71gat), .B(G78gat), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n512_), .A3(KEYINPUT11), .ZN(new_n513_));
  XOR2_X1   g312(.A(G71gat), .B(G78gat), .Z(new_n514_));
  INV_X1    g313(.A(G64gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(G57gat), .ZN(new_n516_));
  INV_X1    g315(.A(G57gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(G64gat), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n516_), .A2(new_n518_), .A3(KEYINPUT11), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n514_), .A2(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n511_), .A2(KEYINPUT11), .ZN(new_n521_));
  OAI211_X1 g320(.A(KEYINPUT12), .B(new_n513_), .C1(new_n520_), .C2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n508_), .A2(new_n510_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G230gat), .A2(G233gat), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n513_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n526_), .B(new_n491_), .C1(new_n505_), .C2(new_n506_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT12), .ZN(new_n528_));
  AND4_X1   g327(.A1(new_n481_), .A2(new_n484_), .A3(new_n489_), .A4(new_n490_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n500_), .A2(new_n501_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(new_n503_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n500_), .A2(new_n501_), .A3(new_n504_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n529_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n528_), .B1(new_n533_), .B2(new_n526_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n524_), .A2(new_n525_), .A3(new_n527_), .A4(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT66), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n525_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n533_), .A2(new_n526_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n527_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n538_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n526_), .ZN(new_n542_));
  AOI21_X1  g341(.A(KEYINPUT12), .B1(new_n507_), .B2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n543_), .A2(new_n540_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n544_), .A2(KEYINPUT66), .A3(new_n525_), .A4(new_n524_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n537_), .A2(new_n541_), .A3(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(G120gat), .B(G148gat), .Z(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G176gat), .B(G204gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n546_), .B(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT13), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n552_), .A2(new_n553_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G29gat), .B(G36gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G43gat), .B(G50gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT73), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G15gat), .B(G22gat), .ZN(new_n562_));
  INV_X1    g361(.A(G1gat), .ZN(new_n563_));
  INV_X1    g362(.A(G8gat), .ZN(new_n564_));
  OAI21_X1  g363(.A(KEYINPUT14), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n562_), .A2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G1gat), .B(G8gat), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n566_), .B(new_n567_), .Z(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n561_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT73), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n560_), .B(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(new_n568_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n570_), .A2(new_n573_), .A3(KEYINPUT74), .ZN(new_n574_));
  OR3_X1    g373(.A1(new_n572_), .A2(KEYINPUT74), .A3(new_n568_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G229gat), .A2(G233gat), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n574_), .A2(new_n575_), .A3(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n560_), .B(KEYINPUT15), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(new_n569_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n573_), .A2(new_n580_), .A3(new_n576_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n578_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G113gat), .B(G141gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G169gat), .B(G197gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT75), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n582_), .B(new_n587_), .Z(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n557_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n568_), .B(new_n526_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G231gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT72), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G127gat), .B(G155gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT16), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G183gat), .B(G211gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT17), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n595_), .B(new_n600_), .ZN(new_n601_));
  OR3_X1    g400(.A1(new_n593_), .A2(KEYINPUT17), .A3(new_n599_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n590_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G232gat), .A2(G233gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT34), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT35), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT71), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n533_), .A2(new_n560_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT68), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT68), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n533_), .A2(new_n613_), .A3(new_n560_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n607_), .A2(new_n608_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n612_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n508_), .A2(new_n510_), .ZN(new_n617_));
  AOI211_X1 g416(.A(new_n610_), .B(new_n616_), .C1(new_n579_), .C2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT69), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n616_), .A2(new_n619_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n612_), .A2(KEYINPUT69), .A3(new_n614_), .A4(new_n615_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n617_), .A2(new_n579_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n620_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n618_), .B1(new_n609_), .B2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(KEYINPUT36), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT36), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n623_), .A2(new_n609_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n626_), .B1(new_n627_), .B2(new_n618_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G190gat), .B(G218gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT70), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(G134gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(G162gat), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n625_), .A2(new_n628_), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT37), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n626_), .B(new_n632_), .C1(new_n627_), .C2(new_n618_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n634_), .A2(new_n635_), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n635_), .B1(new_n634_), .B2(new_n636_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n604_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n477_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT100), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n439_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n477_), .A2(KEYINPUT100), .A3(new_n641_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n644_), .A2(new_n563_), .A3(new_n645_), .A4(new_n646_), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n647_), .A2(KEYINPUT101), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(KEYINPUT101), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT38), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n648_), .A2(KEYINPUT38), .A3(new_n649_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n604_), .B(KEYINPUT102), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n634_), .A2(new_n636_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n476_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n654_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT103), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n654_), .A2(new_n657_), .A3(KEYINPUT103), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n439_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n652_), .B(new_n653_), .C1(new_n563_), .C2(new_n662_), .ZN(G1324gat));
  OAI21_X1  g462(.A(G8gat), .B1(new_n658_), .B2(new_n386_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT39), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n386_), .A2(G8gat), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n644_), .A2(new_n646_), .A3(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT104), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n665_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT40), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n665_), .A2(new_n668_), .A3(KEYINPUT40), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1325gat));
  INV_X1    g472(.A(new_n642_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n674_), .A2(new_n389_), .A3(new_n418_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n660_), .A2(new_n661_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n389_), .B1(new_n676_), .B2(new_n418_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n677_), .A2(KEYINPUT41), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(KEYINPUT41), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n675_), .B1(new_n678_), .B2(new_n679_), .ZN(G1326gat));
  INV_X1    g479(.A(G22gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n674_), .A2(new_n681_), .A3(new_n458_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n281_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n683_), .A2(new_n681_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n684_), .A2(KEYINPUT42), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n684_), .A2(KEYINPUT42), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n682_), .B1(new_n685_), .B2(new_n686_), .ZN(G1327gat));
  INV_X1    g486(.A(new_n603_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n656_), .A2(new_n688_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n689_), .A2(new_n589_), .A3(new_n557_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n458_), .A2(new_n386_), .A3(new_n439_), .ZN(new_n691_));
  AOI22_X1  g490(.A1(new_n691_), .A2(new_n442_), .B1(new_n281_), .B2(new_n473_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n418_), .B1(new_n692_), .B2(new_n459_), .ZN(new_n693_));
  OAI211_X1 g492(.A(KEYINPUT105), .B(new_n690_), .C1(new_n693_), .C2(new_n441_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n590_), .A2(new_n688_), .A3(new_n656_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(new_n476_), .B2(new_n696_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n694_), .A2(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G29gat), .B1(new_n698_), .B2(new_n645_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n640_), .B1(new_n693_), .B2(new_n441_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n603_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  OAI211_X1 g501(.A(KEYINPUT43), .B(new_n640_), .C1(new_n693_), .C2(new_n441_), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n702_), .A2(KEYINPUT44), .A3(new_n590_), .A4(new_n703_), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n704_), .A2(G29gat), .A3(new_n645_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n640_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n701_), .B1(new_n476_), .B2(new_n706_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n703_), .A2(new_n707_), .A3(new_n590_), .A4(new_n688_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n699_), .B1(new_n705_), .B2(new_n710_), .ZN(G1328gat));
  INV_X1    g510(.A(G36gat), .ZN(new_n712_));
  INV_X1    g511(.A(new_n386_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n698_), .A2(new_n712_), .A3(new_n713_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT45), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n704_), .A2(new_n710_), .A3(new_n713_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(G36gat), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT46), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n715_), .A2(new_n717_), .A3(KEYINPUT46), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1329gat));
  XNOR2_X1  g521(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n694_), .A2(new_n697_), .A3(new_n418_), .ZN(new_n725_));
  INV_X1    g524(.A(G43gat), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT106), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n725_), .A2(new_n729_), .A3(new_n726_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n417_), .A2(new_n726_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n704_), .A2(new_n710_), .A3(new_n733_), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n731_), .A2(new_n732_), .A3(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n732_), .B1(new_n731_), .B2(new_n734_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n724_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n729_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n730_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n710_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n733_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n741_));
  OAI22_X1  g540(.A1(new_n738_), .A2(new_n739_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT108), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n731_), .A2(new_n732_), .A3(new_n734_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(new_n744_), .A3(new_n723_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n737_), .A2(new_n745_), .ZN(G1330gat));
  NAND3_X1  g545(.A1(new_n704_), .A2(new_n710_), .A3(new_n458_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(G50gat), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n281_), .A2(G50gat), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT109), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n698_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n748_), .A2(new_n751_), .ZN(G1331gat));
  NOR2_X1   g551(.A1(new_n556_), .A2(new_n588_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n477_), .A2(new_n753_), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n754_), .A2(new_n688_), .A3(new_n640_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n755_), .A2(new_n517_), .A3(new_n645_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n753_), .A2(new_n603_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n476_), .A2(new_n656_), .A3(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(G57gat), .B1(new_n759_), .B2(new_n439_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n756_), .A2(new_n760_), .ZN(G1332gat));
  NAND3_X1  g560(.A1(new_n755_), .A2(new_n515_), .A3(new_n713_), .ZN(new_n762_));
  OAI21_X1  g561(.A(G64gat), .B1(new_n759_), .B2(new_n386_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n763_), .A2(KEYINPUT48), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n763_), .A2(KEYINPUT48), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n762_), .B1(new_n764_), .B2(new_n765_), .ZN(G1333gat));
  INV_X1    g565(.A(G71gat), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n755_), .A2(new_n767_), .A3(new_n418_), .ZN(new_n768_));
  OAI21_X1  g567(.A(G71gat), .B1(new_n759_), .B2(new_n417_), .ZN(new_n769_));
  XOR2_X1   g568(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n770_));
  AND2_X1   g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n769_), .A2(new_n770_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n771_), .B2(new_n772_), .ZN(G1334gat));
  INV_X1    g572(.A(G78gat), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n755_), .A2(new_n774_), .A3(new_n458_), .ZN(new_n775_));
  OAI21_X1  g574(.A(G78gat), .B1(new_n759_), .B2(new_n281_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n776_), .A2(KEYINPUT50), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(KEYINPUT50), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n775_), .B1(new_n777_), .B2(new_n778_), .ZN(G1335gat));
  NAND4_X1  g578(.A1(new_n703_), .A2(new_n707_), .A3(new_n688_), .A4(new_n753_), .ZN(new_n780_));
  OAI21_X1  g579(.A(G85gat), .B1(new_n780_), .B2(new_n439_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n754_), .A2(new_n689_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n782_), .A2(new_n485_), .A3(new_n645_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(G1336gat));
  OAI21_X1  g583(.A(G92gat), .B1(new_n780_), .B2(new_n386_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n782_), .A2(new_n486_), .A3(new_n713_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(G1337gat));
  OAI21_X1  g586(.A(G99gat), .B1(new_n780_), .B2(new_n417_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n782_), .A2(new_n418_), .A3(new_n478_), .A4(new_n480_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g590(.A(G106gat), .B1(new_n780_), .B2(new_n281_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(new_n795_));
  OAI211_X1 g594(.A(G106gat), .B(new_n793_), .C1(new_n780_), .C2(new_n281_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n782_), .A2(new_n479_), .A3(new_n458_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n799_), .B(new_n800_), .ZN(G1339gat));
  NOR3_X1   g600(.A1(new_n554_), .A2(new_n555_), .A3(new_n588_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n603_), .B(new_n802_), .C1(new_n638_), .C2(new_n639_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n803_), .B(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT57), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n582_), .A2(new_n585_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n574_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n585_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT116), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n573_), .A2(new_n580_), .A3(new_n577_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n809_), .A2(KEYINPUT116), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n807_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n814_), .A2(new_n552_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n537_), .A2(new_n817_), .A3(new_n545_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n544_), .A2(new_n524_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n538_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n544_), .A2(KEYINPUT55), .A3(new_n525_), .A4(new_n524_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n822_), .B(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n816_), .B1(new_n821_), .B2(new_n824_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n822_), .B(KEYINPUT113), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n826_), .A2(KEYINPUT114), .A3(new_n818_), .A4(new_n820_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n551_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT56), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n828_), .A2(KEYINPUT56), .A3(new_n551_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n831_), .A2(new_n832_), .A3(new_n833_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n828_), .A2(KEYINPUT115), .A3(KEYINPUT56), .A4(new_n551_), .ZN(new_n835_));
  OR2_X1    g634(.A1(new_n546_), .A2(new_n551_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n588_), .A2(new_n836_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n835_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n815_), .B1(new_n834_), .B2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n806_), .B1(new_n839_), .B2(new_n656_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n835_), .A2(new_n837_), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT56), .B1(new_n828_), .B2(new_n551_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n551_), .ZN(new_n843_));
  AOI211_X1 g642(.A(new_n830_), .B(new_n843_), .C1(new_n825_), .C2(new_n827_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n842_), .A2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n841_), .B1(new_n845_), .B2(new_n832_), .ZN(new_n846_));
  OAI211_X1 g645(.A(KEYINPUT57), .B(new_n655_), .C1(new_n846_), .C2(new_n815_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n831_), .A2(new_n833_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n848_), .A2(KEYINPUT58), .A3(new_n836_), .A4(new_n814_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT58), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n814_), .A2(new_n836_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n845_), .B2(new_n851_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n849_), .A2(new_n852_), .A3(new_n640_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n840_), .A2(new_n847_), .A3(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n805_), .B1(new_n854_), .B2(new_n688_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n387_), .A2(new_n439_), .A3(new_n417_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n855_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(G113gat), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n858_), .A2(new_n859_), .A3(new_n588_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n854_), .A2(new_n688_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n805_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n863_), .A2(KEYINPUT59), .A3(new_n856_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(new_n855_), .B2(new_n857_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n589_), .B1(new_n864_), .B2(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n860_), .B1(new_n867_), .B2(new_n859_), .ZN(G1340gat));
  AOI21_X1  g667(.A(new_n556_), .B1(new_n864_), .B2(new_n866_), .ZN(new_n869_));
  INV_X1    g668(.A(G120gat), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n858_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n870_), .B1(new_n556_), .B2(KEYINPUT60), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(KEYINPUT60), .B2(new_n870_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n872_), .A2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(KEYINPUT117), .B1(new_n871_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT117), .ZN(new_n877_));
  OAI221_X1 g676(.A(new_n877_), .B1(new_n872_), .B2(new_n874_), .C1(new_n869_), .C2(new_n870_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(G1341gat));
  NAND3_X1  g678(.A1(new_n858_), .A2(new_n396_), .A3(new_n603_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n688_), .B1(new_n864_), .B2(new_n866_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n881_), .B2(new_n396_), .ZN(G1342gat));
  NAND3_X1  g681(.A1(new_n858_), .A2(new_n394_), .A3(new_n656_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n706_), .B1(new_n864_), .B2(new_n866_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n884_), .B2(new_n394_), .ZN(G1343gat));
  NOR4_X1   g684(.A1(new_n713_), .A2(new_n281_), .A3(new_n439_), .A4(new_n418_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n863_), .A2(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n589_), .ZN(new_n888_));
  XOR2_X1   g687(.A(new_n888_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g688(.A1(new_n887_), .A2(new_n556_), .ZN(new_n890_));
  XOR2_X1   g689(.A(new_n890_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g690(.A1(new_n887_), .A2(new_n688_), .ZN(new_n892_));
  XOR2_X1   g691(.A(KEYINPUT61), .B(G155gat), .Z(new_n893_));
  XNOR2_X1  g692(.A(new_n892_), .B(new_n893_), .ZN(G1346gat));
  OAI21_X1  g693(.A(G162gat), .B1(new_n887_), .B2(new_n706_), .ZN(new_n895_));
  OR2_X1    g694(.A1(new_n655_), .A2(G162gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n887_), .B2(new_n896_), .ZN(G1347gat));
  INV_X1    g696(.A(KEYINPUT118), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n855_), .A2(new_n458_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n440_), .A2(new_n386_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n899_), .A2(new_n588_), .A3(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n898_), .B1(new_n901_), .B2(G169gat), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n901_), .A2(new_n898_), .A3(G169gat), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n903_), .A2(KEYINPUT62), .A3(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n899_), .A2(new_n900_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n588_), .A2(new_n295_), .ZN(new_n908_));
  XOR2_X1   g707(.A(new_n908_), .B(KEYINPUT119), .Z(new_n909_));
  AOI22_X1  g708(.A1(new_n902_), .A2(new_n906_), .B1(new_n907_), .B2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n905_), .A2(new_n910_), .ZN(G1348gat));
  NAND2_X1  g710(.A1(new_n899_), .A2(new_n900_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n912_), .A2(new_n556_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(new_n296_), .ZN(G1349gat));
  INV_X1    g713(.A(new_n304_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n907_), .A2(new_n915_), .A3(new_n603_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(KEYINPUT120), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n289_), .B1(new_n912_), .B2(new_n688_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT120), .ZN(new_n919_));
  NAND4_X1  g718(.A1(new_n907_), .A2(new_n919_), .A3(new_n915_), .A4(new_n603_), .ZN(new_n920_));
  AND3_X1   g719(.A1(new_n917_), .A2(new_n918_), .A3(new_n920_), .ZN(G1350gat));
  OAI21_X1  g720(.A(G190gat), .B1(new_n912_), .B2(new_n706_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n656_), .A2(new_n303_), .A3(new_n308_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n922_), .B1(new_n912_), .B2(new_n923_), .ZN(G1351gat));
  NAND3_X1  g723(.A1(new_n458_), .A2(new_n439_), .A3(new_n417_), .ZN(new_n925_));
  OR2_X1    g724(.A1(new_n925_), .A2(KEYINPUT121), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n925_), .A2(KEYINPUT121), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n926_), .A2(new_n713_), .A3(new_n927_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n928_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(new_n588_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(KEYINPUT122), .B(G197gat), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n930_), .B(new_n931_), .ZN(G1352gat));
  NAND2_X1  g731(.A1(new_n929_), .A2(new_n557_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n203_), .A2(KEYINPUT123), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n933_), .B(new_n934_), .ZN(G1353gat));
  NAND2_X1  g734(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n603_), .A2(new_n936_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(KEYINPUT124), .ZN(new_n938_));
  NOR3_X1   g737(.A1(new_n855_), .A2(new_n928_), .A3(new_n938_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n939_), .B(new_n940_), .ZN(G1354gat));
  XOR2_X1   g740(.A(KEYINPUT126), .B(G218gat), .Z(new_n942_));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n943_), .B1(new_n929_), .B2(new_n656_), .ZN(new_n944_));
  NOR4_X1   g743(.A1(new_n855_), .A2(KEYINPUT125), .A3(new_n655_), .A4(new_n928_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n942_), .B1(new_n944_), .B2(new_n945_), .ZN(new_n946_));
  INV_X1    g745(.A(KEYINPUT127), .ZN(new_n947_));
  NOR3_X1   g746(.A1(new_n855_), .A2(new_n706_), .A3(new_n928_), .ZN(new_n948_));
  OR2_X1    g747(.A1(new_n948_), .A2(new_n942_), .ZN(new_n949_));
  AND3_X1   g748(.A1(new_n946_), .A2(new_n947_), .A3(new_n949_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n947_), .B1(new_n946_), .B2(new_n949_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n950_), .A2(new_n951_), .ZN(G1355gat));
endmodule


