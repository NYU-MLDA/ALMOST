//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 1 0 1 0 0 0 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n861_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  XOR2_X1   g001(.A(G211gat), .B(G218gat), .Z(new_n203_));
  INV_X1    g002(.A(KEYINPUT21), .ZN(new_n204_));
  INV_X1    g003(.A(G197gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G204gat), .ZN(new_n206_));
  INV_X1    g005(.A(G204gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G197gat), .ZN(new_n208_));
  AND2_X1   g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n203_), .B1(new_n204_), .B2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT86), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n208_), .B1(new_n206_), .B2(new_n211_), .ZN(new_n212_));
  AOI21_X1  g011(.A(KEYINPUT86), .B1(new_n205_), .B2(G204gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT21), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n210_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n209_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(KEYINPUT21), .A3(new_n203_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n218_), .B(KEYINPUT87), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(G183gat), .A3(G190gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT82), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G183gat), .ZN(new_n225_));
  INV_X1    g024(.A(G190gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT23), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT81), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n227_), .A2(KEYINPUT81), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n224_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT77), .B(G183gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n230_), .B1(G190gat), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT22), .B(G169gat), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n236_), .A2(KEYINPUT80), .ZN(new_n237_));
  INV_X1    g036(.A(G176gat), .ZN(new_n238_));
  INV_X1    g037(.A(G169gat), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n239_), .A2(KEYINPUT22), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n238_), .B1(new_n240_), .B2(KEYINPUT80), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n233_), .B(new_n234_), .C1(new_n237_), .C2(new_n241_), .ZN(new_n242_));
  OR2_X1    g041(.A1(new_n227_), .A2(KEYINPUT79), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n227_), .A2(KEYINPUT79), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(new_n222_), .A3(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n234_), .A2(KEYINPUT24), .ZN(new_n246_));
  NOR2_X1   g045(.A1(G169gat), .A2(G176gat), .ZN(new_n247_));
  MUX2_X1   g046(.A(new_n246_), .B(KEYINPUT24), .S(new_n247_), .Z(new_n248_));
  INV_X1    g047(.A(KEYINPUT25), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(new_n225_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n250_), .B1(new_n231_), .B2(new_n249_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT78), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n252_), .A2(new_n249_), .ZN(new_n253_));
  AOI22_X1  g052(.A1(new_n251_), .A2(new_n252_), .B1(new_n231_), .B2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT26), .B(G190gat), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n245_), .B(new_n248_), .C1(new_n254_), .C2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n242_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT83), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n242_), .A2(KEYINPUT83), .A3(new_n257_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n220_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G226gat), .A2(G233gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT19), .ZN(new_n264_));
  XOR2_X1   g063(.A(KEYINPUT25), .B(G183gat), .Z(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT91), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n234_), .A2(KEYINPUT92), .A3(KEYINPUT24), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT92), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n247_), .B1(new_n246_), .B2(new_n268_), .ZN(new_n269_));
  AOI22_X1  g068(.A1(new_n266_), .A2(new_n255_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n247_), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n270_), .B(new_n230_), .C1(KEYINPUT24), .C2(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n245_), .B1(G183gat), .B2(G190gat), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n273_), .B(new_n234_), .C1(G176gat), .C2(new_n236_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT20), .B1(new_n275_), .B2(new_n218_), .ZN(new_n276_));
  OR3_X1    g075(.A1(new_n262_), .A2(new_n264_), .A3(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n260_), .A2(new_n261_), .A3(new_n220_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT20), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n279_), .B1(new_n275_), .B2(new_n218_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(new_n264_), .ZN(new_n282_));
  XOR2_X1   g081(.A(G64gat), .B(G92gat), .Z(new_n283_));
  XNOR2_X1  g082(.A(G8gat), .B(G36gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n286_));
  XOR2_X1   g085(.A(new_n285_), .B(new_n286_), .Z(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n277_), .A2(new_n282_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT97), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n202_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT96), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n292_), .B1(new_n281_), .B2(new_n264_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n264_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n278_), .A2(KEYINPUT96), .A3(new_n294_), .A4(new_n280_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n264_), .B1(new_n262_), .B2(new_n276_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n293_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n287_), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n291_), .B(new_n298_), .C1(new_n290_), .C2(new_n289_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n277_), .A2(new_n282_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(new_n287_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n289_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(new_n202_), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n299_), .A2(new_n303_), .ZN(new_n304_));
  XOR2_X1   g103(.A(G155gat), .B(G162gat), .Z(new_n305_));
  NOR2_X1   g104(.A1(G141gat), .A2(G148gat), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n306_), .B(KEYINPUT3), .Z(new_n307_));
  NAND2_X1  g106(.A1(G141gat), .A2(G148gat), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n308_), .B(KEYINPUT2), .Z(new_n309_));
  OAI21_X1  g108(.A(new_n305_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT1), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n305_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n306_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n312_), .A2(new_n313_), .A3(new_n308_), .A4(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n310_), .A2(new_n315_), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n316_), .A2(KEYINPUT29), .ZN(new_n317_));
  XOR2_X1   g116(.A(G22gat), .B(G50gat), .Z(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT28), .ZN(new_n319_));
  XOR2_X1   g118(.A(new_n317_), .B(new_n319_), .Z(new_n320_));
  NAND2_X1  g119(.A1(new_n316_), .A2(KEYINPUT29), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(new_n218_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n322_), .A2(G228gat), .A3(G233gat), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  AOI22_X1  g123(.A1(new_n316_), .A2(KEYINPUT29), .B1(G228gat), .B2(G233gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n219_), .A2(new_n325_), .ZN(new_n326_));
  OR2_X1    g125(.A1(new_n326_), .A2(KEYINPUT88), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(KEYINPUT88), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n324_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G78gat), .B(G106gat), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n320_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n329_), .A2(new_n331_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n333_), .A2(KEYINPUT90), .A3(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT89), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n327_), .A2(new_n328_), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n336_), .B(new_n330_), .C1(new_n337_), .C2(new_n324_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n320_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n334_), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT89), .B1(new_n329_), .B2(new_n331_), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n338_), .B(new_n339_), .C1(new_n340_), .C2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT90), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n343_), .B1(new_n340_), .B2(new_n332_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n335_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n304_), .A2(new_n346_), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n260_), .A2(new_n261_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT30), .ZN(new_n349_));
  OR2_X1    g148(.A1(new_n349_), .A2(KEYINPUT85), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(KEYINPUT85), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT84), .ZN(new_n353_));
  XOR2_X1   g152(.A(G127gat), .B(G134gat), .Z(new_n354_));
  XOR2_X1   g153(.A(G113gat), .B(G120gat), .Z(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT31), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n353_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n358_), .B1(new_n357_), .B2(new_n356_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G227gat), .A2(G233gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G71gat), .B(G99gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G15gat), .B(G43gat), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n363_), .B(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n352_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n363_), .B(new_n364_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n368_), .A2(new_n351_), .A3(new_n350_), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT94), .ZN(new_n371_));
  INV_X1    g170(.A(new_n356_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n316_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n356_), .A2(new_n310_), .A3(new_n315_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(KEYINPUT4), .A3(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT4), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n316_), .A2(new_n377_), .A3(new_n372_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G225gat), .A2(G233gat), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n371_), .B1(new_n376_), .B2(new_n381_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n375_), .A2(new_n378_), .A3(KEYINPUT94), .A4(new_n380_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n373_), .A2(new_n374_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(new_n379_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n382_), .A2(new_n383_), .A3(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G1gat), .B(G29gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT0), .ZN(new_n389_));
  INV_X1    g188(.A(G57gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(G85gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n387_), .A2(new_n393_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n382_), .A2(new_n392_), .A3(new_n383_), .A4(new_n386_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n370_), .A2(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n347_), .A2(new_n398_), .ZN(new_n399_));
  AND2_X1   g198(.A1(new_n345_), .A2(new_n397_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n304_), .A2(new_n400_), .A3(KEYINPUT98), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n395_), .A2(KEYINPUT33), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n395_), .A2(KEYINPUT33), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n375_), .A2(new_n379_), .A3(new_n378_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n392_), .B1(new_n385_), .B2(new_n380_), .ZN(new_n405_));
  AOI22_X1  g204(.A1(new_n402_), .A2(new_n403_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n301_), .A2(new_n406_), .A3(new_n289_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT95), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n297_), .A2(KEYINPUT32), .A3(new_n288_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n288_), .A2(KEYINPUT32), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n409_), .B(new_n396_), .C1(new_n300_), .C2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT95), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n301_), .A2(new_n406_), .A3(new_n413_), .A4(new_n289_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n408_), .A2(new_n412_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n346_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n299_), .A2(new_n345_), .A3(new_n397_), .A4(new_n303_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT98), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n401_), .A2(new_n416_), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n370_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n399_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT9), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G85gat), .A2(G92gat), .ZN(new_n424_));
  NOR2_X1   g223(.A1(G85gat), .A2(G92gat), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n423_), .B(new_n424_), .C1(new_n425_), .C2(KEYINPUT65), .ZN(new_n426_));
  AND2_X1   g225(.A1(G85gat), .A2(G92gat), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT65), .ZN(new_n428_));
  NOR3_X1   g227(.A1(new_n427_), .A2(new_n425_), .A3(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n426_), .B1(new_n429_), .B2(new_n423_), .ZN(new_n430_));
  AND2_X1   g229(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n431_));
  NOR2_X1   g230(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n432_));
  NOR3_X1   g231(.A1(new_n431_), .A2(new_n432_), .A3(G106gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G99gat), .A2(G106gat), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT6), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n433_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n430_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT7), .ZN(new_n441_));
  INV_X1    g240(.A(G99gat), .ZN(new_n442_));
  INV_X1    g241(.A(G106gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n441_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n444_), .A2(new_n436_), .A3(new_n437_), .A4(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n427_), .A2(new_n425_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT8), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n446_), .A2(KEYINPUT8), .A3(new_n447_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n440_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT12), .ZN(new_n453_));
  XOR2_X1   g252(.A(G71gat), .B(G78gat), .Z(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(G64gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(G57gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n390_), .A2(G64gat), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT67), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n457_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n459_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT11), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n390_), .A2(G64gat), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n456_), .A2(G57gat), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT67), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT11), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n457_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n455_), .B1(new_n462_), .B2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n466_), .B1(new_n465_), .B2(new_n467_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n470_), .A2(new_n454_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n453_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT66), .ZN(new_n474_));
  AOI22_X1  g273(.A1(new_n430_), .A2(new_n439_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n474_), .B1(new_n475_), .B2(new_n451_), .ZN(new_n476_));
  AND4_X1   g275(.A1(new_n474_), .A2(new_n440_), .A3(new_n451_), .A4(new_n450_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NOR3_X1   g277(.A1(new_n460_), .A2(new_n461_), .A3(KEYINPUT11), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n454_), .B1(new_n479_), .B2(new_n470_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n462_), .A2(new_n455_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT68), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n480_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT68), .B1(new_n469_), .B2(new_n471_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n473_), .B1(new_n478_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT12), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n487_), .B1(new_n478_), .B2(new_n485_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G230gat), .A2(G233gat), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n489_), .B(KEYINPUT64), .Z(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n486_), .A2(new_n488_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n452_), .A2(KEYINPUT66), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n475_), .A2(new_n474_), .A3(new_n451_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n485_), .B(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n492_), .B1(new_n491_), .B2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G120gat), .B(G148gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(new_n207_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT5), .B(G176gat), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n499_), .B(new_n500_), .Z(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n497_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT69), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n497_), .A2(new_n502_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n497_), .A2(KEYINPUT69), .A3(new_n502_), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n506_), .A2(KEYINPUT13), .A3(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT13), .B1(new_n506_), .B2(new_n507_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT74), .B(G1gat), .ZN(new_n511_));
  INV_X1    g310(.A(G8gat), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT14), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G15gat), .B(G22gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(G1gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(G8gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n515_), .B(G1gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(new_n512_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G29gat), .B(G36gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G43gat), .B(G50gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n521_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G229gat), .A2(G233gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n524_), .B(KEYINPUT15), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n518_), .A2(new_n520_), .A3(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n525_), .A2(new_n526_), .A3(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n524_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n521_), .B(new_n530_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n529_), .B1(new_n531_), .B2(new_n526_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G113gat), .B(G141gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(G169gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(new_n205_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n532_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT76), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n529_), .B(new_n535_), .C1(new_n531_), .C2(new_n526_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n537_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n532_), .A2(KEYINPUT76), .A3(new_n536_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT37), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G232gat), .A2(G233gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT34), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT35), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT70), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n478_), .A2(new_n524_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n527_), .A2(new_n452_), .B1(new_n547_), .B2(new_n546_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n550_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n548_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n554_), .A2(KEYINPUT70), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n553_), .A2(new_n556_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n551_), .A2(new_n549_), .A3(new_n548_), .A4(new_n552_), .ZN(new_n558_));
  XOR2_X1   g357(.A(G134gat), .B(G162gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(G190gat), .B(G218gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT36), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n557_), .A2(new_n558_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT36), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n561_), .A2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT71), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  AOI211_X1 g367(.A(new_n555_), .B(new_n550_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n558_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n568_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT72), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n557_), .A2(new_n558_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n574_), .A2(KEYINPUT72), .A3(new_n568_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n564_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT73), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  AOI211_X1 g377(.A(KEYINPUT73), .B(new_n564_), .C1(new_n573_), .C2(new_n575_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n543_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(KEYINPUT72), .B1(new_n574_), .B2(new_n568_), .ZN(new_n581_));
  AOI211_X1 g380(.A(new_n572_), .B(new_n567_), .C1(new_n557_), .C2(new_n558_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n563_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT73), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n576_), .A2(new_n577_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(new_n585_), .A3(KEYINPUT37), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n580_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  AND2_X1   g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n521_), .B(new_n589_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n590_), .A2(new_n472_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n472_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G127gat), .B(G155gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT16), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(G183gat), .ZN(new_n595_));
  INV_X1    g394(.A(G211gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT17), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n591_), .A2(new_n592_), .A3(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n483_), .A2(new_n484_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n590_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n590_), .A2(new_n601_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n597_), .B(KEYINPUT17), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n602_), .A2(new_n603_), .A3(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n600_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT75), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT75), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n600_), .A2(new_n605_), .A3(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n588_), .A2(new_n610_), .ZN(new_n611_));
  NOR4_X1   g410(.A1(new_n422_), .A2(new_n510_), .A3(new_n542_), .A4(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n612_), .A2(new_n396_), .A3(new_n511_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT99), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT38), .ZN(new_n615_));
  INV_X1    g414(.A(new_n610_), .ZN(new_n616_));
  NOR3_X1   g415(.A1(new_n422_), .A2(new_n576_), .A3(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n510_), .A2(new_n542_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  OAI21_X1  g418(.A(G1gat), .B1(new_n619_), .B2(new_n397_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n615_), .A2(new_n620_), .ZN(G1324gat));
  INV_X1    g420(.A(new_n304_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n612_), .A2(new_n512_), .A3(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n617_), .A2(new_n618_), .A3(new_n622_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT39), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n624_), .A2(new_n625_), .A3(G8gat), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n625_), .B1(new_n624_), .B2(G8gat), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n623_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g429(.A(G15gat), .B1(new_n619_), .B2(new_n421_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT41), .Z(new_n632_));
  INV_X1    g431(.A(G15gat), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n612_), .A2(new_n633_), .A3(new_n370_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(G1326gat));
  OAI21_X1  g434(.A(G22gat), .B1(new_n619_), .B2(new_n346_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT42), .ZN(new_n637_));
  INV_X1    g436(.A(G22gat), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n612_), .A2(new_n638_), .A3(new_n345_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(G1327gat));
  NOR2_X1   g439(.A1(new_n610_), .A2(new_n583_), .ZN(new_n641_));
  AOI22_X1  g440(.A1(new_n417_), .A2(new_n418_), .B1(new_n415_), .B2(new_n346_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n370_), .B1(new_n642_), .B2(new_n401_), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n618_), .B(new_n641_), .C1(new_n643_), .C2(new_n399_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(G29gat), .B1(new_n645_), .B2(new_n396_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT43), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n647_), .B1(new_n422_), .B2(new_n588_), .ZN(new_n648_));
  OAI211_X1 g447(.A(KEYINPUT43), .B(new_n587_), .C1(new_n643_), .C2(new_n399_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n648_), .A2(new_n618_), .A3(new_n616_), .A4(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT44), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n650_), .A2(KEYINPUT100), .A3(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(KEYINPUT100), .B1(new_n650_), .B2(new_n651_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n650_), .A2(new_n651_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n656_), .A2(G29gat), .A3(new_n396_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n646_), .B1(new_n655_), .B2(new_n657_), .ZN(G1328gat));
  INV_X1    g457(.A(G36gat), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n622_), .A2(new_n659_), .ZN(new_n660_));
  OR3_X1    g459(.A1(new_n644_), .A2(KEYINPUT101), .A3(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(KEYINPUT101), .B1(new_n644_), .B2(new_n660_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n661_), .A2(KEYINPUT45), .A3(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(KEYINPUT45), .B1(new_n661_), .B2(new_n662_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n622_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n650_), .A2(new_n651_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT100), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n650_), .A2(KEYINPUT100), .A3(new_n651_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n666_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n665_), .B1(new_n671_), .B2(new_n659_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT46), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  OAI211_X1 g473(.A(KEYINPUT46), .B(new_n665_), .C1(new_n671_), .C2(new_n659_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1329gat));
  AOI21_X1  g475(.A(G43gat), .B1(new_n645_), .B2(new_n370_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n656_), .A2(G43gat), .A3(new_n370_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n678_), .B1(new_n654_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT47), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT47), .ZN(new_n682_));
  OAI211_X1 g481(.A(new_n682_), .B(new_n678_), .C1(new_n654_), .C2(new_n679_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(G1330gat));
  OR3_X1    g483(.A1(new_n644_), .A2(G50gat), .A3(new_n346_), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n345_), .B(new_n656_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n686_), .A2(new_n687_), .A3(G50gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n686_), .B2(G50gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n685_), .B1(new_n688_), .B2(new_n689_), .ZN(G1331gat));
  INV_X1    g489(.A(new_n422_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n510_), .ZN(new_n692_));
  OAI21_X1  g491(.A(KEYINPUT103), .B1(new_n611_), .B2(new_n692_), .ZN(new_n693_));
  OR3_X1    g492(.A1(new_n611_), .A2(KEYINPUT103), .A3(new_n692_), .ZN(new_n694_));
  AND4_X1   g493(.A1(new_n542_), .A2(new_n691_), .A3(new_n693_), .A4(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n695_), .A2(new_n390_), .A3(new_n396_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n542_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n692_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n617_), .A2(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(G57gat), .B1(new_n699_), .B2(new_n397_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n696_), .A2(new_n700_), .ZN(G1332gat));
  OAI21_X1  g500(.A(G64gat), .B1(new_n699_), .B2(new_n304_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT48), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n622_), .A2(new_n456_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT104), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n695_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n703_), .A2(new_n706_), .ZN(G1333gat));
  OAI21_X1  g506(.A(G71gat), .B1(new_n699_), .B2(new_n421_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT49), .ZN(new_n709_));
  INV_X1    g508(.A(G71gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n695_), .A2(new_n710_), .A3(new_n370_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n711_), .ZN(G1334gat));
  OAI21_X1  g511(.A(G78gat), .B1(new_n699_), .B2(new_n346_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT50), .ZN(new_n714_));
  INV_X1    g513(.A(G78gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n695_), .A2(new_n715_), .A3(new_n345_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1335gat));
  NAND4_X1  g516(.A1(new_n648_), .A2(new_n616_), .A3(new_n649_), .A4(new_n698_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n719_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n720_), .A2(new_n396_), .A3(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(G85gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n691_), .A2(new_n641_), .A3(new_n698_), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n397_), .A2(G85gat), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n723_), .B1(new_n724_), .B2(new_n725_), .ZN(G1336gat));
  INV_X1    g525(.A(new_n724_), .ZN(new_n727_));
  AOI21_X1  g526(.A(G92gat), .B1(new_n727_), .B2(new_n622_), .ZN(new_n728_));
  XOR2_X1   g527(.A(new_n728_), .B(KEYINPUT106), .Z(new_n729_));
  NAND4_X1  g528(.A1(new_n720_), .A2(G92gat), .A3(new_n622_), .A4(new_n721_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1337gat));
  INV_X1    g530(.A(KEYINPUT107), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT51), .ZN(new_n733_));
  OR3_X1    g532(.A1(new_n421_), .A2(new_n432_), .A3(new_n431_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(new_n724_), .B2(new_n734_), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n718_), .A2(new_n421_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n736_), .B2(G99gat), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n732_), .A2(KEYINPUT51), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n737_), .B(new_n738_), .ZN(G1338gat));
  NAND3_X1  g538(.A1(new_n727_), .A2(new_n443_), .A3(new_n345_), .ZN(new_n740_));
  OAI21_X1  g539(.A(G106gat), .B1(new_n718_), .B2(new_n346_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n741_), .A2(KEYINPUT52), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT52), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n743_), .B(G106gat), .C1(new_n718_), .C2(new_n346_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n740_), .B1(new_n742_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT53), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT53), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n748_), .B(new_n740_), .C1(new_n742_), .C2(new_n745_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1339gat));
  INV_X1    g549(.A(KEYINPUT59), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n347_), .A2(new_n421_), .A3(new_n397_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n539_), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n525_), .A2(G229gat), .A3(G233gat), .A4(new_n528_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n531_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n535_), .B1(new_n755_), .B2(new_n526_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n753_), .B1(new_n754_), .B2(new_n756_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n757_), .A2(new_n503_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT55), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n492_), .A2(new_n759_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n486_), .A2(new_n488_), .A3(KEYINPUT55), .A4(new_n491_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n486_), .A2(new_n488_), .ZN(new_n762_));
  AOI21_X1  g561(.A(KEYINPUT109), .B1(new_n762_), .B2(new_n490_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT109), .ZN(new_n764_));
  AOI211_X1 g563(.A(new_n764_), .B(new_n491_), .C1(new_n486_), .C2(new_n488_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n760_), .B(new_n761_), .C1(new_n763_), .C2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT110), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  OAI22_X1  g567(.A1(new_n601_), .A2(new_n495_), .B1(new_n472_), .B2(new_n453_), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT12), .B1(new_n601_), .B2(new_n495_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n490_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n764_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n762_), .A2(KEYINPUT109), .A3(new_n490_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n774_), .A2(KEYINPUT110), .A3(new_n760_), .A4(new_n761_), .ZN(new_n775_));
  AND4_X1   g574(.A1(KEYINPUT56), .A2(new_n768_), .A3(new_n502_), .A4(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n501_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT56), .B1(new_n777_), .B2(new_n775_), .ZN(new_n778_));
  OAI211_X1 g577(.A(KEYINPUT58), .B(new_n758_), .C1(new_n776_), .C2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n587_), .A2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n768_), .A2(new_n775_), .A3(new_n502_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT56), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n777_), .A2(KEYINPUT56), .A3(new_n775_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT58), .B1(new_n785_), .B2(new_n758_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n780_), .A2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n506_), .A2(new_n757_), .A3(new_n507_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n540_), .A2(new_n503_), .A3(new_n541_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n791_), .B1(new_n776_), .B2(new_n778_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT111), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n789_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n790_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT111), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n576_), .B1(new_n794_), .B2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n787_), .B1(new_n797_), .B2(KEYINPUT57), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n788_), .B1(new_n795_), .B2(KEYINPUT111), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n792_), .A2(new_n793_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n583_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT57), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n610_), .B1(new_n798_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n607_), .A2(new_n542_), .A3(new_n609_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n692_), .A2(KEYINPUT108), .A3(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT108), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n610_), .A2(new_n542_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n808_), .B1(new_n809_), .B2(new_n510_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n807_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n805_), .B1(new_n811_), .B2(new_n588_), .ZN(new_n812_));
  AOI211_X1 g611(.A(KEYINPUT54), .B(new_n587_), .C1(new_n807_), .C2(new_n810_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n751_), .B(new_n752_), .C1(new_n804_), .C2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n752_), .ZN(new_n816_));
  OAI21_X1  g615(.A(KEYINPUT112), .B1(new_n797_), .B2(KEYINPUT57), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT112), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n801_), .A2(new_n818_), .A3(new_n802_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n817_), .A2(new_n798_), .A3(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n616_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n814_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n816_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n815_), .B1(new_n823_), .B2(new_n751_), .ZN(new_n824_));
  OAI21_X1  g623(.A(G113gat), .B1(new_n824_), .B2(new_n542_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n821_), .A2(new_n822_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n752_), .ZN(new_n827_));
  OR2_X1    g626(.A1(new_n542_), .A2(G113gat), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n825_), .B1(new_n827_), .B2(new_n828_), .ZN(G1340gat));
  OAI211_X1 g628(.A(new_n510_), .B(new_n815_), .C1(new_n823_), .C2(new_n751_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(G120gat), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT60), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(G120gat), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n692_), .A2(KEYINPUT60), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n823_), .B(new_n833_), .C1(G120gat), .C2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n831_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT113), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n831_), .A2(KEYINPUT113), .A3(new_n835_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(G1341gat));
  OAI21_X1  g639(.A(G127gat), .B1(new_n824_), .B2(new_n616_), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n616_), .A2(G127gat), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n827_), .B2(new_n842_), .ZN(G1342gat));
  INV_X1    g642(.A(G134gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n827_), .B2(new_n583_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n587_), .A2(G134gat), .ZN(new_n846_));
  XOR2_X1   g645(.A(new_n846_), .B(KEYINPUT114), .Z(new_n847_));
  OAI211_X1 g646(.A(new_n815_), .B(new_n847_), .C1(new_n823_), .C2(new_n751_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n845_), .A2(new_n848_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(KEYINPUT115), .ZN(G1343gat));
  INV_X1    g649(.A(KEYINPUT117), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n421_), .A2(new_n396_), .A3(new_n304_), .A4(new_n345_), .ZN(new_n852_));
  XOR2_X1   g651(.A(new_n852_), .B(KEYINPUT116), .Z(new_n853_));
  NAND3_X1  g652(.A1(new_n826_), .A2(new_n851_), .A3(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n814_), .B1(new_n820_), .B2(new_n616_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n853_), .ZN(new_n856_));
  OAI21_X1  g655(.A(KEYINPUT117), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n542_), .B1(new_n854_), .B2(new_n857_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(KEYINPUT118), .B(G141gat), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(G1344gat));
  NAND2_X1  g659(.A1(new_n854_), .A2(new_n857_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n510_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G148gat), .ZN(G1345gat));
  AOI21_X1  g662(.A(new_n616_), .B1(new_n854_), .B2(new_n857_), .ZN(new_n864_));
  XOR2_X1   g663(.A(KEYINPUT119), .B(KEYINPUT61), .Z(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(G155gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(KEYINPUT120), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n864_), .B(new_n867_), .ZN(G1346gat));
  INV_X1    g667(.A(G162gat), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n861_), .A2(new_n869_), .A3(new_n576_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n588_), .B1(new_n854_), .B2(new_n857_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n869_), .B2(new_n871_), .ZN(G1347gat));
  OR2_X1    g671(.A1(new_n804_), .A2(new_n814_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n398_), .A2(new_n304_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n345_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n873_), .A2(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(KEYINPUT121), .B1(new_n877_), .B2(new_n542_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT121), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n873_), .A2(new_n879_), .A3(new_n697_), .A4(new_n876_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n878_), .A2(G169gat), .A3(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT62), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NAND4_X1  g682(.A1(new_n878_), .A2(KEYINPUT62), .A3(G169gat), .A4(new_n880_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n877_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n885_), .A2(new_n697_), .A3(new_n235_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n883_), .A2(new_n884_), .A3(new_n886_), .ZN(G1348gat));
  OAI21_X1  g686(.A(new_n238_), .B1(new_n877_), .B2(new_n692_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n889_));
  OR2_X1    g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n889_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n818_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n892_));
  OAI211_X1 g691(.A(KEYINPUT57), .B(new_n583_), .C1(new_n799_), .C2(new_n800_), .ZN(new_n893_));
  OR2_X1    g692(.A1(new_n780_), .A2(new_n786_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n892_), .A2(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n610_), .B1(new_n896_), .B2(new_n819_), .ZN(new_n897_));
  OAI211_X1 g696(.A(KEYINPUT123), .B(new_n346_), .C1(new_n897_), .C2(new_n814_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n899_), .B1(new_n855_), .B2(new_n345_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n875_), .A2(new_n238_), .A3(new_n692_), .ZN(new_n902_));
  AOI22_X1  g701(.A1(new_n890_), .A2(new_n891_), .B1(new_n901_), .B2(new_n902_), .ZN(G1349gat));
  NOR2_X1   g702(.A1(new_n875_), .A2(new_n616_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n232_), .B1(new_n901_), .B2(new_n904_), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n616_), .A2(new_n266_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n877_), .A2(new_n906_), .ZN(new_n907_));
  OAI21_X1  g706(.A(KEYINPUT124), .B1(new_n905_), .B2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n909_));
  INV_X1    g708(.A(new_n904_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n910_), .B1(new_n898_), .B2(new_n900_), .ZN(new_n911_));
  OAI221_X1 g710(.A(new_n909_), .B1(new_n877_), .B2(new_n906_), .C1(new_n911_), .C2(new_n232_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n908_), .A2(new_n912_), .ZN(G1350gat));
  OAI21_X1  g712(.A(G190gat), .B1(new_n877_), .B2(new_n588_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n576_), .A2(new_n255_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n877_), .B2(new_n915_), .ZN(G1351gat));
  NOR4_X1   g715(.A1(new_n304_), .A2(new_n370_), .A3(new_n396_), .A4(new_n346_), .ZN(new_n917_));
  AND2_X1   g716(.A1(new_n826_), .A2(new_n917_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n918_), .A2(G197gat), .A3(new_n697_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT125), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n919_), .A2(new_n920_), .ZN(new_n922_));
  AOI21_X1  g721(.A(G197gat), .B1(new_n918_), .B2(new_n697_), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n921_), .A2(new_n922_), .A3(new_n923_), .ZN(G1352gat));
  NAND2_X1  g723(.A1(new_n826_), .A2(new_n917_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n925_), .A2(new_n692_), .ZN(new_n926_));
  AND2_X1   g725(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n927_));
  NOR2_X1   g726(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n926_), .B1(new_n927_), .B2(new_n928_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n929_), .B1(new_n926_), .B2(new_n928_), .ZN(G1353gat));
  INV_X1    g729(.A(KEYINPUT63), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n610_), .B1(new_n931_), .B2(new_n596_), .ZN(new_n932_));
  XOR2_X1   g731(.A(new_n932_), .B(KEYINPUT127), .Z(new_n933_));
  NAND2_X1  g732(.A1(new_n918_), .A2(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n931_), .A2(new_n596_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n934_), .B(new_n935_), .ZN(G1354gat));
  OR3_X1    g735(.A1(new_n925_), .A2(G218gat), .A3(new_n583_), .ZN(new_n937_));
  OAI21_X1  g736(.A(G218gat), .B1(new_n925_), .B2(new_n588_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n937_), .A2(new_n938_), .ZN(G1355gat));
endmodule


