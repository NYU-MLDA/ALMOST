//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 1 1 0 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n635_,
    new_n636_, new_n637_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n690_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n842_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n866_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n874_, new_n875_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_;
  NAND2_X1  g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT77), .B(G176gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT76), .ZN(new_n204_));
  INV_X1    g003(.A(G169gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n204_), .B1(new_n205_), .B2(KEYINPUT22), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT22), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n207_), .A2(KEYINPUT76), .A3(G169gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT75), .B1(new_n207_), .B2(G169gat), .ZN(new_n209_));
  NAND4_X1  g008(.A1(new_n203_), .A2(new_n206_), .A3(new_n208_), .A4(new_n209_), .ZN(new_n210_));
  NOR3_X1   g009(.A1(new_n207_), .A2(KEYINPUT75), .A3(G169gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n202_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT78), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT73), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT73), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(G183gat), .A3(G190gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(new_n218_), .A3(KEYINPUT23), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT23), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n215_), .A2(new_n220_), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  OR2_X1    g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  OAI211_X1 g023(.A(KEYINPUT78), .B(new_n202_), .C1(new_n210_), .C2(new_n211_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n214_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n216_), .A2(new_n218_), .A3(new_n220_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n215_), .A2(KEYINPUT23), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT72), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT72), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n215_), .A2(new_n230_), .A3(KEYINPUT23), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n227_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n232_));
  OR3_X1    g031(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT74), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT71), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT25), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n237_), .B1(new_n238_), .B2(G183gat), .ZN(new_n239_));
  XOR2_X1   g038(.A(KEYINPUT25), .B(G183gat), .Z(new_n240_));
  AOI21_X1  g039(.A(new_n239_), .B1(new_n240_), .B2(new_n237_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT26), .B(G190gat), .ZN(new_n242_));
  XOR2_X1   g041(.A(G169gat), .B(G176gat), .Z(new_n243_));
  AOI22_X1  g042(.A1(new_n241_), .A2(new_n242_), .B1(KEYINPUT24), .B2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n232_), .A2(KEYINPUT74), .A3(new_n233_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n236_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n226_), .A2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT30), .ZN(new_n248_));
  INV_X1    g047(.A(G120gat), .ZN(new_n249_));
  INV_X1    g048(.A(G127gat), .ZN(new_n250_));
  INV_X1    g049(.A(G134gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(G113gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G127gat), .A2(G134gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n253_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n249_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n257_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n259_), .A2(G120gat), .A3(new_n255_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  OR2_X1    g060(.A1(new_n248_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n248_), .A2(new_n261_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G15gat), .B(G43gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT31), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  AND3_X1   g065(.A1(new_n262_), .A2(new_n263_), .A3(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n266_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G71gat), .B(G99gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G227gat), .A2(G233gat), .ZN(new_n270_));
  XOR2_X1   g069(.A(new_n269_), .B(new_n270_), .Z(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  OR3_X1    g071(.A1(new_n267_), .A2(new_n268_), .A3(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n272_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT80), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT3), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n279_));
  OAI22_X1  g078(.A1(new_n278_), .A2(new_n279_), .B1(G141gat), .B2(G148gat), .ZN(new_n280_));
  AND3_X1   g079(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n281_));
  AOI21_X1  g080(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(G141gat), .A2(G148gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n284_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n280_), .A2(new_n283_), .A3(new_n285_), .ZN(new_n286_));
  XOR2_X1   g085(.A(G155gat), .B(G162gat), .Z(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT79), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n284_), .A2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT79), .B1(G141gat), .B2(G148gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n293_));
  AND4_X1   g092(.A1(new_n289_), .A2(new_n291_), .A3(new_n292_), .A4(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT1), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n287_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n288_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(new_n261_), .ZN(new_n299_));
  AOI22_X1  g098(.A1(new_n286_), .A2(new_n287_), .B1(new_n294_), .B2(new_n296_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n300_), .A2(new_n260_), .A3(new_n258_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n299_), .A2(new_n301_), .A3(KEYINPUT4), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT4), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n298_), .A2(new_n303_), .A3(new_n261_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT92), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G225gat), .A2(G233gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n298_), .A2(KEYINPUT92), .A3(new_n303_), .A4(new_n261_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n302_), .A2(new_n306_), .A3(new_n308_), .A4(new_n309_), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n299_), .A2(new_n301_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n307_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G1gat), .B(G29gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G57gat), .B(G85gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n310_), .A2(new_n312_), .A3(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n317_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n320_));
  OR3_X1    g119(.A1(new_n319_), .A2(KEYINPUT98), .A3(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT98), .B1(new_n319_), .B2(new_n320_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT86), .ZN(new_n324_));
  XOR2_X1   g123(.A(KEYINPUT85), .B(KEYINPUT29), .Z(new_n325_));
  XOR2_X1   g124(.A(G211gat), .B(G218gat), .Z(new_n326_));
  INV_X1    g125(.A(G197gat), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n327_), .A2(G204gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT83), .B(G197gat), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n328_), .B1(new_n329_), .B2(G204gat), .ZN(new_n330_));
  XOR2_X1   g129(.A(KEYINPUT84), .B(KEYINPUT21), .Z(new_n331_));
  AOI21_X1  g130(.A(new_n326_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(G204gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n329_), .A2(new_n333_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n334_), .B(KEYINPUT21), .C1(new_n327_), .C2(new_n333_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n332_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n326_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n330_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT21), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n298_), .A2(new_n325_), .B1(new_n336_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT82), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(G233gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n341_), .A2(G233gat), .ZN(new_n344_));
  OAI21_X1  g143(.A(G228gat), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n324_), .B1(new_n340_), .B2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n298_), .A2(KEYINPUT81), .A3(KEYINPUT29), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT81), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT29), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n348_), .B1(new_n300_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n336_), .A2(new_n339_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n347_), .A2(new_n350_), .A3(new_n345_), .A4(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n345_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n325_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n300_), .A2(new_n354_), .ZN(new_n355_));
  AOI22_X1  g154(.A1(new_n332_), .A2(new_n335_), .B1(new_n338_), .B2(KEYINPUT21), .ZN(new_n356_));
  OAI211_X1 g155(.A(KEYINPUT86), .B(new_n353_), .C1(new_n355_), .C2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n346_), .A2(new_n352_), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT87), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n346_), .A2(new_n352_), .A3(KEYINPUT87), .A4(new_n357_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(KEYINPUT28), .B1(new_n298_), .B2(KEYINPUT29), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT28), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n300_), .A2(new_n364_), .A3(new_n349_), .ZN(new_n365_));
  XOR2_X1   g164(.A(G22gat), .B(G50gat), .Z(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n363_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n367_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n362_), .A2(new_n371_), .ZN(new_n372_));
  XOR2_X1   g171(.A(G78gat), .B(G106gat), .Z(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n361_), .A2(new_n370_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n372_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n370_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n375_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n373_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n376_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n275_), .A2(new_n323_), .A3(new_n381_), .ZN(new_n382_));
  XOR2_X1   g181(.A(G8gat), .B(G36gat), .Z(new_n383_));
  XNOR2_X1  g182(.A(G64gat), .B(G92gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n385_), .B(new_n386_), .Z(new_n387_));
  NAND2_X1  g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT19), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT97), .ZN(new_n391_));
  INV_X1    g190(.A(new_n240_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n242_), .ZN(new_n393_));
  OR2_X1    g192(.A1(KEYINPUT88), .A2(KEYINPUT24), .ZN(new_n394_));
  NAND2_X1  g193(.A1(KEYINPUT88), .A2(KEYINPUT24), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n243_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n395_), .ZN(new_n397_));
  INV_X1    g196(.A(G176gat), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n397_), .A2(new_n205_), .A3(new_n398_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n393_), .A2(new_n222_), .A3(new_n396_), .A4(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n232_), .A2(new_n223_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT22), .B(G169gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n203_), .A2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n401_), .A2(new_n202_), .A3(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n356_), .A2(new_n400_), .A3(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT96), .B(KEYINPUT20), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n391_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n356_), .B1(new_n226_), .B2(new_n246_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n405_), .A2(new_n391_), .A3(new_n406_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n390_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT20), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n404_), .A2(new_n400_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n412_), .B1(new_n413_), .B2(new_n351_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n226_), .A2(new_n246_), .A3(new_n356_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n416_), .A2(new_n389_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n387_), .B1(new_n411_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n387_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n408_), .A2(new_n412_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n420_), .A2(new_n390_), .A3(new_n405_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT89), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n422_), .B1(new_n416_), .B2(new_n389_), .ZN(new_n423_));
  AOI211_X1 g222(.A(KEYINPUT89), .B(new_n390_), .C1(new_n414_), .C2(new_n415_), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n419_), .B(new_n421_), .C1(new_n423_), .C2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n418_), .A2(KEYINPUT27), .A3(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT99), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT99), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n418_), .A2(new_n428_), .A3(KEYINPUT27), .A4(new_n425_), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n421_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n387_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT91), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(new_n433_), .A3(new_n425_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT27), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n431_), .A2(KEYINPUT91), .A3(new_n387_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n434_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n430_), .A2(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n382_), .A2(new_n438_), .ZN(new_n439_));
  AOI22_X1  g238(.A1(new_n376_), .A2(new_n379_), .B1(new_n322_), .B2(new_n321_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n440_), .A2(new_n437_), .A3(new_n427_), .A4(new_n429_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT100), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n430_), .A2(KEYINPUT100), .A3(new_n440_), .A4(new_n437_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n434_), .A2(new_n436_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n302_), .A2(new_n306_), .A3(new_n307_), .A4(new_n309_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n311_), .A2(new_n308_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n317_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n318_), .A2(KEYINPUT33), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n318_), .A2(KEYINPUT33), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n450_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(KEYINPUT94), .B1(new_n445_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT94), .ZN(new_n456_));
  AOI211_X1 g255(.A(new_n456_), .B(new_n453_), .C1(new_n434_), .C2(new_n436_), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n419_), .A2(KEYINPUT32), .ZN(new_n458_));
  OR3_X1    g257(.A1(new_n431_), .A2(KEYINPUT95), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n417_), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n405_), .A2(new_n391_), .A3(new_n406_), .ZN(new_n461_));
  NOR3_X1   g260(.A1(new_n461_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n460_), .B1(new_n462_), .B2(new_n390_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n320_), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n463_), .A2(new_n458_), .B1(new_n464_), .B2(new_n318_), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT95), .B1(new_n431_), .B2(new_n458_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n459_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n455_), .A2(new_n457_), .A3(new_n468_), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n443_), .B(new_n444_), .C1(new_n469_), .C2(new_n380_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n275_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n439_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(KEYINPUT68), .B(G22gat), .Z(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(G15gat), .ZN(new_n474_));
  INV_X1    g273(.A(G1gat), .ZN(new_n475_));
  INV_X1    g274(.A(G8gat), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT14), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT68), .B(G22gat), .ZN(new_n478_));
  INV_X1    g277(.A(G15gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n474_), .A2(new_n477_), .A3(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT69), .ZN(new_n482_));
  XOR2_X1   g281(.A(G1gat), .B(G8gat), .Z(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n482_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n482_), .A2(new_n484_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G57gat), .B(G64gat), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n489_), .A2(KEYINPUT11), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(KEYINPUT11), .ZN(new_n491_));
  XOR2_X1   g290(.A(G71gat), .B(G78gat), .Z(new_n492_));
  NAND3_X1  g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n491_), .A2(new_n492_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G231gat), .A2(G233gat), .ZN(new_n496_));
  XOR2_X1   g295(.A(new_n495_), .B(new_n496_), .Z(new_n497_));
  XNOR2_X1  g296(.A(new_n488_), .B(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT16), .B(G183gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(G211gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G127gat), .B(G155gat), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n500_), .B(new_n501_), .Z(new_n502_));
  INV_X1    g301(.A(KEYINPUT17), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n502_), .A2(new_n503_), .ZN(new_n505_));
  NOR3_X1   g304(.A1(new_n498_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n506_), .B1(new_n504_), .B2(new_n498_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G230gat), .A2(G233gat), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G99gat), .A2(G106gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT6), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n513_));
  OR3_X1    g312(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n512_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(G85gat), .B(G92gat), .Z(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT8), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n515_), .A2(KEYINPUT8), .A3(new_n516_), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT9), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT64), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n522_), .A2(KEYINPUT64), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n516_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(KEYINPUT10), .B(G99gat), .Z(new_n526_));
  INV_X1    g325(.A(G106gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n522_), .A2(KEYINPUT64), .A3(G85gat), .A4(G92gat), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n525_), .A2(new_n528_), .A3(new_n529_), .A4(new_n512_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n521_), .A2(new_n530_), .A3(new_n495_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n519_), .A2(new_n530_), .A3(new_n520_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n495_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n531_), .A2(new_n534_), .A3(KEYINPUT12), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT12), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n532_), .A2(new_n536_), .A3(new_n533_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n510_), .B1(new_n535_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n531_), .A2(new_n534_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n510_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G120gat), .B(G148gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(new_n333_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT5), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(new_n398_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n542_), .A2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n539_), .A2(new_n541_), .A3(new_n546_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT13), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G113gat), .B(G141gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(new_n205_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(new_n327_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(KEYINPUT65), .B(G43gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(G50gat), .ZN(new_n556_));
  XOR2_X1   g355(.A(G29gat), .B(G36gat), .Z(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT15), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n488_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G229gat), .A2(G233gat), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n558_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n560_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n561_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n558_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n487_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n565_), .B1(new_n566_), .B2(new_n485_), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n486_), .A2(new_n558_), .A3(new_n487_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n564_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n563_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT70), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n554_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n554_), .ZN(new_n573_));
  AOI211_X1 g372(.A(KEYINPUT70), .B(new_n573_), .C1(new_n563_), .C2(new_n569_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n551_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G190gat), .B(G218gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(G134gat), .ZN(new_n579_));
  INV_X1    g378(.A(G162gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n582_), .A2(KEYINPUT36), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n559_), .A2(new_n532_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G232gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT34), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT35), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n521_), .A2(new_n530_), .A3(new_n558_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n584_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n587_), .A2(new_n588_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n592_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n584_), .A2(new_n594_), .A3(new_n589_), .A4(new_n590_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n583_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n582_), .A2(KEYINPUT36), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(KEYINPUT67), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT66), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n593_), .A2(new_n599_), .A3(new_n583_), .A4(new_n595_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n593_), .A2(new_n583_), .A3(new_n595_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT66), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n598_), .A2(new_n600_), .A3(new_n602_), .ZN(new_n603_));
  AOI22_X1  g402(.A1(new_n596_), .A2(new_n597_), .B1(KEYINPUT67), .B2(KEYINPUT37), .ZN(new_n604_));
  OAI21_X1  g403(.A(KEYINPUT37), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n601_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NOR4_X1   g407(.A1(new_n472_), .A2(new_n508_), .A3(new_n577_), .A4(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n323_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n609_), .A2(new_n475_), .A3(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n472_), .A2(new_n577_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n596_), .A2(new_n597_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n601_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n617_), .A2(new_n508_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n614_), .A2(new_n618_), .ZN(new_n619_));
  OAI21_X1  g418(.A(G1gat), .B1(new_n619_), .B2(new_n323_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n613_), .A2(new_n620_), .ZN(G1324gat));
  NAND3_X1  g420(.A1(new_n614_), .A2(new_n618_), .A3(new_n438_), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n622_), .A2(KEYINPUT103), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(KEYINPUT103), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n623_), .A2(G8gat), .A3(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(KEYINPUT104), .B(KEYINPUT39), .Z(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n609_), .A2(new_n476_), .A3(new_n438_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT102), .Z(new_n630_));
  NAND2_X1  g429(.A1(new_n625_), .A2(new_n627_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n628_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT40), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(G1325gat));
  OAI21_X1  g433(.A(G15gat), .B1(new_n619_), .B2(new_n471_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT41), .Z(new_n636_));
  NAND3_X1  g435(.A1(new_n609_), .A2(new_n479_), .A3(new_n275_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(G1326gat));
  INV_X1    g437(.A(G22gat), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n609_), .A2(new_n639_), .A3(new_n380_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G22gat), .B1(new_n619_), .B2(new_n381_), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n641_), .A2(KEYINPUT105), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(KEYINPUT105), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n642_), .A2(KEYINPUT42), .A3(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(KEYINPUT42), .B1(new_n642_), .B2(new_n643_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n640_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT106), .ZN(G1327gat));
  INV_X1    g446(.A(G29gat), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n616_), .A2(new_n507_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n614_), .A2(new_n648_), .A3(new_n610_), .A4(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n651_));
  OAI211_X1 g450(.A(KEYINPUT107), .B(new_n651_), .C1(new_n472_), .C2(new_n607_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n455_), .A2(new_n457_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n380_), .B1(new_n653_), .B2(new_n467_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n443_), .A2(new_n444_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n471_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n439_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n651_), .A2(KEYINPUT107), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n651_), .A2(KEYINPUT107), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n658_), .A2(new_n608_), .A3(new_n659_), .A4(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT108), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n577_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n652_), .A2(new_n661_), .A3(new_n508_), .A4(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n662_), .A2(new_n663_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n667_), .A2(new_n610_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n650_), .B1(new_n668_), .B2(new_n648_), .ZN(G1328gat));
  INV_X1    g468(.A(G36gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n670_), .B1(new_n667_), .B2(new_n438_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n614_), .A2(new_n649_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n438_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n672_), .A2(G36gat), .A3(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT45), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n671_), .A2(new_n675_), .ZN(new_n676_));
  XOR2_X1   g475(.A(KEYINPUT109), .B(KEYINPUT46), .Z(new_n677_));
  OAI21_X1  g476(.A(KEYINPUT110), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(KEYINPUT46), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT110), .ZN(new_n680_));
  INV_X1    g479(.A(new_n677_), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n680_), .B(new_n681_), .C1(new_n671_), .C2(new_n675_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n678_), .A2(new_n679_), .A3(new_n682_), .ZN(G1329gat));
  NAND3_X1  g482(.A1(new_n667_), .A2(G43gat), .A3(new_n275_), .ZN(new_n684_));
  INV_X1    g483(.A(G43gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n685_), .B1(new_n672_), .B2(new_n471_), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT111), .Z(new_n687_));
  NAND2_X1  g486(.A1(new_n684_), .A2(new_n687_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT47), .ZN(G1330gat));
  AND2_X1   g488(.A1(new_n667_), .A2(new_n380_), .ZN(new_n690_));
  INV_X1    g489(.A(G50gat), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n380_), .A2(new_n691_), .ZN(new_n692_));
  OAI22_X1  g491(.A1(new_n690_), .A2(new_n691_), .B1(new_n672_), .B2(new_n692_), .ZN(G1331gat));
  NOR2_X1   g492(.A1(new_n472_), .A2(new_n576_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n551_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n694_), .A2(new_n618_), .A3(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(G57gat), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n696_), .A2(new_n697_), .A3(new_n323_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n694_), .B(KEYINPUT112), .ZN(new_n699_));
  AND4_X1   g498(.A1(new_n507_), .A2(new_n699_), .A3(new_n695_), .A4(new_n607_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n610_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n698_), .B1(new_n701_), .B2(new_n697_), .ZN(G1332gat));
  INV_X1    g501(.A(G64gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n700_), .A2(new_n703_), .A3(new_n438_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G64gat), .B1(new_n696_), .B2(new_n673_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT48), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT113), .Z(G1333gat));
  NOR2_X1   g507(.A1(new_n471_), .A2(G71gat), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT114), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n700_), .A2(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(G71gat), .B1(new_n696_), .B2(new_n471_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT49), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1334gat));
  INV_X1    g513(.A(G78gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n700_), .A2(new_n715_), .A3(new_n380_), .ZN(new_n716_));
  OAI21_X1  g515(.A(G78gat), .B1(new_n696_), .B2(new_n381_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT50), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(G1335gat));
  AND2_X1   g518(.A1(new_n699_), .A2(new_n695_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(new_n610_), .A3(new_n649_), .ZN(new_n721_));
  INV_X1    g520(.A(G85gat), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT115), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n723_), .B(new_n724_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n652_), .A2(new_n661_), .A3(new_n508_), .A4(new_n695_), .ZN(new_n726_));
  OR3_X1    g525(.A1(new_n726_), .A2(KEYINPUT116), .A3(new_n576_), .ZN(new_n727_));
  OAI21_X1  g526(.A(KEYINPUT116), .B1(new_n726_), .B2(new_n576_), .ZN(new_n728_));
  AOI211_X1 g527(.A(new_n722_), .B(new_n323_), .C1(new_n727_), .C2(new_n728_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n725_), .A2(new_n729_), .ZN(G1336gat));
  NAND2_X1  g529(.A1(new_n720_), .A2(new_n649_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n731_), .A2(new_n673_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n732_), .A2(G92gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n673_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(G92gat), .B2(new_n734_), .ZN(G1337gat));
  NAND2_X1  g534(.A1(new_n275_), .A2(new_n526_), .ZN(new_n736_));
  INV_X1    g535(.A(G99gat), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n726_), .A2(new_n576_), .A3(new_n471_), .ZN(new_n738_));
  OAI22_X1  g537(.A1(new_n731_), .A2(new_n736_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g539(.A(KEYINPUT52), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n726_), .A2(new_n576_), .A3(new_n381_), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n742_), .A2(KEYINPUT117), .A3(new_n527_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT117), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n652_), .A2(new_n661_), .A3(new_n508_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n745_), .A2(new_n695_), .A3(new_n575_), .A4(new_n380_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n744_), .B1(new_n746_), .B2(G106gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n741_), .B1(new_n743_), .B2(new_n747_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n720_), .A2(new_n527_), .A3(new_n380_), .A4(new_n649_), .ZN(new_n749_));
  OAI21_X1  g548(.A(KEYINPUT117), .B1(new_n742_), .B2(new_n527_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n746_), .A2(new_n744_), .A3(G106gat), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(new_n751_), .A3(KEYINPUT52), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n748_), .A2(new_n749_), .A3(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT53), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT53), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n748_), .A2(new_n755_), .A3(new_n749_), .A4(new_n752_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(G1339gat));
  NAND3_X1  g556(.A1(new_n535_), .A2(new_n510_), .A3(new_n537_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT118), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n758_), .A2(new_n759_), .A3(KEYINPUT55), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n758_), .B2(KEYINPUT55), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n538_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n758_), .A2(KEYINPUT55), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT118), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n758_), .A2(new_n759_), .A3(KEYINPUT55), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n764_), .A2(new_n539_), .A3(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n762_), .A2(new_n766_), .A3(new_n547_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT56), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n762_), .A2(new_n766_), .A3(KEYINPUT56), .A4(new_n547_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n560_), .A2(new_n564_), .A3(new_n562_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n561_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n554_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n570_), .A2(new_n573_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT119), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT119), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n775_), .A2(new_n776_), .A3(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n771_), .A2(new_n549_), .A3(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT58), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n771_), .A2(KEYINPUT58), .A3(new_n549_), .A4(new_n781_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n784_), .A2(new_n608_), .A3(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n549_), .B1(new_n572_), .B2(new_n574_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n787_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n788_));
  AOI22_X1  g587(.A1(new_n778_), .A2(new_n780_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n616_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT57), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  OAI211_X1 g591(.A(KEYINPUT57), .B(new_n616_), .C1(new_n788_), .C2(new_n789_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n786_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n508_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n607_), .A2(new_n507_), .A3(new_n551_), .A4(new_n575_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT54), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n471_), .A2(new_n380_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n438_), .A2(new_n323_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n798_), .A2(new_n799_), .A3(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(G113gat), .B1(new_n801_), .B2(new_n576_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT59), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n798_), .A2(new_n803_), .A3(new_n799_), .A4(new_n800_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT121), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n801_), .A2(KEYINPUT121), .A3(new_n803_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n798_), .A2(new_n799_), .A3(new_n800_), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n808_), .A2(KEYINPUT120), .A3(KEYINPUT59), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT120), .B1(new_n808_), .B2(KEYINPUT59), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n806_), .B(new_n807_), .C1(new_n809_), .C2(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n811_), .A2(new_n575_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n802_), .B1(new_n812_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g612(.A(KEYINPUT122), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n811_), .B2(new_n551_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n810_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n808_), .A2(KEYINPUT120), .A3(KEYINPUT59), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n804_), .B(KEYINPUT121), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n818_), .A2(new_n819_), .A3(KEYINPUT122), .A4(new_n695_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n815_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(G120gat), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT60), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n551_), .B2(G120gat), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n801_), .B(new_n824_), .C1(new_n823_), .C2(G120gat), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n822_), .A2(new_n825_), .ZN(G1341gat));
  AOI21_X1  g625(.A(G127gat), .B1(new_n801_), .B2(new_n507_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n811_), .A2(new_n250_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n827_), .B1(new_n828_), .B2(new_n507_), .ZN(G1342gat));
  NAND4_X1  g628(.A1(new_n818_), .A2(new_n819_), .A3(G134gat), .A4(new_n608_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n251_), .B1(new_n808_), .B2(new_n616_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT123), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n830_), .A2(KEYINPUT123), .A3(new_n831_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(G1343gat));
  NOR2_X1   g635(.A1(new_n275_), .A2(new_n381_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n798_), .A2(new_n800_), .A3(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n576_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n695_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g642(.A1(new_n838_), .A2(new_n508_), .ZN(new_n844_));
  XOR2_X1   g643(.A(KEYINPUT61), .B(G155gat), .Z(new_n845_));
  XNOR2_X1  g644(.A(new_n844_), .B(new_n845_), .ZN(G1346gat));
  NOR3_X1   g645(.A1(new_n838_), .A2(new_n580_), .A3(new_n607_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n839_), .A2(new_n617_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n847_), .B1(new_n580_), .B2(new_n848_), .ZN(G1347gat));
  NOR2_X1   g648(.A1(new_n673_), .A2(new_n610_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n798_), .A2(new_n576_), .A3(new_n799_), .A4(new_n850_), .ZN(new_n851_));
  OR2_X1    g650(.A1(new_n851_), .A2(KEYINPUT124), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(KEYINPUT124), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(G169gat), .A3(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT62), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n798_), .A2(new_n850_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n857_), .A2(new_n799_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n858_), .A2(new_n576_), .A3(new_n402_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n852_), .A2(KEYINPUT62), .A3(G169gat), .A4(new_n853_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n856_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(KEYINPUT125), .ZN(G1348gat));
  NAND2_X1  g661(.A1(new_n858_), .A2(new_n695_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(new_n398_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n864_), .B1(new_n203_), .B2(new_n863_), .ZN(G1349gat));
  NAND2_X1  g664(.A1(new_n858_), .A2(new_n507_), .ZN(new_n866_));
  MUX2_X1   g665(.A(new_n392_), .B(G183gat), .S(new_n866_), .Z(G1350gat));
  NAND3_X1  g666(.A1(new_n858_), .A2(new_n617_), .A3(new_n242_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n858_), .A2(new_n608_), .ZN(new_n869_));
  INV_X1    g668(.A(G190gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n868_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT126), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n871_), .B(new_n872_), .ZN(G1351gat));
  NAND2_X1  g672(.A1(new_n857_), .A2(new_n837_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n874_), .A2(new_n575_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(new_n327_), .ZN(G1352gat));
  NOR2_X1   g675(.A1(new_n874_), .A2(new_n551_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(new_n333_), .ZN(G1353gat));
  INV_X1    g677(.A(KEYINPUT127), .ZN(new_n879_));
  INV_X1    g678(.A(new_n874_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n507_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n879_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n884_));
  INV_X1    g683(.A(new_n882_), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n880_), .A2(new_n507_), .A3(new_n884_), .A4(new_n885_), .ZN(new_n886_));
  MUX2_X1   g685(.A(new_n879_), .B(new_n883_), .S(new_n886_), .Z(G1354gat));
  AND3_X1   g686(.A1(new_n880_), .A2(G218gat), .A3(new_n608_), .ZN(new_n888_));
  AOI21_X1  g687(.A(G218gat), .B1(new_n880_), .B2(new_n617_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n888_), .A2(new_n889_), .ZN(G1355gat));
endmodule


