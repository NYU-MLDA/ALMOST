//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n797_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n919_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n929_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n956_, new_n957_, new_n958_, new_n960_,
    new_n961_, new_n962_, new_n964_, new_n965_, new_n966_, new_n968_,
    new_n969_, new_n970_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n977_, new_n978_;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT94), .Z(new_n203_));
  INV_X1    g002(.A(G228gat), .ZN(new_n204_));
  INV_X1    g003(.A(G233gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G197gat), .A2(G204gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT90), .B(G204gat), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n208_), .B1(new_n209_), .B2(G197gat), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n210_), .A2(KEYINPUT21), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G211gat), .B(G218gat), .ZN(new_n212_));
  XOR2_X1   g011(.A(KEYINPUT90), .B(G204gat), .Z(new_n213_));
  INV_X1    g012(.A(G197gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT21), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n216_), .B1(G197gat), .B2(G204gat), .ZN(new_n217_));
  AND3_X1   g016(.A1(new_n215_), .A2(KEYINPUT91), .A3(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(KEYINPUT91), .B1(new_n215_), .B2(new_n217_), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n211_), .B(new_n212_), .C1(new_n218_), .C2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT92), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n216_), .B1(new_n212_), .B2(new_n221_), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n210_), .B(new_n222_), .C1(new_n221_), .C2(new_n212_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n220_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G155gat), .A2(G162gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT87), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT3), .ZN(new_n231_));
  INV_X1    g030(.A(G141gat), .ZN(new_n232_));
  INV_X1    g031(.A(G148gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT2), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G141gat), .A2(G148gat), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n234_), .B(new_n235_), .C1(new_n236_), .C2(new_n237_), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n225_), .B(new_n227_), .C1(new_n230_), .C2(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n226_), .B1(KEYINPUT1), .B2(new_n225_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n240_), .B1(KEYINPUT1), .B2(new_n225_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n232_), .A2(new_n233_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n241_), .A2(new_n237_), .A3(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n239_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT88), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT88), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n239_), .A2(new_n246_), .A3(new_n243_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT29), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n207_), .B(new_n224_), .C1(new_n248_), .C2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n244_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n251_), .A2(new_n249_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n224_), .A2(KEYINPUT93), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT93), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n220_), .A2(new_n254_), .A3(new_n223_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n252_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n203_), .B(new_n250_), .C1(new_n256_), .C2(new_n207_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT96), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n248_), .A2(new_n249_), .ZN(new_n260_));
  XOR2_X1   g059(.A(G22gat), .B(G50gat), .Z(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n263_));
  INV_X1    g062(.A(new_n261_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n248_), .A2(new_n249_), .A3(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n262_), .A2(new_n263_), .A3(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n263_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n264_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n268_));
  AOI211_X1 g067(.A(KEYINPUT29), .B(new_n261_), .C1(new_n245_), .C2(new_n247_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n267_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n266_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  AND3_X1   g071(.A1(new_n220_), .A2(new_n254_), .A3(new_n223_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n254_), .B1(new_n220_), .B2(new_n223_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n206_), .B1(new_n275_), .B2(new_n252_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n276_), .A2(KEYINPUT96), .A3(new_n203_), .A4(new_n250_), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n259_), .A2(new_n272_), .A3(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n250_), .B1(new_n256_), .B2(new_n207_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT95), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n276_), .A2(KEYINPUT95), .A3(new_n250_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n281_), .A2(new_n282_), .A3(new_n202_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n203_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n279_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(new_n257_), .ZN(new_n286_));
  AOI22_X1  g085(.A1(new_n278_), .A2(new_n283_), .B1(new_n286_), .B2(new_n271_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n224_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(G169gat), .A2(G176gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT82), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT83), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n291_), .A2(KEYINPUT24), .A3(new_n294_), .ZN(new_n295_));
  AND2_X1   g094(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n296_));
  NOR2_X1   g095(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n297_));
  OAI21_X1  g096(.A(G183gat), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n298_), .A2(KEYINPUT81), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(KEYINPUT81), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT26), .B(G190gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT25), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n302_), .B1(new_n303_), .B2(G183gat), .ZN(new_n304_));
  OAI211_X1 g103(.A(KEYINPUT84), .B(new_n295_), .C1(new_n301_), .C2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT84), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n304_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n295_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n306_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G183gat), .A2(G190gat), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT23), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n291_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT24), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n314_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n305_), .A2(new_n309_), .A3(new_n317_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n312_), .B(new_n313_), .C1(G183gat), .C2(G190gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT22), .B(G169gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n319_), .B(new_n294_), .C1(new_n321_), .C2(G176gat), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n288_), .B1(new_n318_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G226gat), .A2(G233gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT19), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n291_), .A2(KEYINPUT24), .A3(new_n292_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT25), .B(G183gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n302_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n310_), .A2(KEYINPUT23), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n311_), .A2(G183gat), .A3(G190gat), .ZN(new_n331_));
  AOI22_X1  g130(.A1(new_n330_), .A2(new_n331_), .B1(new_n316_), .B2(new_n289_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n327_), .A2(KEYINPUT97), .A3(new_n329_), .A4(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n327_), .A2(new_n329_), .A3(new_n332_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT97), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n294_), .A2(KEYINPUT98), .ZN(new_n337_));
  INV_X1    g136(.A(G176gat), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n320_), .A2(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n292_), .B(KEYINPUT83), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT98), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n319_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(KEYINPUT99), .B1(new_n340_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT99), .ZN(new_n346_));
  NOR4_X1   g145(.A1(new_n343_), .A2(new_n337_), .A3(new_n346_), .A4(new_n339_), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n333_), .B(new_n336_), .C1(new_n345_), .C2(new_n347_), .ZN(new_n348_));
  OAI211_X1 g147(.A(KEYINPUT20), .B(new_n326_), .C1(new_n348_), .C2(new_n224_), .ZN(new_n349_));
  OR2_X1    g148(.A1(new_n323_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT20), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n351_), .B1(new_n348_), .B2(new_n224_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n288_), .A2(new_n318_), .A3(new_n322_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n325_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G8gat), .B(G36gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT18), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G64gat), .B(G92gat), .ZN(new_n358_));
  XOR2_X1   g157(.A(new_n357_), .B(new_n358_), .Z(new_n359_));
  NAND3_X1  g158(.A1(new_n350_), .A2(new_n355_), .A3(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n359_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n323_), .A2(new_n349_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n326_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n361_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n360_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT27), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n340_), .A2(new_n344_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(new_n334_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n253_), .A2(new_n255_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT100), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(new_n372_), .A3(KEYINPUT20), .ZN(new_n373_));
  INV_X1    g172(.A(new_n323_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n372_), .B1(new_n371_), .B2(KEYINPUT20), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n325_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n352_), .A2(new_n353_), .A3(new_n326_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT101), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  OAI211_X1 g179(.A(KEYINPUT101), .B(new_n325_), .C1(new_n375_), .C2(new_n376_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n359_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n360_), .A2(KEYINPUT102), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n362_), .A2(new_n363_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT102), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n384_), .A2(new_n385_), .A3(new_n359_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n383_), .A2(KEYINPUT27), .A3(new_n386_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n287_), .B(new_n367_), .C1(new_n382_), .C2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n318_), .A2(KEYINPUT30), .A3(new_n322_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(KEYINPUT30), .B1(new_n318_), .B2(new_n322_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT86), .ZN(new_n393_));
  INV_X1    g192(.A(new_n391_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n389_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT86), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n393_), .A2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G71gat), .B(G99gat), .ZN(new_n399_));
  INV_X1    g198(.A(G43gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G227gat), .A2(G233gat), .ZN(new_n402_));
  XOR2_X1   g201(.A(new_n401_), .B(new_n402_), .Z(new_n403_));
  XOR2_X1   g202(.A(KEYINPUT85), .B(G15gat), .Z(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n398_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n393_), .A2(new_n405_), .ZN(new_n408_));
  XOR2_X1   g207(.A(G127gat), .B(G134gat), .Z(new_n409_));
  XOR2_X1   g208(.A(G113gat), .B(G120gat), .Z(new_n410_));
  XOR2_X1   g209(.A(new_n409_), .B(new_n410_), .Z(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(KEYINPUT31), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n407_), .A2(new_n408_), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n412_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n405_), .B1(new_n393_), .B2(new_n397_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n395_), .A2(new_n396_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n416_), .A2(new_n406_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n414_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n413_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n245_), .A2(new_n247_), .A3(new_n411_), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n244_), .A2(new_n411_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT4), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G225gat), .A2(G233gat), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n420_), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n423_), .B(new_n425_), .C1(new_n426_), .C2(KEYINPUT4), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n422_), .A2(new_n424_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G1gat), .B(G29gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(G85gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(KEYINPUT0), .B(G57gat), .ZN(new_n432_));
  XOR2_X1   g231(.A(new_n431_), .B(new_n432_), .Z(new_n433_));
  NAND2_X1  g232(.A1(new_n429_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n433_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n427_), .A2(new_n435_), .A3(new_n428_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n419_), .A2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n388_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n359_), .A2(KEYINPUT32), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n381_), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n273_), .A2(new_n274_), .A3(new_n369_), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT100), .B1(new_n444_), .B2(new_n351_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(new_n374_), .A3(new_n373_), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n446_), .A2(new_n325_), .B1(KEYINPUT101), .B2(new_n378_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n442_), .B1(new_n443_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n384_), .A2(new_n441_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n436_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n435_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n449_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT33), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n451_), .B(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n420_), .A2(new_n421_), .A3(new_n425_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n426_), .A2(KEYINPUT4), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n457_), .B1(KEYINPUT4), .B2(new_n422_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n435_), .B(new_n456_), .C1(new_n458_), .C2(new_n425_), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n459_), .A2(new_n360_), .A3(new_n364_), .ZN(new_n460_));
  AOI22_X1  g259(.A1(new_n448_), .A2(new_n453_), .B1(new_n455_), .B2(new_n460_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n283_), .A2(new_n272_), .A3(new_n277_), .A4(new_n259_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n286_), .A2(new_n271_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n367_), .B1(new_n382_), .B2(new_n387_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n438_), .ZN(new_n466_));
  OAI22_X1  g265(.A1(new_n461_), .A2(new_n464_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n419_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n440_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G1gat), .B(G8gat), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  OR2_X1    g270(.A1(KEYINPUT76), .A2(G15gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(KEYINPUT76), .A2(G15gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(G22gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n472_), .A2(G22gat), .A3(new_n473_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT14), .ZN(new_n479_));
  XNOR2_X1  g278(.A(KEYINPUT77), .B(G1gat), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n479_), .B1(new_n480_), .B2(G8gat), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n471_), .B1(new_n478_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(G8gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT14), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n484_), .A2(new_n477_), .A3(new_n476_), .A4(new_n470_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n482_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G29gat), .B(G36gat), .Z(new_n488_));
  XNOR2_X1  g287(.A(G43gat), .B(G50gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n487_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT79), .ZN(new_n492_));
  INV_X1    g291(.A(new_n490_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n486_), .A2(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n492_), .B1(new_n494_), .B2(KEYINPUT78), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n490_), .B1(new_n482_), .B2(new_n485_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT78), .ZN(new_n497_));
  NOR3_X1   g296(.A1(new_n496_), .A2(new_n497_), .A3(KEYINPUT79), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n491_), .B1(new_n495_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G229gat), .A2(G233gat), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n494_), .A2(KEYINPUT78), .A3(new_n492_), .ZN(new_n502_));
  OAI21_X1  g301(.A(KEYINPUT79), .B1(new_n496_), .B2(new_n497_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n502_), .A2(new_n503_), .A3(new_n487_), .A4(new_n490_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n499_), .A2(new_n501_), .A3(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n490_), .B(KEYINPUT15), .Z(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(new_n487_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n507_), .A2(new_n500_), .A3(new_n494_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G113gat), .B(G141gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G169gat), .B(G197gat), .ZN(new_n510_));
  XOR2_X1   g309(.A(new_n509_), .B(new_n510_), .Z(new_n511_));
  AND3_X1   g310(.A1(new_n505_), .A2(new_n508_), .A3(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n511_), .B1(new_n505_), .B2(new_n508_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n469_), .A2(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(G120gat), .B(G148gat), .Z(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT72), .ZN(new_n517_));
  XOR2_X1   g316(.A(G176gat), .B(G204gat), .Z(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n519_), .B(new_n520_), .Z(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(G230gat), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n523_), .A2(new_n205_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G99gat), .A2(G106gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT6), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT6), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n527_), .A2(G99gat), .A3(G106gat), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n526_), .A2(new_n528_), .A3(KEYINPUT66), .ZN(new_n529_));
  AOI21_X1  g328(.A(KEYINPUT66), .B1(new_n526_), .B2(new_n528_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT7), .ZN(new_n531_));
  INV_X1    g330(.A(G99gat), .ZN(new_n532_));
  INV_X1    g331(.A(G106gat), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NOR3_X1   g335(.A1(new_n529_), .A2(new_n530_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT67), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G85gat), .A2(G92gat), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(G85gat), .A2(G92gat), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n538_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(G85gat), .ZN(new_n543_));
  INV_X1    g342(.A(G92gat), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n545_), .A2(KEYINPUT67), .A3(new_n539_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n542_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT8), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(KEYINPUT68), .B1(new_n537_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT66), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n527_), .B1(G99gat), .B2(G106gat), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n525_), .A2(KEYINPUT6), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n551_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n526_), .A2(new_n528_), .A3(KEYINPUT66), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n534_), .A2(new_n535_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n554_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT68), .ZN(new_n558_));
  AOI21_X1  g357(.A(KEYINPUT8), .B1(new_n542_), .B2(new_n546_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n557_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n552_), .A2(new_n553_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n547_), .B1(new_n561_), .B2(new_n536_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT8), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n550_), .A2(new_n560_), .A3(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(KEYINPUT69), .B(G71gat), .ZN(new_n565_));
  INV_X1    g364(.A(G78gat), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n566_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(G64gat), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(G57gat), .ZN(new_n571_));
  INV_X1    g370(.A(G57gat), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(G64gat), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n571_), .A2(new_n573_), .A3(KEYINPUT11), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n569_), .A2(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(KEYINPUT11), .B1(new_n571_), .B2(new_n573_), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n567_), .B(new_n568_), .C1(new_n577_), .C2(new_n574_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT9), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n539_), .A2(KEYINPUT65), .A3(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT65), .B1(new_n539_), .B2(new_n581_), .ZN(new_n583_));
  OAI221_X1 g382(.A(new_n545_), .B1(new_n581_), .B2(new_n539_), .C1(new_n582_), .C2(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(KEYINPUT10), .B(G99gat), .Z(new_n585_));
  XOR2_X1   g384(.A(KEYINPUT64), .B(G106gat), .Z(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n584_), .A2(new_n555_), .A3(new_n554_), .A4(new_n587_), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n564_), .A2(new_n580_), .A3(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n580_), .B1(new_n564_), .B2(new_n588_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n524_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(KEYINPUT70), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT70), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n593_), .B(new_n524_), .C1(new_n589_), .C2(new_n590_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n557_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n558_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n556_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n548_), .B1(new_n598_), .B2(new_n547_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n596_), .A2(new_n597_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n588_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n579_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n564_), .A2(new_n580_), .A3(new_n588_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n602_), .A2(KEYINPUT12), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT12), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n590_), .A2(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n524_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n522_), .B1(new_n595_), .B2(new_n607_), .ZN(new_n608_));
  NOR3_X1   g407(.A1(new_n589_), .A2(new_n590_), .A3(new_n605_), .ZN(new_n609_));
  AOI211_X1 g408(.A(KEYINPUT12), .B(new_n580_), .C1(new_n564_), .C2(new_n588_), .ZN(new_n610_));
  OAI22_X1  g409(.A1(new_n609_), .A2(new_n610_), .B1(new_n523_), .B2(new_n205_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n611_), .A2(new_n594_), .A3(new_n592_), .A4(new_n521_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(KEYINPUT73), .B(KEYINPUT13), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n608_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n608_), .A2(new_n612_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n614_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(G127gat), .B(G155gat), .Z(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT16), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G183gat), .B(G211gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT17), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G231gat), .A2(G233gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n486_), .B(new_n623_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n624_), .A2(new_n579_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n579_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n622_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n624_), .A2(new_n579_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT17), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n621_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n624_), .A2(new_n579_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n628_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n627_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT37), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n506_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n635_));
  XOR2_X1   g434(.A(KEYINPUT74), .B(KEYINPUT34), .Z(new_n636_));
  NAND2_X1  g435(.A1(G232gat), .A2(G233gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n638_), .A2(KEYINPUT35), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n564_), .A2(new_n493_), .A3(new_n588_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n635_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n638_), .A2(KEYINPUT35), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT75), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n635_), .A2(new_n642_), .A3(new_n639_), .A4(new_n640_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n644_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT36), .ZN(new_n648_));
  XNOR2_X1  g447(.A(G190gat), .B(G218gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(G134gat), .B(G162gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n647_), .A2(new_n648_), .A3(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n644_), .A2(new_n651_), .A3(new_n646_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n648_), .B1(new_n647_), .B2(new_n652_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n634_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n656_), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n658_), .A2(KEYINPUT37), .A3(new_n654_), .A4(new_n653_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n515_), .A2(new_n617_), .A3(new_n633_), .A4(new_n660_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n661_), .A2(new_n438_), .A3(new_n480_), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n662_), .A2(KEYINPUT38), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(KEYINPUT38), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n655_), .A2(new_n656_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n469_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n617_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n668_), .A2(new_n514_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n667_), .A2(new_n633_), .A3(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G1gat), .B1(new_n670_), .B2(new_n438_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n663_), .A2(new_n664_), .A3(new_n671_), .ZN(G1324gat));
  NAND2_X1  g471(.A1(new_n380_), .A2(new_n381_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(new_n361_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n387_), .ZN(new_n675_));
  AOI22_X1  g474(.A1(new_n674_), .A2(new_n675_), .B1(new_n366_), .B2(new_n365_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G8gat), .B1(new_n670_), .B2(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT39), .ZN(new_n678_));
  OR3_X1    g477(.A1(new_n661_), .A2(G8gat), .A3(new_n676_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT40), .Z(G1325gat));
  NOR3_X1   g480(.A1(new_n661_), .A2(G15gat), .A3(new_n468_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT103), .Z(new_n683_));
  OAI21_X1  g482(.A(G15gat), .B1(new_n670_), .B2(new_n468_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT41), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n684_), .A2(KEYINPUT41), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n683_), .A2(new_n685_), .A3(new_n686_), .ZN(G1326gat));
  OAI21_X1  g486(.A(G22gat), .B1(new_n670_), .B2(new_n287_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT42), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n464_), .A2(new_n475_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT104), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n689_), .B1(new_n661_), .B2(new_n691_), .ZN(G1327gat));
  INV_X1    g491(.A(new_n440_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n437_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n360_), .A2(new_n364_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n434_), .A2(new_n454_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n451_), .A2(KEYINPUT33), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n695_), .A2(new_n696_), .A3(new_n459_), .A4(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n441_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n698_), .B1(new_n699_), .B2(new_n452_), .ZN(new_n700_));
  AOI22_X1  g499(.A1(new_n676_), .A2(new_n694_), .B1(new_n700_), .B2(new_n287_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n693_), .B1(new_n701_), .B2(new_n419_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n514_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n633_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n666_), .A2(new_n704_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n705_), .A2(new_n668_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n702_), .A2(new_n703_), .A3(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT105), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n515_), .A2(KEYINPUT105), .A3(new_n706_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(G29gat), .B1(new_n711_), .B2(new_n437_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT43), .ZN(new_n713_));
  INV_X1    g512(.A(new_n660_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n702_), .B2(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n452_), .B1(new_n673_), .B2(new_n442_), .ZN(new_n716_));
  AND4_X1   g515(.A1(new_n695_), .A2(new_n696_), .A3(new_n459_), .A4(new_n697_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n287_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n694_), .B(new_n367_), .C1(new_n382_), .C2(new_n387_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n419_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n713_), .B(new_n714_), .C1(new_n720_), .C2(new_n440_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n704_), .B(new_n669_), .C1(new_n715_), .C2(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT44), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n437_), .A2(G29gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n712_), .B1(new_n724_), .B2(new_n725_), .ZN(G1328gat));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n676_), .A2(G36gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n709_), .A2(new_n710_), .A3(new_n728_), .ZN(new_n729_));
  XOR2_X1   g528(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n709_), .A2(new_n710_), .A3(new_n728_), .A4(new_n730_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n723_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n723_), .A2(new_n735_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n736_), .A2(new_n465_), .A3(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n734_), .B1(new_n738_), .B2(G36gat), .ZN(new_n739_));
  XNOR2_X1  g538(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n727_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n740_), .ZN(new_n742_));
  INV_X1    g541(.A(G36gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n724_), .B2(new_n465_), .ZN(new_n744_));
  OAI211_X1 g543(.A(KEYINPUT108), .B(new_n742_), .C1(new_n744_), .C2(new_n734_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n739_), .A2(KEYINPUT46), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n741_), .A2(new_n745_), .A3(new_n746_), .ZN(G1329gat));
  AOI21_X1  g546(.A(G43gat), .B1(new_n711_), .B2(new_n419_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n468_), .A2(new_n400_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n724_), .B2(new_n749_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g550(.A(G50gat), .B1(new_n711_), .B2(new_n464_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n464_), .A2(G50gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n724_), .B2(new_n753_), .ZN(G1331gat));
  NOR2_X1   g553(.A1(new_n469_), .A2(new_n703_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n755_), .A2(new_n668_), .A3(new_n633_), .A4(new_n660_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(G57gat), .B1(new_n757_), .B2(new_n437_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n505_), .A2(new_n508_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n511_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n505_), .A2(new_n508_), .A3(new_n511_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n761_), .A2(new_n633_), .A3(new_n762_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n617_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n667_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n572_), .B1(new_n437_), .B2(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n768_), .B1(new_n767_), .B2(new_n572_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n758_), .B1(new_n766_), .B2(new_n769_), .ZN(G1332gat));
  OAI21_X1  g569(.A(G64gat), .B1(new_n765_), .B2(new_n676_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT48), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n757_), .A2(new_n570_), .A3(new_n465_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(G1333gat));
  OAI21_X1  g573(.A(G71gat), .B1(new_n765_), .B2(new_n468_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n775_), .B(new_n776_), .ZN(new_n777_));
  OR2_X1    g576(.A1(new_n468_), .A2(G71gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n756_), .B2(new_n778_), .ZN(G1334gat));
  OAI21_X1  g578(.A(G78gat), .B1(new_n765_), .B2(new_n287_), .ZN(new_n780_));
  XOR2_X1   g579(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n781_));
  XNOR2_X1  g580(.A(new_n780_), .B(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n464_), .A2(new_n566_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT112), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n782_), .B1(new_n756_), .B2(new_n784_), .ZN(G1335gat));
  NOR2_X1   g584(.A1(new_n705_), .A2(new_n617_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n755_), .A2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n543_), .B1(new_n787_), .B2(new_n438_), .ZN(new_n788_));
  XOR2_X1   g587(.A(new_n788_), .B(KEYINPUT113), .Z(new_n789_));
  NOR3_X1   g588(.A1(new_n617_), .A2(new_n703_), .A3(new_n633_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(KEYINPUT43), .B1(new_n469_), .B2(new_n660_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(new_n721_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n794_), .A2(new_n543_), .A3(new_n438_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n789_), .A2(new_n795_), .ZN(G1336gat));
  OAI21_X1  g595(.A(G92gat), .B1(new_n794_), .B2(new_n676_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n787_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(new_n544_), .A3(new_n465_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n799_), .ZN(G1337gat));
  OAI21_X1  g599(.A(G99gat), .B1(new_n794_), .B2(new_n468_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n798_), .A2(new_n419_), .A3(new_n585_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g603(.A1(new_n798_), .A2(new_n464_), .A3(new_n586_), .ZN(new_n805_));
  AOI211_X1 g604(.A(KEYINPUT52), .B(new_n533_), .C1(new_n793_), .C2(new_n464_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n464_), .B(new_n790_), .C1(new_n715_), .C2(new_n722_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n807_), .B1(new_n808_), .B2(G106gat), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n805_), .B1(new_n806_), .B2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT115), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n812_), .B(new_n805_), .C1(new_n806_), .C2(new_n809_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n811_), .A2(new_n813_), .A3(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n814_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(G1339gat));
  NOR3_X1   g616(.A1(new_n595_), .A2(new_n607_), .A3(new_n522_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n514_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT55), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n589_), .A2(new_n590_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n610_), .B1(new_n822_), .B2(KEYINPUT12), .ZN(new_n823_));
  OAI211_X1 g622(.A(KEYINPUT118), .B(new_n821_), .C1(new_n823_), .C2(new_n524_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n825_), .B1(new_n607_), .B2(KEYINPUT55), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n607_), .A2(KEYINPUT55), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n823_), .A2(new_n524_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n824_), .A2(new_n826_), .A3(new_n827_), .A4(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n522_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT56), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n829_), .A2(KEYINPUT56), .A3(new_n522_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n820_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n499_), .A2(new_n500_), .A3(new_n504_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n496_), .A2(new_n500_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n511_), .B1(new_n507_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n762_), .A2(new_n838_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n615_), .A2(new_n839_), .ZN(new_n840_));
  OAI211_X1 g639(.A(KEYINPUT57), .B(new_n665_), .C1(new_n834_), .C2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT119), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n665_), .B1(new_n834_), .B2(new_n840_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n829_), .A2(KEYINPUT56), .A3(new_n522_), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT56), .B1(new_n829_), .B2(new_n522_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n819_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n840_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n851_), .A2(KEYINPUT119), .A3(KEYINPUT57), .A4(new_n665_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n818_), .A2(new_n839_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  OAI211_X1 g655(.A(KEYINPUT58), .B(new_n853_), .C1(new_n847_), .C2(new_n848_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n856_), .A2(new_n714_), .A3(new_n857_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n843_), .A2(new_n846_), .A3(new_n852_), .A4(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n704_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n763_), .A2(KEYINPUT116), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n514_), .A2(new_n862_), .A3(new_n633_), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n608_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n616_), .B1(new_n608_), .B2(new_n612_), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n861_), .B(new_n863_), .C1(new_n864_), .C2(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n660_), .B1(new_n866_), .B2(KEYINPUT117), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT117), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n862_), .B1(new_n514_), .B2(new_n633_), .ZN(new_n869_));
  AND4_X1   g668(.A1(new_n862_), .A2(new_n761_), .A3(new_n633_), .A4(new_n762_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n868_), .B1(new_n871_), .B2(new_n617_), .ZN(new_n872_));
  OAI21_X1  g671(.A(KEYINPUT54), .B1(new_n867_), .B2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n866_), .A2(KEYINPUT117), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n871_), .A2(new_n617_), .A3(new_n868_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n874_), .A2(new_n875_), .A3(new_n876_), .A4(new_n660_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n873_), .A2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n860_), .A2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(KEYINPUT120), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n860_), .A2(new_n882_), .A3(new_n879_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n883_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n388_), .A2(new_n468_), .A3(new_n438_), .ZN(new_n885_));
  XOR2_X1   g684(.A(new_n885_), .B(KEYINPUT121), .Z(new_n886_));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(G113gat), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n888_), .A2(new_n889_), .A3(new_n703_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n880_), .A2(new_n891_), .A3(new_n886_), .ZN(new_n892_));
  AOI211_X1 g691(.A(new_n514_), .B(new_n892_), .C1(new_n887_), .C2(KEYINPUT59), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n890_), .B1(new_n893_), .B2(new_n889_), .ZN(G1340gat));
  NOR2_X1   g693(.A1(new_n617_), .A2(KEYINPUT60), .ZN(new_n895_));
  INV_X1    g694(.A(G120gat), .ZN(new_n896_));
  MUX2_X1   g695(.A(KEYINPUT60), .B(new_n895_), .S(new_n896_), .Z(new_n897_));
  NAND3_X1  g696(.A1(new_n884_), .A2(new_n886_), .A3(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n898_), .B(new_n899_), .ZN(new_n900_));
  AOI211_X1 g699(.A(new_n617_), .B(new_n892_), .C1(new_n887_), .C2(KEYINPUT59), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n896_), .B2(new_n901_), .ZN(G1341gat));
  AOI21_X1  g701(.A(G127gat), .B1(new_n888_), .B2(new_n633_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n892_), .B1(new_n887_), .B2(KEYINPUT59), .ZN(new_n904_));
  INV_X1    g703(.A(G127gat), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n905_), .B1(new_n633_), .B2(KEYINPUT123), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n906_), .B1(KEYINPUT123), .B2(new_n905_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n903_), .B1(new_n904_), .B2(new_n907_), .ZN(G1342gat));
  AOI21_X1  g707(.A(G134gat), .B1(new_n888_), .B2(new_n666_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(KEYINPUT124), .B(G134gat), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n660_), .A2(new_n910_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n909_), .B1(new_n904_), .B2(new_n911_), .ZN(G1343gat));
  NOR3_X1   g711(.A1(new_n465_), .A2(new_n287_), .A3(new_n438_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n882_), .B1(new_n860_), .B2(new_n879_), .ZN(new_n914_));
  AOI211_X1 g713(.A(KEYINPUT120), .B(new_n878_), .C1(new_n859_), .C2(new_n704_), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n468_), .B(new_n913_), .C1(new_n914_), .C2(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(new_n514_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(new_n232_), .ZN(G1344gat));
  NOR2_X1   g717(.A1(new_n916_), .A2(new_n617_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(new_n233_), .ZN(G1345gat));
  AOI21_X1  g719(.A(new_n419_), .B1(new_n881_), .B2(new_n883_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT125), .ZN(new_n922_));
  NAND4_X1  g721(.A1(new_n921_), .A2(new_n922_), .A3(new_n633_), .A4(new_n913_), .ZN(new_n923_));
  OAI21_X1  g722(.A(KEYINPUT125), .B1(new_n916_), .B2(new_n704_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(KEYINPUT61), .B(G155gat), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n923_), .A2(new_n924_), .A3(new_n925_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n923_), .B2(new_n924_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n926_), .A2(new_n927_), .ZN(G1346gat));
  OAI21_X1  g727(.A(G162gat), .B1(new_n916_), .B2(new_n660_), .ZN(new_n929_));
  OR2_X1    g728(.A1(new_n665_), .A2(G162gat), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n916_), .B2(new_n930_), .ZN(G1347gat));
  NOR2_X1   g730(.A1(new_n676_), .A2(new_n439_), .ZN(new_n932_));
  INV_X1    g731(.A(new_n932_), .ZN(new_n933_));
  AOI211_X1 g732(.A(new_n464_), .B(new_n933_), .C1(new_n860_), .C2(new_n879_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(new_n703_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n935_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n936_), .B1(new_n321_), .B2(new_n935_), .ZN(new_n937_));
  AOI21_X1  g736(.A(KEYINPUT62), .B1(new_n935_), .B2(G169gat), .ZN(new_n938_));
  OR2_X1    g737(.A1(new_n937_), .A2(new_n938_), .ZN(G1348gat));
  NOR3_X1   g738(.A1(new_n933_), .A2(new_n338_), .A3(new_n617_), .ZN(new_n940_));
  AOI21_X1  g739(.A(KEYINPUT126), .B1(new_n884_), .B2(new_n287_), .ZN(new_n941_));
  OAI211_X1 g740(.A(KEYINPUT126), .B(new_n287_), .C1(new_n914_), .C2(new_n915_), .ZN(new_n942_));
  INV_X1    g741(.A(new_n942_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n940_), .B1(new_n941_), .B2(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n945_));
  AOI21_X1  g744(.A(G176gat), .B1(new_n934_), .B2(new_n668_), .ZN(new_n946_));
  INV_X1    g745(.A(new_n946_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n944_), .A2(new_n945_), .A3(new_n947_), .ZN(new_n948_));
  INV_X1    g747(.A(new_n940_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n287_), .B1(new_n914_), .B2(new_n915_), .ZN(new_n950_));
  INV_X1    g749(.A(KEYINPUT126), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n950_), .A2(new_n951_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n949_), .B1(new_n952_), .B2(new_n942_), .ZN(new_n953_));
  OAI21_X1  g752(.A(KEYINPUT127), .B1(new_n953_), .B2(new_n946_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n948_), .A2(new_n954_), .ZN(G1349gat));
  OAI211_X1 g754(.A(new_n633_), .B(new_n932_), .C1(new_n941_), .C2(new_n943_), .ZN(new_n956_));
  INV_X1    g755(.A(G183gat), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n704_), .A2(new_n328_), .ZN(new_n958_));
  AOI22_X1  g757(.A1(new_n956_), .A2(new_n957_), .B1(new_n934_), .B2(new_n958_), .ZN(G1350gat));
  NAND3_X1  g758(.A1(new_n934_), .A2(new_n302_), .A3(new_n666_), .ZN(new_n960_));
  AND2_X1   g759(.A1(new_n934_), .A2(new_n714_), .ZN(new_n961_));
  INV_X1    g760(.A(G190gat), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n960_), .B1(new_n961_), .B2(new_n962_), .ZN(G1351gat));
  NOR2_X1   g762(.A1(new_n676_), .A2(new_n466_), .ZN(new_n964_));
  NAND3_X1  g763(.A1(new_n884_), .A2(new_n468_), .A3(new_n964_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n965_), .A2(new_n514_), .ZN(new_n966_));
  XNOR2_X1  g765(.A(new_n966_), .B(new_n214_), .ZN(G1352gat));
  INV_X1    g766(.A(new_n965_), .ZN(new_n968_));
  AOI21_X1  g767(.A(G204gat), .B1(new_n968_), .B2(new_n668_), .ZN(new_n969_));
  NOR3_X1   g768(.A1(new_n965_), .A2(new_n213_), .A3(new_n617_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(new_n969_), .A2(new_n970_), .ZN(G1353gat));
  NOR2_X1   g770(.A1(new_n965_), .A2(new_n704_), .ZN(new_n972_));
  NOR2_X1   g771(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n973_));
  AND2_X1   g772(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n974_));
  OAI21_X1  g773(.A(new_n972_), .B1(new_n973_), .B2(new_n974_), .ZN(new_n975_));
  OAI21_X1  g774(.A(new_n975_), .B1(new_n972_), .B2(new_n973_), .ZN(G1354gat));
  OAI21_X1  g775(.A(G218gat), .B1(new_n965_), .B2(new_n660_), .ZN(new_n977_));
  OR2_X1    g776(.A1(new_n665_), .A2(G218gat), .ZN(new_n978_));
  OAI21_X1  g777(.A(new_n977_), .B1(new_n965_), .B2(new_n978_), .ZN(G1355gat));
endmodule


