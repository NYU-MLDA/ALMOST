//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n904_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n935_, new_n936_,
    new_n937_, new_n939_, new_n940_, new_n941_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n951_, new_n952_;
  INV_X1    g000(.A(KEYINPUT105), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT104), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G225gat), .A2(G233gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  OR2_X1    g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  AND2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT2), .ZN(new_n209_));
  AND3_X1   g008(.A1(KEYINPUT86), .A2(G141gat), .A3(G148gat), .ZN(new_n210_));
  AOI21_X1  g009(.A(KEYINPUT86), .B1(G141gat), .B2(G148gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n209_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT89), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT89), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n215_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n212_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n219_));
  INV_X1    g018(.A(G141gat), .ZN(new_n220_));
  INV_X1    g019(.A(G148gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT88), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .A4(KEYINPUT88), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n220_), .A2(new_n221_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT3), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n224_), .A2(new_n225_), .A3(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n208_), .B1(new_n218_), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT1), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n207_), .A2(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n231_), .B1(KEYINPUT87), .B2(new_n226_), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n210_), .A2(new_n211_), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n226_), .A2(KEYINPUT87), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n206_), .A2(new_n230_), .A3(new_n207_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .A4(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n229_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(G120gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(G113gat), .ZN(new_n239_));
  INV_X1    g038(.A(G113gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(G120gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT84), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n239_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n242_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n244_));
  OAI21_X1  g043(.A(G127gat), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n240_), .A2(G120gat), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n238_), .A2(G113gat), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT84), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(G127gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n239_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n245_), .A2(G134gat), .A3(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(G134gat), .B1(new_n245_), .B2(new_n251_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n237_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(G134gat), .ZN(new_n255_));
  NOR3_X1   g054(.A1(new_n243_), .A2(new_n244_), .A3(G127gat), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n249_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n255_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n245_), .A2(new_n251_), .A3(G134gat), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n258_), .A2(new_n229_), .A3(new_n236_), .A4(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n254_), .A2(new_n260_), .A3(KEYINPUT4), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n259_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n262_), .A2(KEYINPUT100), .A3(new_n263_), .A4(new_n237_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  AOI22_X1  g064(.A1(new_n258_), .A2(new_n259_), .B1(new_n229_), .B2(new_n236_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT100), .B1(new_n266_), .B2(new_n263_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n205_), .B(new_n261_), .C1(new_n265_), .C2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n254_), .A2(new_n260_), .A3(new_n204_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G1gat), .B(G29gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT0), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(G57gat), .ZN(new_n273_));
  OR2_X1    g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n273_), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n274_), .A2(G85gat), .A3(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(G85gat), .B1(new_n274_), .B2(new_n275_), .ZN(new_n277_));
  OR2_X1    g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n268_), .A2(new_n269_), .A3(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n278_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n280_));
  NOR3_X1   g079(.A1(new_n279_), .A2(new_n280_), .A3(KEYINPUT102), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n268_), .A2(KEYINPUT102), .A3(new_n269_), .A4(new_n278_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n203_), .B1(new_n281_), .B2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G15gat), .B(G43gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G71gat), .B(G99gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n258_), .A2(KEYINPUT31), .A3(new_n259_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(KEYINPUT31), .B1(new_n258_), .B2(new_n259_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n286_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT31), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n262_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n286_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n292_), .A2(new_n287_), .A3(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G227gat), .A2(G233gat), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n295_), .B(KEYINPUT83), .Z(new_n296_));
  AND3_X1   g095(.A1(new_n290_), .A2(new_n294_), .A3(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n296_), .B1(new_n290_), .B2(new_n294_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n285_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n290_), .A2(new_n294_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n296_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n285_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n290_), .A2(new_n294_), .A3(new_n296_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n302_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  NOR3_X1   g104(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n306_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT26), .B(G190gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT25), .B(G183gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT81), .B(KEYINPUT23), .ZN(new_n314_));
  INV_X1    g113(.A(G183gat), .ZN(new_n315_));
  INV_X1    g114(.A(G190gat), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n314_), .A2(new_n317_), .ZN(new_n318_));
  NOR3_X1   g117(.A1(new_n315_), .A2(new_n316_), .A3(KEYINPUT23), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n310_), .B(new_n313_), .C1(new_n318_), .C2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT22), .B(G169gat), .ZN(new_n321_));
  INV_X1    g120(.A(G176gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT82), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n321_), .A2(KEYINPUT82), .A3(new_n322_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT23), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n329_), .B1(G183gat), .B2(G190gat), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n330_), .B1(new_n314_), .B2(new_n317_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(G183gat), .A2(G190gat), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n309_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n320_), .B1(new_n328_), .B2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT30), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT85), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n299_), .A2(new_n305_), .A3(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n336_), .B1(new_n299_), .B2(new_n305_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n237_), .B(new_n263_), .C1(new_n252_), .C2(new_n253_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT100), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n342_), .A2(new_n264_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n261_), .A2(new_n205_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n269_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n278_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT102), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n268_), .A2(new_n269_), .A3(new_n278_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n347_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n350_), .A2(KEYINPUT104), .A3(new_n282_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n284_), .A2(new_n339_), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n237_), .A2(KEYINPUT29), .ZN(new_n353_));
  NOR2_X1   g152(.A1(G197gat), .A2(G204gat), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G197gat), .A2(G204gat), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n355_), .A2(KEYINPUT21), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT21), .ZN(new_n358_));
  INV_X1    g157(.A(new_n356_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n358_), .B1(new_n359_), .B2(new_n354_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G211gat), .B(G218gat), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n357_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n355_), .A2(KEYINPUT91), .A3(new_n356_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT91), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n364_), .B1(new_n359_), .B2(new_n354_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT92), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n361_), .A2(new_n358_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n366_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n367_), .B1(new_n366_), .B2(new_n368_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n362_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT90), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(G233gat), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n373_), .A2(G233gat), .ZN(new_n376_));
  OAI21_X1  g175(.A(G228gat), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n353_), .A2(new_n372_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n377_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n362_), .ZN(new_n380_));
  AOI21_X1  g179(.A(KEYINPUT91), .B1(new_n355_), .B2(new_n356_), .ZN(new_n381_));
  NOR3_X1   g180(.A1(new_n359_), .A2(new_n354_), .A3(new_n364_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n368_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT92), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n380_), .B1(new_n384_), .B2(new_n369_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT29), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n386_), .B1(new_n229_), .B2(new_n236_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n379_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G78gat), .B(G106gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n378_), .A2(new_n388_), .A3(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n390_), .B1(new_n378_), .B2(new_n388_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n391_), .B1(new_n392_), .B2(KEYINPUT93), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT93), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n378_), .A2(new_n388_), .A3(new_n394_), .A4(new_n390_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n229_), .A2(new_n386_), .A3(new_n236_), .ZN(new_n397_));
  XOR2_X1   g196(.A(G22gat), .B(G50gat), .Z(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT28), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n397_), .B(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(KEYINPUT94), .B1(new_n396_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT94), .ZN(new_n402_));
  INV_X1    g201(.A(new_n400_), .ZN(new_n403_));
  AOI211_X1 g202(.A(new_n402_), .B(new_n403_), .C1(new_n393_), .C2(new_n395_), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n401_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT20), .ZN(new_n406_));
  INV_X1    g205(.A(new_n309_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n407_), .A2(new_n307_), .ZN(new_n408_));
  NOR3_X1   g207(.A1(new_n331_), .A2(new_n408_), .A3(new_n306_), .ZN(new_n409_));
  OR2_X1    g208(.A1(new_n312_), .A2(KEYINPUT96), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n312_), .A2(KEYINPUT96), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(new_n311_), .A3(new_n411_), .ZN(new_n412_));
  OAI22_X1  g211(.A1(new_n318_), .A2(new_n319_), .B1(G183gat), .B2(G190gat), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n407_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n414_));
  AOI22_X1  g213(.A1(new_n409_), .A2(new_n412_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n406_), .B1(new_n385_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n334_), .A2(new_n372_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G226gat), .A2(G233gat), .ZN(new_n418_));
  XOR2_X1   g217(.A(new_n418_), .B(KEYINPUT19), .Z(new_n419_));
  NAND3_X1  g218(.A1(new_n416_), .A2(new_n417_), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT97), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n327_), .B(new_n309_), .C1(new_n331_), .C2(new_n332_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n385_), .A2(new_n423_), .A3(new_n320_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n409_), .A2(new_n412_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n413_), .A2(new_n414_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n372_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n424_), .A2(new_n428_), .A3(KEYINPUT20), .ZN(new_n429_));
  XOR2_X1   g228(.A(new_n419_), .B(KEYINPUT95), .Z(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n416_), .A2(new_n417_), .A3(KEYINPUT97), .A4(new_n419_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n422_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G64gat), .B(G92gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G8gat), .B(G36gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n433_), .A2(new_n439_), .ZN(new_n440_));
  AOI22_X1  g239(.A1(new_n421_), .A2(new_n420_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n441_), .A2(new_n432_), .A3(new_n438_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT27), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n416_), .A2(new_n417_), .ZN(new_n445_));
  OAI22_X1  g244(.A1(new_n445_), .A2(new_n419_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n444_), .B1(new_n446_), .B2(new_n439_), .ZN(new_n447_));
  AOI22_X1  g246(.A1(new_n443_), .A2(new_n444_), .B1(new_n442_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n392_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(new_n403_), .A3(new_n391_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n405_), .A2(new_n448_), .A3(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n202_), .B1(new_n352_), .B2(new_n451_), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n350_), .A2(KEYINPUT104), .A3(new_n282_), .ZN(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT104), .B1(new_n350_), .B2(new_n282_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n450_), .B1(new_n401_), .B2(new_n404_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n438_), .B1(new_n441_), .B2(new_n432_), .ZN(new_n457_));
  AND4_X1   g256(.A1(new_n432_), .A2(new_n422_), .A3(new_n431_), .A4(new_n438_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n444_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n447_), .A2(new_n442_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n456_), .A2(new_n461_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n455_), .A2(new_n462_), .A3(KEYINPUT105), .A4(new_n339_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n452_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n438_), .A2(KEYINPUT32), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n429_), .A2(new_n430_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n419_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n466_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n422_), .A2(new_n431_), .A3(new_n432_), .A4(new_n465_), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n350_), .A2(new_n282_), .A3(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT103), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n350_), .A2(KEYINPUT103), .A3(new_n282_), .A4(new_n471_), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT99), .B1(new_n457_), .B2(new_n458_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n349_), .A2(KEYINPUT33), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT33), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n268_), .A2(new_n478_), .A3(new_n269_), .A4(new_n278_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n254_), .A2(new_n260_), .A3(new_n205_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n278_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n261_), .A2(new_n204_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n482_), .B1(new_n343_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT101), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT101), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n482_), .B(new_n486_), .C1(new_n343_), .C2(new_n483_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT99), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n440_), .A2(new_n442_), .A3(new_n489_), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n476_), .A2(new_n480_), .A3(new_n488_), .A4(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n474_), .A2(new_n475_), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n456_), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n456_), .A2(new_n448_), .ZN(new_n494_));
  AOI22_X1  g293(.A1(new_n492_), .A2(new_n493_), .B1(new_n494_), .B2(new_n455_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n464_), .B1(new_n495_), .B2(new_n339_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G230gat), .A2(G233gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT64), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G71gat), .B(G78gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G57gat), .B(G64gat), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT67), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT11), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n499_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n500_), .B(KEYINPUT67), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT11), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(KEYINPUT11), .A3(new_n499_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT7), .ZN(new_n511_));
  INV_X1    g310(.A(G99gat), .ZN(new_n512_));
  INV_X1    g311(.A(G106gat), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n511_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G99gat), .A2(G106gat), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT66), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n519_), .A2(KEYINPUT6), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT6), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n521_), .A2(KEYINPUT66), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n518_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(KEYINPUT66), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n519_), .A2(KEYINPUT6), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n524_), .A2(new_n525_), .A3(new_n517_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n516_), .B1(new_n523_), .B2(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(G85gat), .B(G92gat), .Z(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT8), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT8), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n524_), .A2(new_n525_), .A3(new_n517_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n517_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n531_), .B(new_n528_), .C1(new_n534_), .C2(new_n516_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n530_), .A2(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n537_));
  XOR2_X1   g336(.A(KEYINPUT65), .B(G85gat), .Z(new_n538_));
  INV_X1    g337(.A(G92gat), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n537_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(KEYINPUT10), .B(G99gat), .Z(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n513_), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n542_), .B(new_n544_), .C1(new_n533_), .C2(new_n532_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n536_), .A2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n510_), .A2(new_n546_), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n536_), .A2(new_n545_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n548_), .A2(new_n509_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n498_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT68), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(KEYINPUT71), .B(KEYINPUT12), .Z(new_n553_));
  OAI21_X1  g352(.A(new_n553_), .B1(new_n548_), .B2(new_n509_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n547_), .A2(new_n498_), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n536_), .A2(KEYINPUT69), .A3(new_n545_), .ZN(new_n556_));
  AOI21_X1  g355(.A(KEYINPUT69), .B1(new_n536_), .B2(new_n545_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n507_), .A2(KEYINPUT12), .A3(new_n508_), .ZN(new_n559_));
  AOI21_X1  g358(.A(KEYINPUT70), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT69), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n546_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n536_), .A2(KEYINPUT69), .A3(new_n545_), .ZN(new_n563_));
  AND4_X1   g362(.A1(KEYINPUT70), .A2(new_n562_), .A3(new_n559_), .A4(new_n563_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n554_), .B(new_n555_), .C1(new_n560_), .C2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n552_), .A2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G120gat), .B(G148gat), .ZN(new_n567_));
  INV_X1    g366(.A(G204gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT5), .B(G176gat), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n569_), .B(new_n570_), .Z(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n566_), .A2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n552_), .A2(new_n565_), .A3(new_n571_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n573_), .A2(KEYINPUT13), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(KEYINPUT13), .B1(new_n573_), .B2(new_n574_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(G36gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(G29gat), .ZN(new_n581_));
  INV_X1    g380(.A(G29gat), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(G36gat), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n581_), .A2(new_n583_), .A3(KEYINPUT72), .ZN(new_n584_));
  AOI21_X1  g383(.A(KEYINPUT72), .B1(new_n581_), .B2(new_n583_), .ZN(new_n585_));
  OAI21_X1  g384(.A(G43gat), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n581_), .A2(new_n583_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT72), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(G43gat), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n581_), .A2(new_n583_), .A3(KEYINPUT72), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n589_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n586_), .A2(new_n592_), .A3(G50gat), .ZN(new_n593_));
  AOI21_X1  g392(.A(G50gat), .B1(new_n586_), .B2(new_n592_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G15gat), .B(G22gat), .ZN(new_n596_));
  INV_X1    g395(.A(G1gat), .ZN(new_n597_));
  INV_X1    g396(.A(G8gat), .ZN(new_n598_));
  OAI21_X1  g397(.A(KEYINPUT14), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G1gat), .B(G8gat), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n600_), .B(new_n601_), .Z(new_n602_));
  NAND2_X1  g401(.A1(new_n595_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G229gat), .A2(G233gat), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT77), .Z(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n603_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n602_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT15), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n593_), .A2(new_n594_), .A3(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n586_), .A2(new_n592_), .ZN(new_n611_));
  INV_X1    g410(.A(G50gat), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n586_), .A2(new_n592_), .A3(G50gat), .ZN(new_n614_));
  AOI21_X1  g413(.A(KEYINPUT15), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n608_), .B1(new_n610_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT76), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n609_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n613_), .A2(KEYINPUT15), .A3(new_n614_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(KEYINPUT76), .A3(new_n608_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n607_), .B1(new_n618_), .B2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n595_), .B(new_n602_), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n624_), .A2(G229gat), .A3(G233gat), .ZN(new_n625_));
  OAI21_X1  g424(.A(KEYINPUT80), .B1(new_n623_), .B2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G113gat), .B(G141gat), .ZN(new_n627_));
  INV_X1    g426(.A(G197gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(KEYINPUT79), .B(G169gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n632_), .A2(KEYINPUT78), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT80), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n624_), .A2(G229gat), .A3(G233gat), .ZN(new_n635_));
  AOI21_X1  g434(.A(KEYINPUT76), .B1(new_n621_), .B2(new_n608_), .ZN(new_n636_));
  AOI211_X1 g435(.A(new_n617_), .B(new_n602_), .C1(new_n619_), .C2(new_n620_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n634_), .B(new_n635_), .C1(new_n638_), .C2(new_n607_), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n626_), .A2(new_n633_), .A3(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n633_), .B1(new_n626_), .B2(new_n639_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n579_), .A2(new_n642_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n496_), .A2(new_n643_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n602_), .B(KEYINPUT75), .Z(new_n645_));
  NAND2_X1  g444(.A1(G231gat), .A2(G233gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(new_n510_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(G127gat), .B(G155gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT16), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(new_n315_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(G211gat), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT17), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n652_), .A2(new_n653_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n648_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n656_), .B1(new_n654_), .B2(new_n648_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT37), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n562_), .A2(new_n621_), .A3(new_n563_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(G232gat), .A2(G233gat), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT34), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n661_), .A2(KEYINPUT35), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n662_), .B1(new_n548_), .B2(new_n595_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n659_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n661_), .A2(KEYINPUT35), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(G190gat), .B(G218gat), .ZN(new_n667_));
  XNOR2_X1  g466(.A(G134gat), .B(G162gat), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(KEYINPUT73), .B(KEYINPUT36), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n666_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT74), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n666_), .A2(KEYINPUT74), .A3(new_n671_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n669_), .B(KEYINPUT36), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n666_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n658_), .B1(new_n676_), .B2(new_n679_), .ZN(new_n680_));
  AOI211_X1 g479(.A(KEYINPUT37), .B(new_n678_), .C1(new_n674_), .C2(new_n675_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n657_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n644_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n455_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n685_), .A2(new_n597_), .A3(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT38), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n643_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n657_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n678_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n496_), .A2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n692_), .A2(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(G1gat), .B1(new_n696_), .B2(new_n455_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n687_), .A2(new_n688_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n689_), .A2(new_n697_), .A3(new_n698_), .ZN(G1324gat));
  NAND3_X1  g498(.A1(new_n685_), .A2(new_n598_), .A3(new_n461_), .ZN(new_n700_));
  OAI21_X1  g499(.A(G8gat), .B1(new_n696_), .B2(new_n448_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n701_), .A2(KEYINPUT39), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(KEYINPUT39), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n700_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g504(.A(new_n339_), .ZN(new_n706_));
  OAI21_X1  g505(.A(G15gat), .B1(new_n696_), .B2(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT41), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n684_), .A2(G15gat), .A3(new_n706_), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1326gat));
  OAI21_X1  g509(.A(G22gat), .B1(new_n696_), .B2(new_n493_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT42), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n493_), .A2(G22gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n712_), .B1(new_n684_), .B2(new_n713_), .ZN(G1327gat));
  NOR2_X1   g513(.A1(new_n690_), .A2(new_n657_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n680_), .A2(new_n681_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n452_), .A2(new_n463_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n492_), .A2(new_n493_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n494_), .A2(new_n455_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n339_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n716_), .B(new_n717_), .C1(new_n718_), .C2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n496_), .B2(new_n717_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n715_), .B1(new_n723_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n715_), .B(KEYINPUT44), .C1(new_n723_), .C2(new_n726_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n730_), .A2(new_n455_), .A3(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n691_), .A2(new_n693_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT107), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n644_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n686_), .A2(new_n582_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT108), .ZN(new_n738_));
  OAI22_X1  g537(.A1(new_n733_), .A2(new_n582_), .B1(new_n736_), .B2(new_n738_), .ZN(G1328gat));
  NAND4_X1  g538(.A1(new_n644_), .A2(new_n580_), .A3(new_n461_), .A4(new_n735_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT45), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n448_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n742_));
  AOI211_X1 g541(.A(KEYINPUT109), .B(new_n580_), .C1(new_n742_), .C2(new_n731_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT109), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n729_), .A2(new_n461_), .A3(new_n731_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n745_), .B2(G36gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n741_), .B1(new_n743_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT46), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  OAI211_X1 g548(.A(KEYINPUT46), .B(new_n741_), .C1(new_n743_), .C2(new_n746_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1329gat));
  OAI21_X1  g550(.A(new_n590_), .B1(new_n736_), .B2(new_n706_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n729_), .A2(G43gat), .A3(new_n339_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n752_), .B1(new_n753_), .B2(new_n732_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g554(.A1(new_n730_), .A2(new_n612_), .A3(new_n493_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n644_), .A2(new_n456_), .A3(new_n735_), .ZN(new_n757_));
  AOI22_X1  g556(.A1(new_n756_), .A2(new_n731_), .B1(new_n612_), .B2(new_n757_), .ZN(G1331gat));
  INV_X1    g557(.A(new_n642_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n578_), .A2(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n695_), .A2(new_n657_), .A3(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(G57gat), .B1(new_n761_), .B2(new_n455_), .ZN(new_n762_));
  AND2_X1   g561(.A1(new_n496_), .A2(new_n760_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n683_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n686_), .A2(new_n273_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n762_), .B1(new_n764_), .B2(new_n765_), .ZN(G1332gat));
  OAI21_X1  g565(.A(G64gat), .B1(new_n761_), .B2(new_n448_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT48), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n448_), .A2(G64gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n768_), .B1(new_n764_), .B2(new_n769_), .ZN(G1333gat));
  OAI21_X1  g569(.A(G71gat), .B1(new_n761_), .B2(new_n706_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT49), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n706_), .A2(G71gat), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT110), .Z(new_n774_));
  OAI21_X1  g573(.A(new_n772_), .B1(new_n764_), .B2(new_n774_), .ZN(G1334gat));
  OAI21_X1  g574(.A(G78gat), .B1(new_n761_), .B2(new_n493_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n776_), .B(new_n777_), .ZN(new_n778_));
  OR2_X1    g577(.A1(new_n493_), .A2(G78gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n778_), .B1(new_n764_), .B2(new_n779_), .ZN(G1335gat));
  NAND2_X1  g579(.A1(new_n763_), .A2(new_n735_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(G85gat), .B1(new_n782_), .B2(new_n686_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n723_), .A2(new_n726_), .ZN(new_n784_));
  NOR4_X1   g583(.A1(new_n784_), .A2(new_n657_), .A3(new_n578_), .A4(new_n759_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n455_), .A2(new_n538_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n783_), .B1(new_n785_), .B2(new_n786_), .ZN(G1336gat));
  OAI21_X1  g586(.A(new_n539_), .B1(new_n781_), .B2(new_n448_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT112), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n448_), .A2(new_n539_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT113), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n789_), .B1(new_n785_), .B2(new_n791_), .ZN(G1337gat));
  NAND3_X1  g591(.A1(new_n782_), .A2(new_n543_), .A3(new_n339_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n578_), .A2(new_n657_), .A3(new_n759_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n339_), .B(new_n794_), .C1(new_n723_), .C2(new_n726_), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n795_), .A2(KEYINPUT114), .A3(G99gat), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT114), .B1(new_n795_), .B2(G99gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n793_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g598(.A1(new_n782_), .A2(new_n513_), .A3(new_n456_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(KEYINPUT115), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n456_), .B(new_n794_), .C1(new_n723_), .C2(new_n726_), .ZN(new_n802_));
  XOR2_X1   g601(.A(KEYINPUT116), .B(KEYINPUT52), .Z(new_n803_));
  AND3_X1   g602(.A1(new_n802_), .A2(G106gat), .A3(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n803_), .B1(new_n802_), .B2(G106gat), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n801_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT53), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n801_), .B(new_n808_), .C1(new_n804_), .C2(new_n805_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(G1339gat));
  XNOR2_X1  g609(.A(new_n693_), .B(new_n658_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n576_), .A2(new_n759_), .A3(new_n577_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n811_), .A2(new_n812_), .A3(new_n813_), .A4(new_n657_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n577_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n815_), .A2(new_n575_), .A3(new_n642_), .ZN(new_n816_));
  OAI21_X1  g615(.A(KEYINPUT54), .B1(new_n682_), .B2(new_n816_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n814_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n573_), .A2(new_n574_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n632_), .B(new_n635_), .C1(new_n638_), .C2(new_n607_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n603_), .B(new_n605_), .C1(new_n636_), .C2(new_n637_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n632_), .B1(new_n624_), .B2(new_n606_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT118), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n823_), .B(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n819_), .A2(new_n820_), .A3(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n574_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT117), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n829_), .B(new_n574_), .C1(new_n640_), .C2(new_n641_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n547_), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n554_), .B(new_n832_), .C1(new_n560_), .C2(new_n564_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n498_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n565_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n558_), .A2(KEYINPUT70), .A3(new_n559_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n562_), .A2(new_n559_), .A3(new_n563_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT70), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n837_), .A2(new_n840_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n841_), .A2(KEYINPUT55), .A3(new_n554_), .A4(new_n555_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n834_), .A2(new_n836_), .A3(new_n842_), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n843_), .A2(KEYINPUT56), .A3(new_n572_), .ZN(new_n844_));
  AOI21_X1  g643(.A(KEYINPUT56), .B1(new_n843_), .B2(new_n572_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n826_), .B1(new_n831_), .B2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n847_), .A2(KEYINPUT57), .A3(new_n694_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n825_), .A2(new_n574_), .A3(new_n820_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT58), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n849_), .B(KEYINPUT58), .C1(new_n844_), .C2(new_n845_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(new_n717_), .A3(new_n853_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n828_), .B(new_n830_), .C1(new_n845_), .C2(new_n844_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n693_), .B1(new_n855_), .B2(new_n826_), .ZN(new_n856_));
  XOR2_X1   g655(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n857_));
  OAI211_X1 g656(.A(new_n848_), .B(new_n854_), .C1(new_n856_), .C2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n818_), .B1(new_n858_), .B2(new_n691_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n455_), .A2(new_n706_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n462_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n859_), .A2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(G113gat), .B1(new_n862_), .B2(new_n759_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT120), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n863_), .B(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT59), .B1(new_n859_), .B2(new_n861_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n858_), .A2(new_n691_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n818_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT59), .ZN(new_n871_));
  INV_X1    g670(.A(new_n861_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n870_), .A2(new_n871_), .A3(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT121), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n862_), .A2(KEYINPUT121), .A3(new_n871_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n867_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n642_), .A2(new_n240_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n865_), .B1(new_n877_), .B2(new_n878_), .ZN(G1340gat));
  AOI21_X1  g678(.A(KEYINPUT60), .B1(new_n579_), .B2(new_n238_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n880_), .B1(KEYINPUT60), .B2(new_n238_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n862_), .A2(new_n881_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(KEYINPUT122), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n866_), .A2(new_n579_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n884_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n885_));
  OAI21_X1  g684(.A(G120gat), .B1(new_n885_), .B2(KEYINPUT123), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n866_), .A2(new_n579_), .ZN(new_n887_));
  AOI21_X1  g686(.A(KEYINPUT121), .B1(new_n862_), .B2(new_n871_), .ZN(new_n888_));
  NOR4_X1   g687(.A1(new_n859_), .A2(new_n874_), .A3(KEYINPUT59), .A4(new_n861_), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n887_), .B(KEYINPUT123), .C1(new_n888_), .C2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n883_), .B1(new_n886_), .B2(new_n891_), .ZN(G1341gat));
  NAND2_X1  g691(.A1(new_n877_), .A2(new_n657_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(G127gat), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n862_), .A2(new_n249_), .A3(new_n657_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1342gat));
  NAND2_X1  g695(.A1(new_n877_), .A2(new_n717_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(G134gat), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n862_), .A2(new_n255_), .A3(new_n693_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1343gat));
  NAND4_X1  g699(.A1(new_n870_), .A2(new_n686_), .A3(new_n494_), .A4(new_n706_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n901_), .A2(new_n642_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(new_n220_), .ZN(G1344gat));
  NOR2_X1   g702(.A1(new_n901_), .A2(new_n578_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(new_n221_), .ZN(G1345gat));
  NOR2_X1   g704(.A1(new_n901_), .A2(new_n691_), .ZN(new_n906_));
  XOR2_X1   g705(.A(KEYINPUT61), .B(G155gat), .Z(new_n907_));
  XNOR2_X1  g706(.A(new_n906_), .B(new_n907_), .ZN(G1346gat));
  OAI21_X1  g707(.A(G162gat), .B1(new_n901_), .B2(new_n811_), .ZN(new_n909_));
  OR2_X1    g708(.A1(new_n694_), .A2(G162gat), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n909_), .B1(new_n901_), .B2(new_n910_), .ZN(G1347gat));
  NOR3_X1   g710(.A1(new_n352_), .A2(new_n456_), .A3(new_n448_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n870_), .A2(new_n912_), .ZN(new_n913_));
  OAI211_X1 g712(.A(KEYINPUT62), .B(G169gat), .C1(new_n913_), .C2(new_n642_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT62), .ZN(new_n915_));
  INV_X1    g714(.A(new_n912_), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n859_), .A2(new_n642_), .A3(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(G169gat), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n915_), .B1(new_n917_), .B2(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n321_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n914_), .A2(new_n919_), .A3(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT124), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n921_), .B(new_n922_), .ZN(G1348gat));
  NOR2_X1   g722(.A1(new_n322_), .A2(KEYINPUT125), .ZN(new_n924_));
  XNOR2_X1  g723(.A(KEYINPUT125), .B(G176gat), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n913_), .A2(new_n578_), .ZN(new_n926_));
  MUX2_X1   g725(.A(new_n924_), .B(new_n925_), .S(new_n926_), .Z(G1349gat));
  INV_X1    g726(.A(new_n913_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n410_), .A2(new_n411_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n928_), .A2(new_n657_), .A3(new_n929_), .ZN(new_n930_));
  AND2_X1   g729(.A1(new_n930_), .A2(KEYINPUT126), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n930_), .A2(KEYINPUT126), .ZN(new_n932_));
  AOI21_X1  g731(.A(G183gat), .B1(new_n928_), .B2(new_n657_), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n931_), .A2(new_n932_), .A3(new_n933_), .ZN(G1350gat));
  OAI21_X1  g733(.A(G190gat), .B1(new_n913_), .B2(new_n811_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n693_), .A2(new_n311_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(KEYINPUT127), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n935_), .B1(new_n913_), .B2(new_n937_), .ZN(G1351gat));
  NOR4_X1   g737(.A1(new_n686_), .A2(new_n493_), .A3(new_n448_), .A4(new_n339_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n870_), .A2(new_n939_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n940_), .A2(new_n642_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(new_n628_), .ZN(G1352gat));
  NOR2_X1   g741(.A1(new_n940_), .A2(new_n578_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(new_n568_), .ZN(G1353gat));
  INV_X1    g743(.A(new_n940_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n945_), .A2(new_n657_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n947_));
  AND2_X1   g746(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n948_));
  NOR3_X1   g747(.A1(new_n946_), .A2(new_n947_), .A3(new_n948_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n949_), .B1(new_n946_), .B2(new_n947_), .ZN(G1354gat));
  OR3_X1    g749(.A1(new_n940_), .A2(G218gat), .A3(new_n694_), .ZN(new_n951_));
  OAI21_X1  g750(.A(G218gat), .B1(new_n940_), .B2(new_n811_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n951_), .A2(new_n952_), .ZN(G1355gat));
endmodule


