//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 1 1 0 1 1 1 1 0 0 1 1 0 0 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n632_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n824_, new_n825_,
    new_n827_, new_n828_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n835_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT72), .B(KEYINPUT73), .Z(new_n203_));
  XNOR2_X1  g002(.A(G43gat), .B(G50gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(G43gat), .B(G50gat), .Z(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G29gat), .B(G36gat), .ZN(new_n209_));
  AND3_X1   g008(.A1(new_n205_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n209_), .B1(new_n205_), .B2(new_n208_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G15gat), .B(G22gat), .ZN(new_n213_));
  INV_X1    g012(.A(G1gat), .ZN(new_n214_));
  INV_X1    g013(.A(G8gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT14), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G1gat), .B(G8gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n212_), .B(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G229gat), .A2(G233gat), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT82), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT15), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n225_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n205_), .A2(new_n208_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n209_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n205_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(KEYINPUT15), .A3(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n220_), .B1(new_n226_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT83), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n212_), .A2(new_n220_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n232_), .A2(new_n233_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n234_), .A2(new_n222_), .A3(new_n235_), .A4(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n221_), .A2(new_n223_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n224_), .B1(new_n239_), .B2(KEYINPUT82), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G169gat), .B(G197gat), .ZN(new_n241_));
  INV_X1    g040(.A(G141gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT84), .B(G113gat), .ZN(new_n244_));
  XOR2_X1   g043(.A(new_n243_), .B(new_n244_), .Z(new_n245_));
  AOI21_X1  g044(.A(new_n202_), .B1(new_n240_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT82), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n247_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n245_), .ZN(new_n249_));
  NOR4_X1   g048(.A1(new_n248_), .A2(KEYINPUT85), .A3(new_n224_), .A4(new_n249_), .ZN(new_n250_));
  OAI22_X1  g049(.A1(new_n246_), .A2(new_n250_), .B1(new_n240_), .B2(new_n245_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT7), .ZN(new_n252_));
  INV_X1    g051(.A(G99gat), .ZN(new_n253_));
  INV_X1    g052(.A(G106gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G99gat), .A2(G106gat), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT6), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n255_), .A2(new_n258_), .A3(new_n259_), .A4(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G85gat), .B(G92gat), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT8), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n267_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT69), .B1(new_n266_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n261_), .A2(new_n265_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT8), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n264_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n258_), .A2(new_n259_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n273_), .A2(KEYINPUT68), .A3(new_n260_), .A4(new_n255_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n272_), .A2(new_n274_), .A3(new_n275_), .A4(new_n267_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n269_), .A2(new_n271_), .A3(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT66), .B(G85gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(G92gat), .ZN(new_n279_));
  NOR2_X1   g078(.A1(G85gat), .A2(G92gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n279_), .B1(KEYINPUT67), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT9), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n281_), .B(new_n282_), .C1(KEYINPUT67), .C2(new_n279_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n265_), .A2(KEYINPUT67), .A3(KEYINPUT9), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT10), .B(G99gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT65), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(new_n254_), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n283_), .A2(new_n284_), .A3(new_n288_), .A4(new_n273_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n277_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n226_), .A2(new_n231_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT76), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n277_), .A2(new_n212_), .A3(new_n289_), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n292_), .A2(KEYINPUT74), .A3(new_n293_), .A4(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G232gat), .A2(G233gat), .ZN(new_n296_));
  XOR2_X1   g095(.A(new_n296_), .B(KEYINPUT34), .Z(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n294_), .A2(new_n293_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n297_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n299_), .A2(KEYINPUT74), .A3(new_n292_), .A4(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT35), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n299_), .A2(new_n303_), .A3(new_n292_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT75), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n298_), .A2(new_n301_), .A3(KEYINPUT35), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n306_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G190gat), .B(G218gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G134gat), .B(G162gat), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n310_), .B(new_n311_), .Z(new_n312_));
  NAND3_X1  g111(.A1(new_n309_), .A2(KEYINPUT36), .A3(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n312_), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n298_), .A2(new_n301_), .A3(KEYINPUT35), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n304_), .B1(new_n298_), .B2(new_n301_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n314_), .B1(new_n317_), .B2(new_n307_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n306_), .A2(new_n308_), .A3(new_n314_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT36), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  OAI211_X1 g120(.A(KEYINPUT37), .B(new_n313_), .C1(new_n318_), .C2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NOR3_X1   g122(.A1(new_n315_), .A2(new_n316_), .A3(KEYINPUT75), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n320_), .B(new_n319_), .C1(new_n324_), .C2(new_n314_), .ZN(new_n325_));
  AOI21_X1  g124(.A(KEYINPUT37), .B1(new_n325_), .B2(new_n313_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G231gat), .A2(G233gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT77), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n219_), .B(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G57gat), .B(G64gat), .ZN(new_n330_));
  AND2_X1   g129(.A1(new_n330_), .A2(KEYINPUT11), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n330_), .A2(KEYINPUT11), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G71gat), .B(G78gat), .ZN(new_n333_));
  OR3_X1    g132(.A1(new_n331_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n330_), .A2(new_n333_), .A3(KEYINPUT11), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n329_), .B(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT80), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G183gat), .B(G211gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  XOR2_X1   g141(.A(G127gat), .B(G155gat), .Z(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  OR2_X1    g143(.A1(new_n344_), .A2(KEYINPUT17), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(KEYINPUT17), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n339_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT81), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n346_), .B(KEYINPUT79), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n350_), .A2(new_n337_), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  NOR3_X1   g151(.A1(new_n323_), .A2(new_n326_), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(G183gat), .ZN(new_n354_));
  INV_X1    g153(.A(G190gat), .ZN(new_n355_));
  NOR3_X1   g154(.A1(new_n354_), .A2(new_n355_), .A3(KEYINPUT23), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT23), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n358_), .B1(G183gat), .B2(G190gat), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n359_), .A2(KEYINPUT87), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n359_), .A2(KEYINPUT87), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n357_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n362_), .B1(G183gat), .B2(G190gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G169gat), .A2(G176gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT22), .B(G169gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT97), .ZN(new_n366_));
  INV_X1    g165(.A(G176gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n363_), .A2(new_n364_), .A3(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(G169gat), .A2(G176gat), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT86), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n372_), .A2(KEYINPUT24), .A3(new_n364_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n370_), .B(KEYINPUT86), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT24), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT25), .B(G183gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT26), .B(G190gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n356_), .A2(new_n359_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n373_), .A2(new_n376_), .A3(new_n379_), .A4(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n369_), .A2(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(G211gat), .B(G218gat), .Z(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(G204gat), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n386_), .A2(G197gat), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n386_), .A2(G197gat), .ZN(new_n388_));
  OAI21_X1  g187(.A(KEYINPUT21), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(KEYINPUT92), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT92), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n391_), .B1(G197gat), .B2(new_n386_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n390_), .B1(new_n392_), .B2(new_n388_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n385_), .B(new_n389_), .C1(new_n393_), .C2(KEYINPUT21), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n393_), .A2(KEYINPUT21), .A3(new_n384_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n383_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n396_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n362_), .A2(new_n379_), .A3(new_n373_), .A4(new_n376_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n365_), .A2(new_n367_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(G183gat), .A2(G190gat), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n364_), .B(new_n400_), .C1(new_n380_), .C2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n398_), .A2(new_n399_), .A3(new_n402_), .ZN(new_n403_));
  AND3_X1   g202(.A1(new_n397_), .A2(KEYINPUT20), .A3(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G226gat), .A2(G233gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT19), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n404_), .A2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT20), .B1(new_n383_), .B2(new_n396_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n398_), .B1(new_n399_), .B2(new_n402_), .ZN(new_n410_));
  NOR3_X1   g209(.A1(new_n409_), .A2(new_n406_), .A3(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n408_), .A2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G64gat), .B(G92gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  XOR2_X1   g214(.A(G8gat), .B(G36gat), .Z(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n412_), .B(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G225gat), .A2(G233gat), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT91), .ZN(new_n421_));
  INV_X1    g220(.A(G148gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n421_), .B1(new_n242_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT2), .ZN(new_n424_));
  OR3_X1    g223(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT2), .ZN(new_n426_));
  OAI211_X1 g225(.A(new_n421_), .B(new_n426_), .C1(new_n242_), .C2(new_n422_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n424_), .A2(new_n425_), .A3(new_n427_), .A4(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(KEYINPUT90), .B1(G155gat), .B2(G162gat), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(KEYINPUT90), .A2(G155gat), .A3(G162gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n429_), .B(new_n433_), .C1(G155gat), .C2(G162gat), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT1), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n431_), .A2(new_n435_), .A3(new_n432_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n432_), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT1), .B1(new_n437_), .B2(new_n430_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n436_), .B(new_n438_), .C1(G155gat), .C2(G162gat), .ZN(new_n439_));
  XOR2_X1   g238(.A(G141gat), .B(G148gat), .Z(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n434_), .A2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G127gat), .B(G134gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G113gat), .B(G120gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n442_), .A2(new_n446_), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n447_), .A2(KEYINPUT4), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n434_), .A2(new_n441_), .A3(new_n445_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n445_), .B1(new_n434_), .B2(new_n441_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(KEYINPUT99), .B1(new_n451_), .B2(KEYINPUT4), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n434_), .A2(new_n441_), .A3(new_n445_), .ZN(new_n453_));
  AND4_X1   g252(.A1(KEYINPUT99), .A2(new_n447_), .A3(KEYINPUT4), .A4(new_n453_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n420_), .B(new_n448_), .C1(new_n452_), .C2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT100), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  XOR2_X1   g256(.A(G1gat), .B(G29gat), .Z(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(G85gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(KEYINPUT0), .B(G57gat), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n459_), .B(new_n460_), .Z(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n451_), .A2(new_n419_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n451_), .A2(KEYINPUT99), .A3(KEYINPUT4), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n447_), .A2(KEYINPUT4), .A3(new_n453_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT99), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n464_), .A2(new_n467_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n468_), .A2(KEYINPUT100), .A3(new_n420_), .A4(new_n448_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n457_), .A2(new_n462_), .A3(new_n463_), .A4(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT33), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n468_), .A2(new_n419_), .A3(new_n448_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n451_), .A2(new_n420_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(new_n461_), .A3(new_n474_), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n470_), .A2(new_n475_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n418_), .B(new_n472_), .C1(new_n476_), .C2(new_n471_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n457_), .A2(new_n463_), .A3(new_n469_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n461_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(new_n470_), .ZN(new_n480_));
  AND4_X1   g279(.A1(KEYINPUT20), .A2(new_n397_), .A3(new_n407_), .A4(new_n403_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT101), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n410_), .B1(new_n409_), .B2(new_n482_), .ZN(new_n483_));
  OAI211_X1 g282(.A(KEYINPUT101), .B(KEYINPUT20), .C1(new_n383_), .C2(new_n396_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n481_), .B1(new_n485_), .B2(new_n406_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n417_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT32), .ZN(new_n488_));
  OR2_X1    g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n412_), .A2(new_n488_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n480_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n477_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT30), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n399_), .A2(new_n493_), .A3(new_n402_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n493_), .B1(new_n399_), .B2(new_n402_), .ZN(new_n496_));
  NOR3_X1   g295(.A1(new_n495_), .A2(KEYINPUT89), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT89), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n399_), .A2(new_n402_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT30), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n499_), .B1(new_n501_), .B2(new_n494_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G71gat), .B(G99gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT88), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G15gat), .B(G43gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G227gat), .A2(G233gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT31), .B1(new_n502_), .B2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT89), .B1(new_n495_), .B2(new_n496_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n507_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n506_), .B(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT31), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n510_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n509_), .A2(new_n446_), .A3(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n446_), .B1(new_n509_), .B2(new_n514_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n498_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n509_), .A2(new_n514_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(new_n445_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n509_), .A2(new_n514_), .A3(new_n446_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n519_), .A2(new_n497_), .A3(new_n520_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n517_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n442_), .A2(KEYINPUT29), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G228gat), .A2(G233gat), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n524_), .A2(new_n396_), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT29), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n527_), .B1(new_n434_), .B2(new_n441_), .ZN(new_n528_));
  OAI211_X1 g327(.A(G228gat), .B(G233gat), .C1(new_n528_), .C2(new_n398_), .ZN(new_n529_));
  XOR2_X1   g328(.A(G78gat), .B(G106gat), .Z(new_n530_));
  NAND3_X1  g329(.A1(new_n526_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n531_), .A2(KEYINPUT93), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n526_), .A2(new_n529_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n530_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT94), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n531_), .A2(KEYINPUT93), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n533_), .A2(KEYINPUT94), .A3(new_n534_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n532_), .A2(new_n537_), .A3(new_n538_), .A4(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(G50gat), .B1(new_n442_), .B2(KEYINPUT29), .ZN(new_n541_));
  INV_X1    g340(.A(G50gat), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n434_), .A2(new_n441_), .A3(new_n527_), .A4(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT28), .B(G22gat), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n541_), .A2(new_n545_), .A3(new_n543_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n540_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT96), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT95), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n552_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n553_));
  AOI211_X1 g352(.A(KEYINPUT95), .B(new_n530_), .C1(new_n526_), .C2(new_n529_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n531_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n551_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n535_), .A2(KEYINPUT95), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n533_), .A2(new_n552_), .A3(new_n534_), .ZN(new_n559_));
  AND4_X1   g358(.A1(new_n551_), .A2(new_n556_), .A3(new_n558_), .A4(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n550_), .B1(new_n557_), .B2(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n523_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n492_), .A2(new_n562_), .ZN(new_n563_));
  OR3_X1    g362(.A1(new_n409_), .A2(new_n406_), .A3(new_n410_), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n564_), .B(new_n487_), .C1(new_n407_), .C2(new_n404_), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n565_), .B(KEYINPUT27), .C1(new_n486_), .C2(new_n487_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT27), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n412_), .B(new_n487_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n567_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n480_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n522_), .A2(new_n561_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n522_), .A2(new_n561_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n570_), .B(new_n571_), .C1(new_n572_), .C2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n563_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n336_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n290_), .A2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n277_), .A2(new_n289_), .A3(new_n336_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n577_), .A2(KEYINPUT70), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G230gat), .A2(G233gat), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n580_), .B(KEYINPUT64), .Z(new_n581_));
  OR2_X1    g380(.A1(new_n578_), .A2(KEYINPUT70), .ZN(new_n582_));
  AND3_X1   g381(.A1(new_n579_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n577_), .A2(KEYINPUT12), .A3(new_n578_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT12), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n290_), .A2(new_n585_), .A3(new_n576_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n581_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n583_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(KEYINPUT71), .B(G204gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(KEYINPUT5), .B(G176gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G120gat), .B(G148gat), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n591_), .B(new_n592_), .Z(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n588_), .B(new_n594_), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n595_), .A2(KEYINPUT13), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(KEYINPUT13), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  AND4_X1   g398(.A1(new_n251_), .A2(new_n353_), .A3(new_n575_), .A4(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n600_), .A2(new_n214_), .A3(new_n480_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT38), .ZN(new_n602_));
  INV_X1    g401(.A(new_n251_), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n598_), .A2(new_n352_), .A3(new_n603_), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n604_), .A2(KEYINPUT102), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n313_), .B1(new_n318_), .B2(new_n321_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n607_), .B1(new_n604_), .B2(KEYINPUT102), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n605_), .A2(new_n608_), .A3(new_n575_), .ZN(new_n609_));
  OAI21_X1  g408(.A(G1gat), .B1(new_n609_), .B2(new_n571_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n602_), .A2(new_n610_), .ZN(G1324gat));
  INV_X1    g410(.A(new_n570_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n600_), .A2(new_n215_), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT39), .ZN(new_n614_));
  INV_X1    g413(.A(new_n609_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n612_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n614_), .B1(new_n616_), .B2(G8gat), .ZN(new_n617_));
  AOI211_X1 g416(.A(KEYINPUT39), .B(new_n215_), .C1(new_n615_), .C2(new_n612_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n613_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n619_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g419(.A(G15gat), .B1(new_n609_), .B2(new_n522_), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n621_), .B(KEYINPUT41), .Z(new_n622_));
  INV_X1    g421(.A(G15gat), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n600_), .A2(new_n623_), .A3(new_n523_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(G1326gat));
  INV_X1    g424(.A(new_n561_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G22gat), .B1(new_n609_), .B2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT42), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n626_), .A2(G22gat), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT103), .Z(new_n630_));
  NAND2_X1  g429(.A1(new_n600_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n628_), .A2(new_n631_), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n632_), .B(KEYINPUT104), .Z(G1327gat));
  AOI21_X1  g432(.A(new_n606_), .B1(new_n563_), .B2(new_n574_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n349_), .A2(new_n351_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n598_), .A2(new_n635_), .A3(new_n603_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  OR3_X1    g436(.A1(new_n637_), .A2(G29gat), .A3(new_n571_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT105), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n639_), .B1(new_n323_), .B2(new_n326_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT37), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n606_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n642_), .A2(KEYINPUT105), .A3(new_n322_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n575_), .A2(new_n640_), .A3(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT43), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT43), .B1(new_n563_), .B2(new_n574_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n323_), .A2(new_n326_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n645_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT106), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n651_), .A2(KEYINPUT44), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n650_), .A2(new_n653_), .A3(new_n636_), .ZN(new_n654_));
  AOI22_X1  g453(.A1(new_n644_), .A2(KEYINPUT43), .B1(new_n648_), .B2(new_n646_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n636_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n652_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n654_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G29gat), .B1(new_n659_), .B2(new_n571_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n660_), .A2(KEYINPUT107), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n660_), .A2(KEYINPUT107), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n638_), .B1(new_n661_), .B2(new_n662_), .ZN(G1328gat));
  NOR3_X1   g462(.A1(new_n637_), .A2(G36gat), .A3(new_n570_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n654_), .A2(new_n657_), .A3(new_n612_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT108), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n667_), .A2(new_n668_), .A3(G36gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n667_), .B2(G36gat), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n666_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT46), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  OAI211_X1 g472(.A(KEYINPUT46), .B(new_n666_), .C1(new_n669_), .C2(new_n670_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1329gat));
  INV_X1    g474(.A(KEYINPUT110), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n654_), .A2(new_n657_), .A3(new_n523_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G43gat), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n637_), .A2(G43gat), .A3(new_n522_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n676_), .B1(new_n678_), .B2(new_n680_), .ZN(new_n681_));
  AOI211_X1 g480(.A(KEYINPUT110), .B(new_n679_), .C1(new_n677_), .C2(G43gat), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT47), .ZN(new_n683_));
  OR3_X1    g482(.A1(new_n681_), .A2(new_n682_), .A3(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n683_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1330gat));
  OAI21_X1  g485(.A(G50gat), .B1(new_n659_), .B2(new_n626_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n561_), .A2(new_n542_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n687_), .B1(new_n637_), .B2(new_n688_), .ZN(G1331gat));
  NAND2_X1  g488(.A1(new_n598_), .A2(new_n603_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n690_), .B1(new_n563_), .B2(new_n574_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n691_), .A2(new_n635_), .A3(new_n606_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT111), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n694_), .A2(G57gat), .A3(new_n480_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT112), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(G57gat), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n691_), .A2(new_n353_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n698_), .B1(new_n699_), .B2(new_n571_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n694_), .A2(KEYINPUT112), .A3(G57gat), .A4(new_n480_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n697_), .A2(new_n700_), .A3(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT113), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n697_), .A2(KEYINPUT113), .A3(new_n700_), .A4(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1332gat));
  OAI21_X1  g505(.A(G64gat), .B1(new_n693_), .B2(new_n570_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT48), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n570_), .A2(G64gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n708_), .B1(new_n699_), .B2(new_n709_), .ZN(G1333gat));
  OAI21_X1  g509(.A(G71gat), .B1(new_n693_), .B2(new_n522_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT49), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n522_), .A2(G71gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n712_), .B1(new_n699_), .B2(new_n713_), .ZN(G1334gat));
  OR3_X1    g513(.A1(new_n699_), .A2(G78gat), .A3(new_n626_), .ZN(new_n715_));
  OAI21_X1  g514(.A(G78gat), .B1(new_n693_), .B2(new_n626_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n716_), .A2(KEYINPUT50), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(KEYINPUT50), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n715_), .B1(new_n717_), .B2(new_n718_), .ZN(G1335gat));
  NAND4_X1  g518(.A1(new_n634_), .A2(new_n603_), .A3(new_n598_), .A4(new_n352_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT114), .ZN(new_n721_));
  AOI21_X1  g520(.A(G85gat), .B1(new_n721_), .B2(new_n480_), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n655_), .A2(new_n635_), .A3(new_n690_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n480_), .A2(new_n278_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n722_), .B1(new_n723_), .B2(new_n724_), .ZN(G1336gat));
  AOI21_X1  g524(.A(G92gat), .B1(new_n721_), .B2(new_n612_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT115), .Z(new_n727_));
  AND2_X1   g526(.A1(new_n612_), .A2(G92gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n723_), .B2(new_n728_), .ZN(G1337gat));
  AOI21_X1  g528(.A(new_n253_), .B1(new_n723_), .B2(new_n523_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n523_), .A2(new_n287_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n721_), .B2(new_n731_), .ZN(new_n732_));
  XOR2_X1   g531(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n733_));
  XNOR2_X1  g532(.A(new_n732_), .B(new_n733_), .ZN(G1338gat));
  AOI21_X1  g533(.A(new_n254_), .B1(new_n723_), .B2(new_n561_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT52), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n735_), .B(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n721_), .A2(new_n254_), .A3(new_n561_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n737_), .A2(new_n738_), .A3(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1339gat));
  INV_X1    g541(.A(KEYINPUT54), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n353_), .A2(new_n743_), .A3(new_n603_), .A4(new_n599_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n642_), .A2(new_n603_), .A3(new_n635_), .A4(new_n322_), .ZN(new_n745_));
  OAI21_X1  g544(.A(KEYINPUT54), .B1(new_n745_), .B2(new_n598_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n588_), .A2(new_n593_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n234_), .A2(new_n223_), .A3(new_n235_), .A4(new_n236_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n221_), .A2(new_n222_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n749_), .A2(new_n249_), .A3(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n246_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n250_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n752_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT119), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n584_), .A2(new_n581_), .A3(new_n586_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT118), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n584_), .A2(KEYINPUT118), .A3(new_n581_), .A4(new_n586_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n581_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n578_), .A2(KEYINPUT12), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n336_), .B1(new_n277_), .B2(new_n289_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n586_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n762_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n587_), .A2(KEYINPUT55), .ZN(new_n770_));
  AND4_X1   g569(.A1(new_n756_), .A2(new_n761_), .A3(new_n769_), .A4(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n584_), .A2(new_n586_), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT55), .B1(new_n772_), .B2(new_n762_), .ZN(new_n773_));
  AOI211_X1 g572(.A(new_n768_), .B(new_n581_), .C1(new_n584_), .C2(new_n586_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n756_), .B1(new_n775_), .B2(new_n761_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n771_), .A2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT56), .B1(new_n777_), .B2(new_n594_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n759_), .A2(new_n760_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n769_), .A2(new_n770_), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT119), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n775_), .A2(new_n756_), .A3(new_n761_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n781_), .A2(KEYINPUT56), .A3(new_n594_), .A4(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n748_), .B(new_n755_), .C1(new_n778_), .C2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT58), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n781_), .A2(new_n594_), .A3(new_n782_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT56), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n783_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n791_), .A2(KEYINPUT58), .A3(new_n748_), .A4(new_n755_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n787_), .A2(new_n648_), .A3(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n251_), .A2(new_n748_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n794_), .B1(new_n790_), .B2(new_n783_), .ZN(new_n795_));
  AOI211_X1 g594(.A(new_n752_), .B(new_n595_), .C1(new_n753_), .C2(new_n754_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n606_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT57), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  OAI211_X1 g598(.A(KEYINPUT57), .B(new_n606_), .C1(new_n795_), .C2(new_n796_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n793_), .A2(new_n799_), .A3(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n747_), .B1(new_n801_), .B2(new_n352_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n573_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n612_), .A2(new_n571_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n802_), .A2(new_n803_), .A3(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(G113gat), .B1(new_n806_), .B2(new_n251_), .ZN(new_n807_));
  OR2_X1    g606(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  XOR2_X1   g609(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NOR4_X1   g611(.A1(new_n802_), .A2(new_n803_), .A3(new_n805_), .A4(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n603_), .B1(new_n810_), .B2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n807_), .B1(new_n815_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g615(.A(KEYINPUT60), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n599_), .B2(G120gat), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n806_), .A2(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n598_), .B(new_n819_), .C1(new_n809_), .C2(new_n813_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(G120gat), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n806_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(G1341gat));
  AOI21_X1  g622(.A(G127gat), .B1(new_n806_), .B2(new_n635_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n352_), .B1(new_n810_), .B2(new_n814_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n824_), .B1(new_n825_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g625(.A(G134gat), .B1(new_n806_), .B2(new_n607_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n647_), .B1(new_n810_), .B2(new_n814_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n827_), .B1(new_n828_), .B2(G134gat), .ZN(G1343gat));
  NOR3_X1   g628(.A1(new_n802_), .A2(new_n626_), .A3(new_n523_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n804_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n831_), .A2(new_n603_), .ZN(new_n832_));
  XOR2_X1   g631(.A(KEYINPUT121), .B(G141gat), .Z(new_n833_));
  XNOR2_X1  g632(.A(new_n832_), .B(new_n833_), .ZN(G1344gat));
  NOR2_X1   g633(.A1(new_n831_), .A2(new_n599_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(new_n422_), .ZN(G1345gat));
  NOR2_X1   g635(.A1(new_n831_), .A2(new_n352_), .ZN(new_n837_));
  XOR2_X1   g636(.A(KEYINPUT61), .B(G155gat), .Z(new_n838_));
  XNOR2_X1  g637(.A(new_n837_), .B(new_n838_), .ZN(G1346gat));
  AND3_X1   g638(.A1(new_n640_), .A2(G162gat), .A3(new_n643_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n830_), .A2(new_n804_), .A3(new_n840_), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n787_), .A2(new_n648_), .A3(new_n792_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n799_), .A2(new_n800_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n352_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n747_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  AND4_X1   g645(.A1(new_n607_), .A2(new_n846_), .A3(new_n572_), .A4(new_n804_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n841_), .B1(new_n847_), .B2(G162gat), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT122), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n841_), .B(KEYINPUT122), .C1(new_n847_), .C2(G162gat), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1347gat));
  NOR2_X1   g651(.A1(new_n802_), .A2(new_n803_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n570_), .A2(new_n480_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n853_), .A2(new_n251_), .A3(new_n366_), .A4(new_n854_), .ZN(new_n855_));
  AND3_X1   g654(.A1(new_n853_), .A2(new_n251_), .A3(new_n854_), .ZN(new_n856_));
  INV_X1    g655(.A(G169gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n855_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(KEYINPUT62), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT62), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n861_), .ZN(G1348gat));
  NAND2_X1  g661(.A1(new_n853_), .A2(new_n854_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(new_n599_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(new_n367_), .ZN(G1349gat));
  NOR2_X1   g664(.A1(new_n863_), .A2(new_n352_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n377_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n867_), .B1(new_n354_), .B2(new_n866_), .ZN(G1350gat));
  AND3_X1   g667(.A1(new_n853_), .A2(new_n648_), .A3(new_n854_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n607_), .A2(new_n378_), .ZN(new_n870_));
  OAI22_X1  g669(.A1(new_n869_), .A2(new_n355_), .B1(new_n863_), .B2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(KEYINPUT123), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT123), .ZN(new_n873_));
  OAI221_X1 g672(.A(new_n873_), .B1(new_n863_), .B2(new_n870_), .C1(new_n869_), .C2(new_n355_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n872_), .A2(new_n874_), .ZN(G1351gat));
  NAND2_X1  g674(.A1(new_n854_), .A2(new_n572_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n876_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n251_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(KEYINPUT124), .B(G197gat), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(G1352gat));
  NAND2_X1  g679(.A1(new_n877_), .A2(new_n598_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g681(.A1(new_n877_), .A2(new_n635_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n884_));
  AND2_X1   g683(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n883_), .A2(new_n884_), .A3(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n886_), .B1(new_n883_), .B2(new_n884_), .ZN(G1354gat));
  INV_X1    g686(.A(KEYINPUT125), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n888_), .B1(new_n877_), .B2(new_n607_), .ZN(new_n889_));
  NOR4_X1   g688(.A1(new_n802_), .A2(KEYINPUT125), .A3(new_n606_), .A4(new_n876_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n889_), .A2(new_n890_), .A3(G218gat), .ZN(new_n891_));
  INV_X1    g690(.A(new_n876_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n846_), .A2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(G218gat), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n647_), .A2(new_n894_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(KEYINPUT126), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n893_), .A2(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(KEYINPUT127), .B1(new_n891_), .B2(new_n897_), .ZN(new_n898_));
  OAI21_X1  g697(.A(KEYINPUT125), .B1(new_n893_), .B2(new_n606_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n877_), .A2(new_n888_), .A3(new_n607_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n899_), .A2(new_n894_), .A3(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT127), .ZN(new_n902_));
  INV_X1    g701(.A(new_n897_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n901_), .A2(new_n902_), .A3(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n898_), .A2(new_n904_), .ZN(G1355gat));
endmodule


