//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 1 0 1 1 1 1 1 0 1 0 0 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n589_, new_n590_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n596_, new_n597_, new_n598_, new_n599_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n791_, new_n792_, new_n794_, new_n795_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n812_,
    new_n813_, new_n814_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n826_,
    new_n827_, new_n828_, new_n830_, new_n831_, new_n833_, new_n834_,
    new_n835_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT15), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G85gat), .B(G92gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT9), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT10), .B(G99gat), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n209_), .A2(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT6), .ZN(new_n212_));
  INV_X1    g011(.A(G85gat), .ZN(new_n213_));
  INV_X1    g012(.A(G92gat), .ZN(new_n214_));
  OR3_X1    g013(.A1(new_n213_), .A2(new_n214_), .A3(KEYINPUT9), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n208_), .A2(new_n210_), .A3(new_n212_), .A4(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT8), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT6), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n211_), .B(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT65), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n212_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT7), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT64), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G99gat), .A2(G106gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n220_), .A2(new_n222_), .A3(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n217_), .B1(new_n227_), .B2(new_n207_), .ZN(new_n228_));
  AOI211_X1 g027(.A(KEYINPUT8), .B(new_n206_), .C1(new_n226_), .C2(new_n212_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n216_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  MUX2_X1   g029(.A(new_n204_), .B(new_n205_), .S(new_n230_), .Z(new_n231_));
  NAND2_X1  g030(.A1(G232gat), .A2(G233gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT34), .ZN(new_n233_));
  XOR2_X1   g032(.A(new_n233_), .B(KEYINPUT35), .Z(new_n234_));
  NAND2_X1  g033(.A1(new_n231_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT69), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n231_), .A2(KEYINPUT69), .A3(new_n234_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n233_), .A2(KEYINPUT35), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n237_), .B(new_n238_), .C1(new_n239_), .C2(new_n231_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G190gat), .B(G218gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(G162gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT67), .B(G134gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT36), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT68), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n240_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT70), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n244_), .B(KEYINPUT36), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n240_), .A2(new_n251_), .ZN(new_n252_));
  OR3_X1    g051(.A1(new_n240_), .A2(new_n249_), .A3(new_n247_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n250_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT37), .ZN(new_n255_));
  AND2_X1   g054(.A1(new_n240_), .A2(KEYINPUT71), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n251_), .B1(new_n240_), .B2(KEYINPUT71), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n248_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n258_), .A2(KEYINPUT37), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n255_), .A2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G1gat), .B(G8gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT72), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G15gat), .B(G22gat), .ZN(new_n263_));
  INV_X1    g062(.A(G1gat), .ZN(new_n264_));
  INV_X1    g063(.A(G8gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT14), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n263_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n262_), .B(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G231gat), .A2(G233gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT73), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n268_), .B(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G57gat), .B(G64gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT11), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(KEYINPUT11), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G71gat), .B(G78gat), .ZN(new_n275_));
  MUX2_X1   g074(.A(new_n273_), .B(new_n274_), .S(new_n275_), .Z(new_n276_));
  XOR2_X1   g075(.A(new_n271_), .B(new_n276_), .Z(new_n277_));
  XOR2_X1   g076(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n278_));
  XNOR2_X1  g077(.A(G127gat), .B(G155gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G183gat), .B(G211gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT17), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n282_), .A2(new_n283_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n277_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n286_), .B1(new_n284_), .B2(new_n277_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n260_), .A2(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(new_n288_), .B(KEYINPUT75), .Z(new_n289_));
  INV_X1    g088(.A(KEYINPUT81), .ZN(new_n290_));
  INV_X1    g089(.A(G183gat), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n291_), .A2(KEYINPUT23), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G183gat), .A2(G190gat), .ZN(new_n293_));
  AOI22_X1  g092(.A1(new_n292_), .A2(G190gat), .B1(KEYINPUT23), .B2(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(G183gat), .A2(G190gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n290_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT22), .B(G169gat), .ZN(new_n299_));
  INV_X1    g098(.A(G176gat), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n298_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n293_), .A2(KEYINPUT23), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT23), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n303_), .A2(G183gat), .A3(G190gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n305_), .B(KEYINPUT81), .C1(G183gat), .C2(G190gat), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n296_), .A2(new_n301_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(G169gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(new_n300_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n309_), .A2(KEYINPUT24), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(KEYINPUT24), .A3(new_n297_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n310_), .B1(new_n311_), .B2(KEYINPUT79), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT25), .B(G183gat), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT78), .ZN(new_n314_));
  INV_X1    g113(.A(G190gat), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT26), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n315_), .A2(KEYINPUT26), .ZN(new_n317_));
  OAI211_X1 g116(.A(new_n313_), .B(new_n316_), .C1(new_n317_), .C2(new_n314_), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n293_), .A2(KEYINPUT80), .A3(KEYINPUT23), .ZN(new_n319_));
  AOI21_X1  g118(.A(KEYINPUT80), .B1(new_n293_), .B2(KEYINPUT23), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n304_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n297_), .A2(KEYINPUT24), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT79), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n322_), .A2(new_n323_), .A3(new_n309_), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n312_), .A2(new_n318_), .A3(new_n321_), .A4(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n307_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT30), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G227gat), .A2(G233gat), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n329_), .B(KEYINPUT82), .Z(new_n330_));
  XNOR2_X1  g129(.A(new_n328_), .B(new_n330_), .ZN(new_n331_));
  XOR2_X1   g130(.A(G15gat), .B(G43gat), .Z(new_n332_));
  XNOR2_X1  g131(.A(G71gat), .B(G99gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n331_), .A2(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n331_), .A2(new_n334_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT83), .ZN(new_n337_));
  OR3_X1    g136(.A1(new_n335_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n337_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G127gat), .B(G134gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G113gat), .B(G120gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT31), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n338_), .A2(new_n339_), .A3(new_n344_), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n339_), .A2(new_n344_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  XOR2_X1   g146(.A(G64gat), .B(G92gat), .Z(new_n348_));
  XNOR2_X1  g147(.A(G8gat), .B(G36gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n351_));
  XOR2_X1   g150(.A(new_n350_), .B(new_n351_), .Z(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G226gat), .A2(G233gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT95), .B1(new_n294_), .B2(new_n310_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT26), .B(G190gat), .ZN(new_n359_));
  AOI22_X1  g158(.A1(new_n313_), .A2(new_n359_), .B1(new_n322_), .B2(new_n309_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT95), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n305_), .B(new_n361_), .C1(KEYINPUT24), .C2(new_n309_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n358_), .A2(new_n360_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n304_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT80), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n302_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n293_), .A2(KEYINPUT80), .A3(KEYINPUT23), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n364_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n301_), .B1(new_n368_), .B2(new_n295_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n363_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT96), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G211gat), .B(G218gat), .ZN(new_n372_));
  AND2_X1   g171(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n373_));
  NOR2_X1   g172(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n374_));
  OAI21_X1  g173(.A(G197gat), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(G197gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(G204gat), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n372_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT21), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT21), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n375_), .A2(new_n380_), .A3(new_n377_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n372_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT88), .ZN(new_n383_));
  INV_X1    g182(.A(G204gat), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n383_), .B1(G197gat), .B2(new_n384_), .ZN(new_n385_));
  NOR3_X1   g184(.A1(new_n376_), .A2(KEYINPUT88), .A3(G204gat), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n374_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(new_n376_), .A3(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n380_), .B1(new_n387_), .B2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n379_), .B1(new_n382_), .B2(new_n391_), .ZN(new_n392_));
  AND3_X1   g191(.A1(new_n370_), .A2(new_n371_), .A3(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n371_), .B1(new_n370_), .B2(new_n392_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT20), .B1(new_n326_), .B2(new_n392_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n357_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n370_), .A2(new_n392_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n326_), .A2(new_n392_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n399_), .A2(KEYINPUT20), .A3(new_n357_), .A4(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n353_), .B1(new_n398_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT98), .ZN(new_n404_));
  NOR3_X1   g203(.A1(new_n393_), .A2(new_n396_), .A3(new_n394_), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n352_), .B(new_n401_), .C1(new_n405_), .C2(new_n357_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n403_), .A2(new_n404_), .A3(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n394_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n370_), .A2(new_n371_), .A3(new_n392_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n397_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(new_n356_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(new_n401_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n412_), .A2(KEYINPUT98), .A3(new_n353_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n407_), .A2(new_n413_), .ZN(new_n414_));
  OR2_X1    g213(.A1(new_n414_), .A2(KEYINPUT27), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n400_), .A2(KEYINPUT20), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n357_), .B1(new_n416_), .B2(new_n399_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT102), .ZN(new_n418_));
  OAI22_X1  g217(.A1(new_n417_), .A2(new_n418_), .B1(new_n356_), .B2(new_n410_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n405_), .A2(KEYINPUT102), .A3(new_n357_), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  OAI211_X1 g220(.A(KEYINPUT27), .B(new_n406_), .C1(new_n421_), .C2(new_n352_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n415_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT3), .ZN(new_n424_));
  INV_X1    g223(.A(G141gat), .ZN(new_n425_));
  INV_X1    g224(.A(G148gat), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G141gat), .A2(G148gat), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT2), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n427_), .A2(new_n430_), .A3(new_n431_), .A4(new_n432_), .ZN(new_n433_));
  OR2_X1    g232(.A1(G155gat), .A2(G162gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G155gat), .A2(G162gat), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n434_), .A2(KEYINPUT85), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(KEYINPUT85), .B1(new_n434_), .B2(new_n435_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n433_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n435_), .A2(KEYINPUT1), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT1), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n440_), .A2(G155gat), .A3(G162gat), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n439_), .A2(new_n441_), .A3(new_n434_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n425_), .A2(new_n426_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(new_n428_), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n438_), .A2(new_n444_), .ZN(new_n445_));
  XOR2_X1   g244(.A(new_n340_), .B(new_n341_), .Z(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n342_), .A2(new_n438_), .A3(new_n444_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(KEYINPUT4), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G225gat), .A2(G233gat), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT4), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n445_), .A2(new_n446_), .A3(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n449_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n447_), .A2(new_n450_), .A3(new_n448_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(KEYINPUT99), .B(KEYINPUT0), .Z(new_n457_));
  XNOR2_X1  g256(.A(G1gat), .B(G29gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G57gat), .B(G85gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n456_), .A2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n454_), .A2(new_n455_), .A3(new_n461_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n445_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT29), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n392_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(G228gat), .A3(G233gat), .ZN(new_n469_));
  OR2_X1    g268(.A1(new_n469_), .A2(KEYINPUT90), .ZN(new_n470_));
  OR3_X1    g269(.A1(new_n466_), .A2(KEYINPUT87), .A3(new_n467_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G228gat), .A2(G233gat), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT87), .B1(new_n466_), .B2(new_n467_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n471_), .A2(new_n472_), .A3(new_n473_), .A4(new_n392_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n469_), .A2(KEYINPUT90), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n470_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G78gat), .B(G106gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT91), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT92), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n476_), .B(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n445_), .A2(KEYINPUT29), .ZN(new_n482_));
  XOR2_X1   g281(.A(G22gat), .B(G50gat), .Z(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n485_));
  XOR2_X1   g284(.A(new_n484_), .B(new_n485_), .Z(new_n486_));
  NAND2_X1  g285(.A1(new_n481_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n476_), .A2(new_n478_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT93), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n476_), .A2(new_n480_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n486_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT93), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n476_), .A2(new_n492_), .A3(new_n478_), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n489_), .A2(new_n490_), .A3(new_n491_), .A4(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n487_), .A2(new_n494_), .ZN(new_n495_));
  NOR4_X1   g294(.A1(new_n347_), .A2(new_n423_), .A3(new_n465_), .A4(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT103), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n464_), .A2(KEYINPUT33), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT33), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n454_), .A2(new_n499_), .A3(new_n455_), .A4(new_n461_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n447_), .A2(new_n451_), .A3(new_n448_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n462_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT100), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n449_), .A2(new_n450_), .A3(new_n453_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT100), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n462_), .A2(new_n506_), .A3(new_n502_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n504_), .A2(new_n505_), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n501_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT101), .B1(new_n414_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT101), .ZN(new_n512_));
  AOI211_X1 g311(.A(new_n512_), .B(new_n509_), .C1(new_n407_), .C2(new_n413_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n412_), .B1(KEYINPUT32), .B2(new_n352_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n352_), .A2(KEYINPUT32), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n515_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n465_), .ZN(new_n517_));
  NOR3_X1   g316(.A1(new_n514_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n511_), .A2(new_n513_), .A3(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n497_), .B1(new_n519_), .B2(new_n495_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n423_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n521_), .A2(new_n517_), .A3(new_n495_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n406_), .A2(new_n404_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n352_), .B1(new_n411_), .B2(new_n401_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  AOI211_X1 g324(.A(new_n404_), .B(new_n352_), .C1(new_n411_), .C2(new_n401_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n510_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n512_), .ZN(new_n528_));
  OR3_X1    g327(.A1(new_n514_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n414_), .A2(KEYINPUT101), .A3(new_n510_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n487_), .A2(new_n494_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(KEYINPUT103), .A3(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n520_), .A2(new_n522_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT84), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n347_), .B(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n496_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n230_), .A2(new_n276_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n230_), .A2(new_n276_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n538_), .A2(KEYINPUT12), .A3(new_n539_), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n539_), .A2(KEYINPUT12), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G230gat), .A2(G233gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n538_), .A2(new_n539_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n544_), .B1(new_n543_), .B2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT5), .B(G176gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(G204gat), .ZN(new_n548_));
  XOR2_X1   g347(.A(G120gat), .B(G148gat), .Z(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n546_), .B(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT66), .B(KEYINPUT13), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT66), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n551_), .B1(new_n554_), .B2(KEYINPUT13), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  MUX2_X1   g355(.A(new_n204_), .B(new_n205_), .S(new_n268_), .Z(new_n557_));
  NAND2_X1  g356(.A1(G229gat), .A2(G233gat), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n268_), .B(new_n204_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n558_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n559_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT76), .B(G113gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(G141gat), .ZN(new_n565_));
  XOR2_X1   g364(.A(G169gat), .B(G197gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n563_), .B(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n568_), .B(KEYINPUT77), .Z(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n556_), .A2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n537_), .A2(new_n571_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n289_), .A2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n573_), .A2(new_n264_), .A3(new_n465_), .ZN(new_n574_));
  XOR2_X1   g373(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n575_));
  XOR2_X1   g374(.A(new_n574_), .B(new_n575_), .Z(new_n576_));
  XOR2_X1   g375(.A(new_n258_), .B(KEYINPUT105), .Z(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n287_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n572_), .A2(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n264_), .B1(new_n581_), .B2(new_n465_), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n576_), .A2(new_n582_), .ZN(G1324gat));
  AOI21_X1  g382(.A(new_n265_), .B1(new_n581_), .B2(new_n423_), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n584_), .B(KEYINPUT39), .Z(new_n585_));
  NAND3_X1  g384(.A1(new_n573_), .A2(new_n265_), .A3(new_n423_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n587_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g387(.A(G15gat), .ZN(new_n589_));
  INV_X1    g388(.A(new_n536_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n573_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n591_), .B(KEYINPUT106), .Z(new_n592_));
  AOI21_X1  g391(.A(new_n589_), .B1(new_n581_), .B2(new_n590_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT41), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(G1326gat));
  INV_X1    g394(.A(G22gat), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n596_), .B1(new_n581_), .B2(new_n495_), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n597_), .B(KEYINPUT42), .Z(new_n598_));
  NAND3_X1  g397(.A1(new_n573_), .A2(new_n596_), .A3(new_n495_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(G1327gat));
  NOR2_X1   g399(.A1(new_n577_), .A2(new_n287_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NOR3_X1   g401(.A1(new_n602_), .A2(new_n571_), .A3(new_n537_), .ZN(new_n603_));
  AOI21_X1  g402(.A(G29gat), .B1(new_n603_), .B2(new_n465_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n556_), .A2(new_n570_), .A3(new_n579_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT43), .ZN(new_n607_));
  INV_X1    g406(.A(new_n496_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n531_), .A2(KEYINPUT103), .A3(new_n532_), .ZN(new_n609_));
  AOI21_X1  g408(.A(KEYINPUT103), .B1(new_n531_), .B2(new_n532_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n423_), .A2(new_n532_), .A3(new_n465_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n609_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n608_), .B1(new_n612_), .B2(new_n590_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n260_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n607_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n537_), .A2(KEYINPUT43), .A3(new_n260_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n606_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(KEYINPUT107), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT44), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n613_), .A2(new_n607_), .A3(new_n614_), .ZN(new_n620_));
  OAI21_X1  g419(.A(KEYINPUT43), .B1(new_n537_), .B2(new_n260_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n605_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT107), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n618_), .A2(new_n619_), .A3(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n622_), .A2(KEYINPUT44), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n627_), .A2(new_n465_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n604_), .B1(new_n628_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g428(.A(KEYINPUT46), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT108), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n521_), .B1(new_n622_), .B2(KEYINPUT44), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n625_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n631_), .B1(new_n625_), .B2(new_n632_), .ZN(new_n634_));
  INV_X1    g433(.A(G36gat), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n633_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n603_), .A2(new_n635_), .A3(new_n423_), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n637_), .B(KEYINPUT45), .Z(new_n638_));
  OAI21_X1  g437(.A(new_n630_), .B1(new_n636_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n634_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n625_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(G36gat), .A3(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n638_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n642_), .A2(KEYINPUT46), .A3(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n639_), .A2(new_n644_), .ZN(G1329gat));
  INV_X1    g444(.A(new_n347_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n627_), .A2(G43gat), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(G43gat), .ZN(new_n648_));
  INV_X1    g447(.A(new_n603_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n648_), .B1(new_n649_), .B2(new_n536_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n647_), .A2(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n647_), .A2(new_n650_), .A3(new_n652_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1330gat));
  AOI21_X1  g455(.A(G50gat), .B1(new_n603_), .B2(new_n495_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n627_), .A2(new_n495_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n658_), .B2(G50gat), .ZN(G1331gat));
  NOR2_X1   g458(.A1(new_n537_), .A2(new_n570_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT110), .ZN(new_n661_));
  INV_X1    g460(.A(new_n556_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n663_), .A2(new_n289_), .ZN(new_n664_));
  AOI21_X1  g463(.A(G57gat), .B1(new_n664_), .B2(new_n465_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n580_), .A2(new_n569_), .A3(new_n662_), .A4(new_n613_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n666_), .A2(new_n517_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n665_), .B1(G57gat), .B2(new_n667_), .ZN(G1332gat));
  INV_X1    g467(.A(G64gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n664_), .A2(new_n669_), .A3(new_n423_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G64gat), .B1(new_n666_), .B2(new_n521_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT48), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(G1333gat));
  INV_X1    g472(.A(G71gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n664_), .A2(new_n674_), .A3(new_n590_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G71gat), .B1(new_n666_), .B2(new_n536_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT49), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(G1334gat));
  INV_X1    g477(.A(G78gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n664_), .A2(new_n679_), .A3(new_n495_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G78gat), .B1(new_n666_), .B2(new_n532_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT50), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(G1335gat));
  AND3_X1   g482(.A1(new_n661_), .A2(new_n662_), .A3(new_n601_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n213_), .B1(new_n685_), .B2(new_n517_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n620_), .A2(new_n621_), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n687_), .A2(KEYINPUT111), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n556_), .A2(new_n570_), .A3(new_n287_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(KEYINPUT111), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n688_), .A2(new_n689_), .A3(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n691_), .A2(G85gat), .A3(new_n465_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n686_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(G1336gat));
  OAI21_X1  g493(.A(new_n214_), .B1(new_n685_), .B2(new_n521_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n691_), .A2(G92gat), .A3(new_n423_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(G1337gat));
  NAND4_X1  g497(.A1(new_n688_), .A2(new_n590_), .A3(new_n689_), .A4(new_n690_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n347_), .A2(new_n209_), .ZN(new_n700_));
  AOI22_X1  g499(.A1(new_n699_), .A2(G99gat), .B1(new_n684_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT51), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(KEYINPUT112), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT112), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n704_), .A2(KEYINPUT51), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n703_), .B(new_n705_), .ZN(G1338gat));
  OR3_X1    g505(.A1(new_n685_), .A2(G106gat), .A3(new_n532_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n687_), .A2(new_n495_), .A3(new_n689_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(KEYINPUT113), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT113), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n687_), .A2(new_n710_), .A3(new_n495_), .A4(new_n689_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n709_), .A2(G106gat), .A3(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT52), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT52), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n709_), .A2(new_n714_), .A3(G106gat), .A4(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n707_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT53), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT53), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n707_), .A2(new_n719_), .A3(new_n716_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1339gat));
  INV_X1    g520(.A(KEYINPUT120), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n546_), .A2(new_n550_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT55), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n544_), .A2(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n542_), .A2(KEYINPUT55), .A3(new_n543_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n725_), .B(new_n726_), .C1(new_n543_), .C2(new_n542_), .ZN(new_n727_));
  AOI21_X1  g526(.A(KEYINPUT56), .B1(new_n727_), .B2(new_n550_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n723_), .B1(new_n728_), .B2(KEYINPUT116), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n550_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT56), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n727_), .A2(KEYINPUT56), .A3(new_n550_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n570_), .B(new_n729_), .C1(new_n734_), .C2(KEYINPUT116), .ZN(new_n735_));
  INV_X1    g534(.A(new_n563_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n560_), .A2(new_n558_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n567_), .B1(new_n557_), .B2(new_n561_), .ZN(new_n738_));
  AOI22_X1  g537(.A1(new_n736_), .A2(new_n567_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n551_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n735_), .A2(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n741_), .A2(new_n577_), .A3(KEYINPUT57), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT117), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n741_), .A2(new_n577_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT57), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n734_), .B(new_n739_), .C1(new_n546_), .C2(new_n550_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT58), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n749_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(new_n614_), .A3(new_n751_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n741_), .A2(new_n577_), .A3(KEYINPUT117), .A4(KEYINPUT57), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n744_), .A2(new_n747_), .A3(new_n752_), .A4(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(new_n579_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n569_), .A2(new_n287_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n756_), .A2(KEYINPUT114), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n662_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(KEYINPUT114), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n758_), .A2(new_n260_), .A3(new_n759_), .ZN(new_n760_));
  XOR2_X1   g559(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n758_), .A2(new_n260_), .A3(new_n759_), .A4(new_n761_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n755_), .A2(new_n766_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n646_), .A2(new_n521_), .A3(new_n465_), .A4(new_n532_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT118), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT119), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n770_), .A2(KEYINPUT59), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n770_), .A2(KEYINPUT59), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n767_), .B(new_n769_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n765_), .B1(new_n754_), .B2(new_n579_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n769_), .ZN(new_n775_));
  OAI22_X1  g574(.A1(new_n774_), .A2(new_n775_), .B1(new_n770_), .B2(KEYINPUT59), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n773_), .A2(new_n776_), .A3(new_n570_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(G113gat), .ZN(new_n778_));
  NOR4_X1   g577(.A1(new_n774_), .A2(G113gat), .A3(new_n569_), .A4(new_n775_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n722_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n781_));
  AOI211_X1 g580(.A(KEYINPUT120), .B(new_n779_), .C1(new_n777_), .C2(G113gat), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n781_), .A2(new_n782_), .ZN(G1340gat));
  NOR2_X1   g582(.A1(new_n774_), .A2(new_n775_), .ZN(new_n784_));
  INV_X1    g583(.A(G120gat), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n785_), .B1(new_n556_), .B2(KEYINPUT60), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n784_), .B(new_n786_), .C1(KEYINPUT60), .C2(new_n785_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT121), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n773_), .A2(new_n662_), .A3(new_n776_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n788_), .B1(new_n785_), .B2(new_n789_), .ZN(G1341gat));
  AOI21_X1  g589(.A(G127gat), .B1(new_n784_), .B2(new_n287_), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n773_), .A2(new_n287_), .A3(new_n776_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g592(.A(G134gat), .B1(new_n784_), .B2(new_n578_), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n773_), .A2(G134gat), .A3(new_n776_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(new_n795_), .B2(new_n614_), .ZN(G1343gat));
  NOR3_X1   g595(.A1(new_n774_), .A2(new_n517_), .A3(new_n590_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n423_), .A2(new_n532_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n799_), .A2(new_n569_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(new_n425_), .ZN(G1344gat));
  NOR2_X1   g600(.A1(new_n799_), .A2(new_n556_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(new_n426_), .ZN(G1345gat));
  NOR2_X1   g602(.A1(new_n590_), .A2(new_n517_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n767_), .A2(new_n798_), .A3(new_n287_), .A4(new_n804_), .ZN(new_n805_));
  OR2_X1    g604(.A1(new_n805_), .A2(G155gat), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(G155gat), .ZN(new_n807_));
  XNOR2_X1  g606(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n806_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n808_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n809_), .A2(new_n810_), .ZN(G1346gat));
  INV_X1    g610(.A(G162gat), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n799_), .A2(new_n812_), .A3(new_n260_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n797_), .A2(new_n798_), .A3(new_n578_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n813_), .B1(new_n812_), .B2(new_n814_), .ZN(G1347gat));
  NOR2_X1   g614(.A1(new_n774_), .A2(new_n495_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n590_), .A2(new_n517_), .A3(new_n423_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(KEYINPUT123), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(G169gat), .B1(new_n819_), .B2(new_n569_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT62), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n816_), .A2(new_n570_), .A3(new_n299_), .A4(new_n818_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n820_), .A2(new_n821_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n822_), .A2(new_n823_), .A3(new_n824_), .ZN(G1348gat));
  OAI22_X1  g624(.A1(new_n819_), .A2(new_n556_), .B1(KEYINPUT124), .B2(new_n300_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n300_), .A2(KEYINPUT124), .ZN(new_n827_));
  XOR2_X1   g626(.A(new_n827_), .B(KEYINPUT125), .Z(new_n828_));
  XOR2_X1   g627(.A(new_n826_), .B(new_n828_), .Z(G1349gat));
  NOR2_X1   g628(.A1(new_n819_), .A2(new_n579_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n313_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(new_n830_), .B2(new_n291_), .ZN(G1350gat));
  OAI21_X1  g631(.A(G190gat), .B1(new_n819_), .B2(new_n260_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n578_), .A2(new_n359_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(KEYINPUT126), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n833_), .B1(new_n819_), .B2(new_n835_), .ZN(G1351gat));
  NOR3_X1   g635(.A1(new_n521_), .A2(new_n465_), .A3(new_n532_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n767_), .A2(new_n536_), .A3(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n838_), .A2(new_n569_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(new_n376_), .ZN(G1352gat));
  INV_X1    g639(.A(new_n838_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n662_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(G204gat), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n373_), .A2(new_n374_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(new_n842_), .ZN(G1353gat));
  NOR2_X1   g644(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT127), .ZN(new_n848_));
  NAND2_X1  g647(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n849_));
  AND4_X1   g648(.A1(new_n848_), .A2(new_n841_), .A3(new_n287_), .A4(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n838_), .A2(new_n579_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n848_), .B1(new_n851_), .B2(new_n849_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n847_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n841_), .A2(new_n287_), .A3(new_n849_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(KEYINPUT127), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n851_), .A2(new_n848_), .A3(new_n849_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(new_n846_), .A3(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n853_), .A2(new_n857_), .ZN(G1354gat));
  AND3_X1   g657(.A1(new_n841_), .A2(G218gat), .A3(new_n614_), .ZN(new_n859_));
  AOI21_X1  g658(.A(G218gat), .B1(new_n841_), .B2(new_n578_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n859_), .A2(new_n860_), .ZN(G1355gat));
endmodule


