//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 0 1 0 0 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 0 0 1 1 0 0 1 0 1 0 1 1 1 1 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n801_, new_n802_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n924_,
    new_n925_, new_n927_, new_n928_, new_n930_, new_n931_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n947_, new_n948_, new_n949_, new_n951_, new_n952_, new_n954_,
    new_n955_, new_n957_, new_n958_, new_n959_, new_n960_, new_n962_,
    new_n963_, new_n965_, new_n966_, new_n967_, new_n968_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XOR2_X1   g002(.A(KEYINPUT10), .B(G99gat), .Z(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  XOR2_X1   g005(.A(G85gat), .B(G92gat), .Z(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT9), .ZN(new_n208_));
  INV_X1    g007(.A(G85gat), .ZN(new_n209_));
  INV_X1    g008(.A(G92gat), .ZN(new_n210_));
  OR3_X1    g009(.A1(new_n209_), .A2(new_n210_), .A3(KEYINPUT9), .ZN(new_n211_));
  AND3_X1   g010(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n212_));
  AOI21_X1  g011(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n206_), .A2(new_n208_), .A3(new_n211_), .A4(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n217_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT6), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(KEYINPUT66), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n218_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n225_));
  INV_X1    g024(.A(G99gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n226_), .A3(new_n205_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT7), .ZN(new_n230_));
  NOR2_X1   g029(.A1(G99gat), .A2(G106gat), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n230_), .B1(new_n231_), .B2(KEYINPUT64), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n229_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n227_), .A2(new_n228_), .A3(new_n230_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n224_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n207_), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT8), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n214_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n238_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT8), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n207_), .A2(new_n240_), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n216_), .B1(new_n237_), .B2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G57gat), .B(G64gat), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n244_), .A2(KEYINPUT11), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(KEYINPUT11), .ZN(new_n246_));
  XOR2_X1   g045(.A(G71gat), .B(G78gat), .Z(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n246_), .A2(new_n247_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n243_), .A2(KEYINPUT67), .A3(new_n250_), .ZN(new_n251_));
  NOR3_X1   g050(.A1(new_n212_), .A2(new_n213_), .A3(new_n217_), .ZN(new_n252_));
  AOI21_X1  g051(.A(KEYINPUT66), .B1(new_n221_), .B2(new_n222_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n226_), .A2(new_n205_), .ZN(new_n255_));
  OAI21_X1  g054(.A(KEYINPUT7), .B1(new_n255_), .B2(new_n228_), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT64), .B1(new_n231_), .B2(new_n225_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n234_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n254_), .A2(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n240_), .B1(new_n259_), .B2(new_n207_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n239_), .A2(new_n241_), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n215_), .B(new_n250_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT67), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n251_), .A2(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n243_), .A2(new_n250_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n203_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n203_), .B1(new_n243_), .B2(new_n250_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT12), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n236_), .B1(new_n254_), .B2(new_n258_), .ZN(new_n270_));
  OAI22_X1  g069(.A1(new_n270_), .A2(new_n240_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n215_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n250_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n269_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  AOI211_X1 g073(.A(KEYINPUT12), .B(new_n250_), .C1(new_n271_), .C2(new_n215_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n268_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G120gat), .B(G148gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT5), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G176gat), .B(G204gat), .ZN(new_n279_));
  XOR2_X1   g078(.A(new_n278_), .B(new_n279_), .Z(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n267_), .A2(new_n276_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n281_), .B1(new_n267_), .B2(new_n276_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n285_), .A2(KEYINPUT13), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(KEYINPUT13), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT68), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G232gat), .A2(G233gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT34), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n292_), .A2(KEYINPUT35), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G29gat), .B(G36gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G43gat), .B(G50gat), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n295_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT15), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n293_), .B1(new_n272_), .B2(new_n299_), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n243_), .A2(KEYINPUT70), .A3(new_n298_), .ZN(new_n301_));
  AOI21_X1  g100(.A(KEYINPUT70), .B1(new_n243_), .B2(new_n298_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n300_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n292_), .A2(KEYINPUT35), .ZN(new_n304_));
  XOR2_X1   g103(.A(new_n304_), .B(KEYINPUT69), .Z(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n303_), .A2(new_n306_), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n300_), .B(new_n305_), .C1(new_n301_), .C2(new_n302_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n307_), .A2(KEYINPUT72), .A3(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G190gat), .B(G218gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT71), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G134gat), .B(G162gat), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n311_), .B(new_n312_), .Z(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n309_), .A2(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n315_), .A2(KEYINPUT36), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT37), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n307_), .A2(new_n308_), .A3(new_n313_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT36), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n315_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n317_), .A2(new_n318_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n318_), .B1(new_n317_), .B2(new_n322_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G231gat), .A2(G233gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n250_), .B(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G1gat), .A2(G8gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT14), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT73), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT73), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n329_), .A2(new_n332_), .A3(KEYINPUT14), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G15gat), .B(G22gat), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n331_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT74), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n331_), .A2(new_n337_), .A3(new_n334_), .A4(new_n333_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(G1gat), .B(G8gat), .Z(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n336_), .A2(new_n340_), .A3(new_n338_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n328_), .B(new_n344_), .Z(new_n345_));
  INV_X1    g144(.A(KEYINPUT17), .ZN(new_n346_));
  XOR2_X1   g145(.A(G127gat), .B(G155gat), .Z(new_n347_));
  XNOR2_X1  g146(.A(G183gat), .B(G211gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  NOR3_X1   g150(.A1(new_n345_), .A2(new_n346_), .A3(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(KEYINPUT17), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n345_), .A2(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n326_), .A2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n290_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G169gat), .A2(G176gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT81), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n359_), .B(KEYINPUT24), .C1(G169gat), .C2(G176gat), .ZN(new_n360_));
  NOR3_X1   g159(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G183gat), .A2(G190gat), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT23), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT82), .B(KEYINPUT23), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n366_), .B1(new_n367_), .B2(new_n364_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n360_), .A2(new_n362_), .A3(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT26), .B(G190gat), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT79), .ZN(new_n372_));
  INV_X1    g171(.A(G183gat), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT25), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  OR2_X1    g173(.A1(new_n373_), .A2(KEYINPUT25), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n371_), .B(new_n374_), .C1(new_n375_), .C2(new_n372_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT80), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n370_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n363_), .A2(new_n365_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n379_), .B1(new_n367_), .B2(new_n363_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  OR2_X1    g180(.A1(G183gat), .A2(G190gat), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT83), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT83), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n381_), .A2(new_n385_), .A3(new_n382_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT22), .B(G169gat), .ZN(new_n387_));
  INV_X1    g186(.A(G176gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  AND2_X1   g188(.A1(new_n389_), .A2(new_n359_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n384_), .A2(new_n386_), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n378_), .A2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(KEYINPUT30), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G71gat), .B(G99gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT31), .ZN(new_n396_));
  OR2_X1    g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n396_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  XOR2_X1   g198(.A(KEYINPUT85), .B(G15gat), .Z(new_n400_));
  NAND2_X1  g199(.A1(G227gat), .A2(G233gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT84), .B(G43gat), .ZN(new_n403_));
  XOR2_X1   g202(.A(new_n402_), .B(new_n403_), .Z(new_n404_));
  XNOR2_X1  g203(.A(G127gat), .B(G134gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G113gat), .B(G120gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n407_), .A2(KEYINPUT86), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT86), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n405_), .A2(new_n406_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n408_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n404_), .B(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n399_), .A2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n397_), .A2(new_n398_), .A3(new_n412_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT102), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G8gat), .B(G36gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT18), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G64gat), .B(G92gat), .ZN(new_n420_));
  XOR2_X1   g219(.A(new_n419_), .B(new_n420_), .Z(new_n421_));
  XNOR2_X1  g220(.A(G197gat), .B(G204gat), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT21), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n423_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G211gat), .B(G218gat), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  OR3_X1    g226(.A1(new_n422_), .A2(new_n426_), .A3(new_n423_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT92), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT96), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n390_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n368_), .A2(new_n382_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n389_), .A2(new_n359_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT96), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n432_), .A2(new_n433_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT92), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n427_), .A2(new_n437_), .A3(new_n428_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n430_), .A2(new_n436_), .A3(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(KEYINPUT94), .B1(new_n358_), .B2(KEYINPUT24), .ZN(new_n440_));
  INV_X1    g239(.A(G169gat), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n440_), .B1(new_n441_), .B2(new_n388_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n358_), .A2(KEYINPUT94), .A3(KEYINPUT24), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT25), .B(G183gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n371_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT95), .B1(new_n380_), .B2(new_n361_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT95), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n381_), .A2(new_n449_), .A3(new_n362_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n447_), .B1(new_n448_), .B2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT20), .B1(new_n439_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT100), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT100), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n454_), .B(KEYINPUT20), .C1(new_n439_), .C2(new_n451_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n392_), .A2(new_n429_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n453_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G226gat), .A2(G233gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT19), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n451_), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n435_), .A2(new_n433_), .ZN(new_n462_));
  AOI21_X1  g261(.A(KEYINPUT97), .B1(new_n462_), .B2(new_n432_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT97), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n436_), .A2(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n461_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n429_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n459_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT20), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n434_), .B1(new_n383_), .B2(KEYINPUT83), .ZN(new_n470_));
  AOI22_X1  g269(.A1(new_n470_), .A2(new_n386_), .B1(new_n370_), .B2(new_n377_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n429_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n469_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n467_), .A2(new_n468_), .A3(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n421_), .B1(new_n460_), .B2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n462_), .A2(KEYINPUT97), .A3(new_n432_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n436_), .A2(new_n464_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n472_), .B1(new_n478_), .B2(new_n461_), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT20), .B1(new_n392_), .B2(new_n429_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n459_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n478_), .A2(new_n472_), .A3(new_n461_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n468_), .A2(KEYINPUT20), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n483_), .B1(new_n392_), .B2(new_n429_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n482_), .A2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n481_), .A2(new_n421_), .A3(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT27), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n475_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT101), .ZN(new_n490_));
  INV_X1    g289(.A(new_n421_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n468_), .B1(new_n467_), .B2(new_n473_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n485_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n491_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(new_n486_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT27), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n490_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  AOI211_X1 g296(.A(KEYINPUT101), .B(KEYINPUT27), .C1(new_n494_), .C2(new_n486_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n489_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G155gat), .A2(G162gat), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n500_), .A2(KEYINPUT1), .ZN(new_n501_));
  NOR2_X1   g300(.A1(G155gat), .A2(G162gat), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n503_), .B1(KEYINPUT1), .B2(new_n500_), .ZN(new_n504_));
  AND2_X1   g303(.A1(G141gat), .A2(G148gat), .ZN(new_n505_));
  NOR2_X1   g304(.A1(G141gat), .A2(G148gat), .ZN(new_n506_));
  NOR3_X1   g305(.A1(new_n504_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n500_), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n509_), .A2(new_n502_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT90), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n506_), .B(KEYINPUT3), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n505_), .A2(KEYINPUT2), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT88), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT87), .B(KEYINPUT2), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n515_), .B1(new_n516_), .B2(new_n505_), .ZN(new_n517_));
  OR3_X1    g316(.A1(new_n516_), .A2(new_n515_), .A3(new_n505_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n514_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT89), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n511_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  AOI211_X1 g320(.A(KEYINPUT89), .B(new_n514_), .C1(new_n518_), .C2(new_n517_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n508_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT28), .B1(new_n523_), .B2(KEYINPUT29), .ZN(new_n524_));
  INV_X1    g323(.A(new_n519_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT89), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n519_), .A2(new_n520_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n526_), .A2(new_n527_), .A3(new_n511_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT28), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT29), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .A4(new_n508_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G22gat), .B(G50gat), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n524_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n532_), .B1(new_n524_), .B2(new_n531_), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT93), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n524_), .A2(new_n531_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n532_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT93), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n539_), .A2(new_n540_), .A3(new_n533_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G78gat), .B(G106gat), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n430_), .A2(new_n438_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n544_), .B1(new_n523_), .B2(KEYINPUT29), .ZN(new_n545_));
  INV_X1    g344(.A(G233gat), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT91), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n547_), .A2(G228gat), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(G228gat), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n546_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n545_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n523_), .A2(KEYINPUT29), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n554_), .A2(new_n429_), .A3(new_n552_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n543_), .B1(new_n553_), .B2(new_n555_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n555_), .B(new_n543_), .C1(new_n545_), .C2(new_n552_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n536_), .B(new_n541_), .C1(new_n556_), .C2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n556_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n540_), .B1(new_n539_), .B2(new_n533_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n560_), .A2(new_n561_), .A3(new_n557_), .ZN(new_n562_));
  AOI21_X1  g361(.A(KEYINPUT4), .B1(new_n523_), .B2(new_n411_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n528_), .A2(new_n407_), .A3(new_n508_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n523_), .A2(new_n411_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n563_), .B1(new_n566_), .B2(KEYINPUT4), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G225gat), .A2(G233gat), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(G1gat), .B(G29gat), .Z(new_n571_));
  XNOR2_X1  g370(.A(G57gat), .B(G85gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT98), .B(KEYINPUT0), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n573_), .B(new_n574_), .Z(new_n575_));
  AOI21_X1  g374(.A(new_n569_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n570_), .A2(new_n575_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n575_), .ZN(new_n579_));
  AOI211_X1 g378(.A(new_n568_), .B(new_n563_), .C1(new_n566_), .C2(KEYINPUT4), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n579_), .B1(new_n580_), .B2(new_n576_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n559_), .A2(new_n562_), .A3(new_n578_), .A4(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n417_), .B1(new_n499_), .B2(new_n582_), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n481_), .A2(new_n421_), .A3(new_n485_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n421_), .B1(new_n481_), .B2(new_n485_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n496_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT101), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n495_), .A2(new_n490_), .A3(new_n496_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n488_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n559_), .A2(new_n562_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n581_), .A2(new_n578_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n589_), .A2(KEYINPUT102), .A3(new_n590_), .A4(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n583_), .A2(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n575_), .B1(new_n570_), .B2(new_n577_), .ZN(new_n595_));
  OAI21_X1  g394(.A(KEYINPUT99), .B1(new_n595_), .B2(KEYINPUT33), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT99), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT33), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n581_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n567_), .A2(new_n569_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n575_), .B1(new_n566_), .B2(new_n568_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n602_), .A2(new_n495_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n595_), .A2(KEYINPUT33), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n596_), .A2(new_n599_), .A3(new_n603_), .A4(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n421_), .A2(KEYINPUT32), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n481_), .A2(new_n606_), .A3(new_n485_), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n460_), .A2(new_n474_), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n591_), .B(new_n607_), .C1(new_n608_), .C2(new_n606_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n590_), .B1(new_n605_), .B2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n416_), .B1(new_n594_), .B2(new_n610_), .ZN(new_n611_));
  NOR4_X1   g410(.A1(new_n416_), .A2(new_n499_), .A3(new_n590_), .A4(new_n591_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G229gat), .A2(G233gat), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n296_), .A2(KEYINPUT76), .A3(new_n297_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT76), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n298_), .A2(new_n618_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n342_), .A2(new_n617_), .A3(new_n619_), .A4(new_n343_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  AOI22_X1  g420(.A1(new_n342_), .A2(new_n343_), .B1(new_n617_), .B2(new_n619_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n616_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n622_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n299_), .A2(new_n343_), .A3(new_n342_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n624_), .A2(new_n625_), .A3(new_n615_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G113gat), .B(G141gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT77), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G169gat), .B(G197gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n623_), .A2(new_n626_), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT78), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n623_), .A2(new_n626_), .A3(KEYINPUT78), .A4(new_n631_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n623_), .A2(new_n626_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(new_n630_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(KEYINPUT103), .B1(new_n614_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT103), .ZN(new_n641_));
  INV_X1    g440(.A(new_n639_), .ZN(new_n642_));
  AOI211_X1 g441(.A(new_n641_), .B(new_n642_), .C1(new_n611_), .C2(new_n613_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n357_), .B1(new_n640_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT104), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  OAI211_X1 g445(.A(KEYINPUT104), .B(new_n357_), .C1(new_n640_), .C2(new_n643_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n592_), .A2(G1gat), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n646_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT38), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n605_), .A2(new_n609_), .ZN(new_n652_));
  OAI211_X1 g451(.A(new_n583_), .B(new_n593_), .C1(new_n652_), .C2(new_n590_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n612_), .B1(new_n653_), .B2(new_n416_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n317_), .A2(new_n322_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n288_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(new_n639_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n355_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n656_), .A2(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G1gat), .B1(new_n661_), .B2(new_n592_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n649_), .A2(new_n650_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n651_), .A2(new_n662_), .A3(new_n663_), .ZN(G1324gat));
  NOR2_X1   g463(.A1(new_n589_), .A2(G8gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n646_), .A2(new_n647_), .A3(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(KEYINPUT106), .A2(KEYINPUT39), .ZN(new_n667_));
  INV_X1    g466(.A(new_n655_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n614_), .A2(new_n499_), .A3(new_n668_), .A4(new_n660_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(KEYINPUT105), .A3(G8gat), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(KEYINPUT105), .B1(new_n669_), .B2(G8gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n667_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n672_), .ZN(new_n674_));
  XOR2_X1   g473(.A(KEYINPUT106), .B(KEYINPUT39), .Z(new_n675_));
  NAND3_X1  g474(.A1(new_n674_), .A2(new_n670_), .A3(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n666_), .A2(new_n673_), .A3(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n666_), .A2(new_n673_), .A3(new_n676_), .A4(new_n678_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1325gat));
  OAI21_X1  g481(.A(G15gat), .B1(new_n661_), .B2(new_n416_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT41), .Z(new_n684_));
  NOR2_X1   g483(.A1(new_n416_), .A2(G15gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n646_), .A2(new_n647_), .A3(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(G1326gat));
  NAND3_X1  g486(.A1(new_n656_), .A2(new_n590_), .A3(new_n660_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(G22gat), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(KEYINPUT108), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT108), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n688_), .A2(new_n691_), .A3(G22gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n690_), .A2(KEYINPUT42), .A3(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n590_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n694_), .A2(G22gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n646_), .A2(new_n647_), .A3(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n693_), .A2(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT42), .B1(new_n690_), .B2(new_n692_), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n697_), .A2(new_n698_), .ZN(G1327gat));
  NOR2_X1   g498(.A1(new_n668_), .A2(new_n355_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(new_n657_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n641_), .B1(new_n654_), .B2(new_n642_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n614_), .A2(KEYINPUT103), .A3(new_n639_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n701_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(G29gat), .B1(new_n704_), .B2(new_n591_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n658_), .A2(new_n355_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n325_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(new_n323_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT109), .ZN(new_n710_));
  OAI21_X1  g509(.A(KEYINPUT43), .B1(new_n654_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n614_), .A2(new_n712_), .A3(new_n709_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n707_), .B1(new_n711_), .B2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT44), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n715_), .A2(G29gat), .A3(new_n591_), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n714_), .A2(KEYINPUT44), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n705_), .B1(new_n716_), .B2(new_n717_), .ZN(G1328gat));
  NOR2_X1   g517(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n719_));
  INV_X1    g518(.A(G36gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n589_), .B1(new_n714_), .B2(KEYINPUT44), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n717_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT45), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n589_), .A2(G36gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n704_), .A2(new_n723_), .A3(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n723_), .B1(new_n704_), .B2(new_n724_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n719_), .B1(new_n722_), .B2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n715_), .A2(new_n499_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n714_), .A2(KEYINPUT44), .ZN(new_n731_));
  OAI21_X1  g530(.A(G36gat), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n727_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(new_n725_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n719_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n732_), .A2(new_n734_), .A3(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n729_), .A2(new_n736_), .ZN(G1329gat));
  INV_X1    g536(.A(G43gat), .ZN(new_n738_));
  INV_X1    g537(.A(new_n704_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(new_n416_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n416_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n715_), .A2(G43gat), .A3(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n740_), .B1(new_n742_), .B2(new_n731_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT47), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT47), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n740_), .B(new_n745_), .C1(new_n742_), .C2(new_n731_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(G1330gat));
  NAND2_X1  g546(.A1(new_n715_), .A2(new_n590_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G50gat), .B1(new_n748_), .B2(new_n731_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n694_), .A2(G50gat), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT111), .Z(new_n751_));
  OAI21_X1  g550(.A(new_n749_), .B1(new_n739_), .B2(new_n751_), .ZN(G1331gat));
  INV_X1    g551(.A(KEYINPUT112), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n753_), .B1(new_n654_), .B2(new_n639_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n614_), .A2(KEYINPUT112), .A3(new_n642_), .ZN(new_n755_));
  AOI211_X1 g554(.A(new_n657_), .B(new_n356_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(G57gat), .B1(new_n756_), .B2(new_n591_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n642_), .A2(new_n355_), .ZN(new_n758_));
  NOR4_X1   g557(.A1(new_n654_), .A2(new_n289_), .A3(new_n655_), .A4(new_n758_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n592_), .A2(KEYINPUT113), .ZN(new_n760_));
  MUX2_X1   g559(.A(KEYINPUT113), .B(new_n760_), .S(G57gat), .Z(new_n761_));
  AOI21_X1  g560(.A(new_n757_), .B1(new_n759_), .B2(new_n761_), .ZN(G1332gat));
  INV_X1    g561(.A(G64gat), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n763_), .B1(new_n759_), .B2(new_n499_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT48), .Z(new_n765_));
  NAND3_X1  g564(.A1(new_n756_), .A2(new_n763_), .A3(new_n499_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(G1333gat));
  INV_X1    g566(.A(G71gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n768_), .B1(new_n759_), .B2(new_n741_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT49), .Z(new_n770_));
  NAND2_X1  g569(.A1(new_n741_), .A2(new_n768_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT114), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n756_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n770_), .A2(new_n773_), .ZN(G1334gat));
  INV_X1    g573(.A(G78gat), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n756_), .A2(new_n775_), .A3(new_n590_), .ZN(new_n776_));
  AOI211_X1 g575(.A(KEYINPUT50), .B(new_n775_), .C1(new_n759_), .C2(new_n590_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT50), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n759_), .A2(new_n590_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n779_), .B2(G78gat), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n776_), .B1(new_n777_), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT115), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n776_), .B(new_n783_), .C1(new_n780_), .C2(new_n777_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(G1335gat));
  NOR2_X1   g584(.A1(new_n355_), .A2(new_n639_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n288_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT116), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n326_), .B(KEYINPUT109), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n712_), .B1(new_n614_), .B2(new_n789_), .ZN(new_n790_));
  AOI211_X1 g589(.A(KEYINPUT43), .B(new_n326_), .C1(new_n611_), .C2(new_n613_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n788_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n711_), .A2(KEYINPUT116), .A3(new_n713_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n787_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(G85gat), .B1(new_n795_), .B2(new_n592_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n290_), .A2(new_n700_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n797_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(new_n209_), .A3(new_n591_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n796_), .A2(new_n799_), .ZN(G1336gat));
  OAI21_X1  g599(.A(G92gat), .B1(new_n795_), .B2(new_n589_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n798_), .A2(new_n210_), .A3(new_n499_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(G1337gat));
  AOI21_X1  g602(.A(new_n226_), .B1(new_n794_), .B2(new_n741_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n741_), .A2(new_n204_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n798_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n798_), .A2(new_n806_), .A3(new_n807_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n805_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n810_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n814_), .A2(new_n808_), .ZN(new_n815_));
  OAI21_X1  g614(.A(KEYINPUT51), .B1(new_n815_), .B2(new_n804_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n813_), .A2(new_n816_), .ZN(G1338gat));
  NAND3_X1  g616(.A1(new_n798_), .A2(new_n205_), .A3(new_n590_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n711_), .A2(new_n713_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n787_), .A2(new_n694_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n819_), .B1(new_n822_), .B2(G106gat), .ZN(new_n823_));
  AOI211_X1 g622(.A(KEYINPUT52), .B(new_n205_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n818_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT53), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n827_), .B(new_n818_), .C1(new_n823_), .C2(new_n824_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(G1339gat));
  NAND2_X1  g628(.A1(new_n589_), .A2(new_n591_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n830_), .A2(new_n416_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n264_), .B(new_n251_), .C1(new_n274_), .C2(new_n275_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n276_), .A2(KEYINPUT55), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT12), .B1(new_n243_), .B2(new_n250_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n272_), .A2(new_n269_), .A3(new_n273_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT55), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(new_n838_), .A3(new_n268_), .ZN(new_n839_));
  AOI221_X4 g638(.A(KEYINPUT118), .B1(new_n833_), .B2(new_n203_), .C1(new_n834_), .C2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n834_), .A2(new_n839_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n833_), .A2(new_n203_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n841_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n280_), .B1(new_n840_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT56), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n838_), .B1(new_n837_), .B2(new_n268_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n262_), .A2(new_n202_), .ZN(new_n849_));
  AOI211_X1 g648(.A(KEYINPUT55), .B(new_n849_), .C1(new_n835_), .C2(new_n836_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n843_), .B1(new_n848_), .B2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(KEYINPUT118), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n842_), .A2(new_n841_), .A3(new_n843_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n854_), .A2(KEYINPUT56), .A3(new_n280_), .ZN(new_n855_));
  AND3_X1   g654(.A1(new_n847_), .A2(KEYINPUT121), .A3(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n615_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n858_), .A2(KEYINPUT119), .A3(new_n630_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n624_), .A2(new_n625_), .A3(new_n616_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n858_), .A2(new_n630_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n861_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  AOI22_X1  g663(.A1(new_n859_), .A2(new_n864_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n857_), .B1(new_n865_), .B2(new_n282_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n862_), .A2(new_n863_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n868_));
  AND4_X1   g667(.A1(new_n857_), .A2(new_n636_), .A3(new_n868_), .A4(new_n282_), .ZN(new_n869_));
  OAI22_X1  g668(.A1(new_n847_), .A2(KEYINPUT121), .B1(new_n866_), .B2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n832_), .B1(new_n856_), .B2(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n871_), .A2(KEYINPUT122), .A3(new_n709_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n866_), .A2(new_n869_), .ZN(new_n874_));
  AOI21_X1  g673(.A(KEYINPUT56), .B1(new_n854_), .B2(new_n280_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT121), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n874_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n847_), .A2(KEYINPUT121), .A3(new_n855_), .ZN(new_n878_));
  AOI21_X1  g677(.A(KEYINPUT58), .B1(new_n877_), .B2(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n873_), .B1(new_n879_), .B2(new_n326_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n877_), .A2(KEYINPUT58), .A3(new_n878_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n872_), .A2(new_n880_), .A3(new_n881_), .ZN(new_n882_));
  AOI211_X1 g681(.A(new_n846_), .B(new_n281_), .C1(new_n852_), .C2(new_n853_), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n639_), .B(new_n282_), .C1(new_n875_), .C2(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n865_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(KEYINPUT57), .B1(new_n886_), .B2(new_n668_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT57), .ZN(new_n888_));
  AOI211_X1 g687(.A(new_n888_), .B(new_n655_), .C1(new_n884_), .C2(new_n885_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n887_), .A2(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n355_), .B1(new_n882_), .B2(new_n890_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n709_), .A2(new_n288_), .A3(new_n758_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(KEYINPUT54), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n694_), .B(new_n831_), .C1(new_n891_), .C2(new_n893_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(KEYINPUT123), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n639_), .ZN(new_n896_));
  INV_X1    g695(.A(G113gat), .ZN(new_n897_));
  XOR2_X1   g696(.A(new_n894_), .B(KEYINPUT59), .Z(new_n898_));
  AOI21_X1  g697(.A(new_n897_), .B1(new_n639_), .B2(KEYINPUT124), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n899_), .B1(KEYINPUT124), .B2(new_n897_), .ZN(new_n900_));
  AOI22_X1  g699(.A1(new_n896_), .A2(new_n897_), .B1(new_n898_), .B2(new_n900_), .ZN(G1340gat));
  XNOR2_X1  g700(.A(new_n894_), .B(KEYINPUT59), .ZN(new_n902_));
  OAI21_X1  g701(.A(G120gat), .B1(new_n902_), .B2(new_n289_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT60), .ZN(new_n904_));
  AOI21_X1  g703(.A(G120gat), .B1(new_n288_), .B2(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n905_), .B1(new_n904_), .B2(G120gat), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n895_), .A2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n903_), .A2(new_n907_), .ZN(G1341gat));
  OAI21_X1  g707(.A(G127gat), .B1(new_n902_), .B2(new_n659_), .ZN(new_n909_));
  INV_X1    g708(.A(G127gat), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n895_), .A2(new_n910_), .A3(new_n355_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n911_), .ZN(G1342gat));
  OAI21_X1  g711(.A(G134gat), .B1(new_n902_), .B2(new_n326_), .ZN(new_n913_));
  INV_X1    g712(.A(G134gat), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n895_), .A2(new_n914_), .A3(new_n655_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n913_), .A2(new_n915_), .ZN(G1343gat));
  OR2_X1    g715(.A1(new_n891_), .A2(new_n893_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n830_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n741_), .A2(new_n694_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n917_), .A2(new_n918_), .A3(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(new_n642_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(KEYINPUT125), .B(G141gat), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n921_), .B(new_n922_), .ZN(G1344gat));
  NOR2_X1   g722(.A1(new_n920_), .A2(new_n289_), .ZN(new_n924_));
  INV_X1    g723(.A(G148gat), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n924_), .B(new_n925_), .ZN(G1345gat));
  NOR2_X1   g725(.A1(new_n920_), .A2(new_n659_), .ZN(new_n927_));
  XOR2_X1   g726(.A(KEYINPUT61), .B(G155gat), .Z(new_n928_));
  XNOR2_X1  g727(.A(new_n927_), .B(new_n928_), .ZN(G1346gat));
  INV_X1    g728(.A(G162gat), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n920_), .A2(new_n930_), .A3(new_n710_), .ZN(new_n931_));
  OR2_X1    g730(.A1(new_n920_), .A2(new_n668_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n931_), .B1(new_n930_), .B2(new_n932_), .ZN(G1347gat));
  NOR3_X1   g732(.A1(new_n416_), .A2(new_n591_), .A3(new_n589_), .ZN(new_n934_));
  AND2_X1   g733(.A1(new_n934_), .A2(new_n639_), .ZN(new_n935_));
  OAI211_X1 g734(.A(new_n694_), .B(new_n935_), .C1(new_n891_), .C2(new_n893_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(G169gat), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT62), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n937_), .A2(new_n938_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n936_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n940_));
  NAND4_X1  g739(.A1(new_n917_), .A2(new_n387_), .A3(new_n694_), .A4(new_n935_), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n939_), .A2(new_n940_), .A3(new_n941_), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(new_n944_));
  NAND4_X1  g743(.A1(new_n939_), .A2(KEYINPUT126), .A3(new_n940_), .A4(new_n941_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(G1348gat));
  NAND3_X1  g745(.A1(new_n917_), .A2(new_n694_), .A3(new_n934_), .ZN(new_n947_));
  OAI21_X1  g746(.A(G176gat), .B1(new_n947_), .B2(new_n289_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n288_), .A2(new_n388_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n948_), .B1(new_n947_), .B2(new_n949_), .ZN(G1349gat));
  NOR3_X1   g749(.A1(new_n947_), .A2(new_n445_), .A3(new_n659_), .ZN(new_n951_));
  OR2_X1    g750(.A1(new_n947_), .A2(new_n659_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n951_), .B1(new_n373_), .B2(new_n952_), .ZN(G1350gat));
  OAI21_X1  g752(.A(G190gat), .B1(new_n947_), .B2(new_n326_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n655_), .A2(new_n371_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n954_), .B1(new_n947_), .B2(new_n955_), .ZN(G1351gat));
  NOR2_X1   g755(.A1(new_n589_), .A2(new_n591_), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n917_), .A2(new_n919_), .A3(new_n957_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n958_), .A2(new_n642_), .ZN(new_n959_));
  INV_X1    g758(.A(G197gat), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n959_), .B(new_n960_), .ZN(G1352gat));
  NOR2_X1   g760(.A1(new_n958_), .A2(new_n289_), .ZN(new_n962_));
  INV_X1    g761(.A(G204gat), .ZN(new_n963_));
  XNOR2_X1  g762(.A(new_n962_), .B(new_n963_), .ZN(G1353gat));
  NOR2_X1   g763(.A1(new_n958_), .A2(new_n659_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n966_));
  AND2_X1   g765(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n967_));
  OAI21_X1  g766(.A(new_n965_), .B1(new_n966_), .B2(new_n967_), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n968_), .B1(new_n965_), .B2(new_n966_), .ZN(G1354gat));
  INV_X1    g768(.A(new_n958_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n970_), .A2(new_n655_), .ZN(new_n971_));
  INV_X1    g770(.A(G218gat), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n709_), .A2(G218gat), .ZN(new_n973_));
  XNOR2_X1  g772(.A(new_n973_), .B(KEYINPUT127), .ZN(new_n974_));
  AOI22_X1  g773(.A1(new_n971_), .A2(new_n972_), .B1(new_n970_), .B2(new_n974_), .ZN(G1355gat));
endmodule


