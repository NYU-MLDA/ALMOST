//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 1 0 0 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n579_, new_n580_, new_n581_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n587_, new_n588_,
    new_n589_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n621_,
    new_n622_, new_n623_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n644_, new_n645_, new_n646_, new_n648_, new_n649_, new_n650_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n813_, new_n815_, new_n816_, new_n818_,
    new_n819_, new_n820_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n843_, new_n844_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  OR2_X1    g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204_));
  AOI22_X1  g003(.A1(new_n203_), .A2(new_n204_), .B1(G169gat), .B2(G176gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT82), .B(G176gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT22), .B(G169gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n205_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G169gat), .ZN(new_n210_));
  INV_X1    g009(.A(G176gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n212_), .A2(KEYINPUT24), .ZN(new_n213_));
  AND2_X1   g012(.A1(new_n203_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT25), .B(G183gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT26), .B(G190gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n214_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n212_), .A2(KEYINPUT24), .A3(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT81), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n209_), .B1(new_n218_), .B2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G71gat), .B(G99gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(G43gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n222_), .B(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G227gat), .A2(G233gat), .ZN(new_n226_));
  XOR2_X1   g025(.A(new_n226_), .B(G15gat), .Z(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT30), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n225_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n225_), .A2(new_n228_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT83), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n229_), .A2(KEYINPUT83), .A3(new_n230_), .ZN(new_n234_));
  XOR2_X1   g033(.A(G127gat), .B(G134gat), .Z(new_n235_));
  XOR2_X1   g034(.A(G113gat), .B(G120gat), .Z(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(new_n237_), .B(KEYINPUT31), .Z(new_n238_));
  NAND3_X1  g037(.A1(new_n233_), .A2(new_n234_), .A3(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n234_), .A2(new_n238_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n241_), .A2(KEYINPUT84), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT84), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n243_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT92), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT28), .B(G22gat), .ZN(new_n247_));
  INV_X1    g046(.A(G50gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G155gat), .A2(G162gat), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(G155gat), .A2(G162gat), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT85), .ZN(new_n256_));
  NOR2_X1   g055(.A1(G141gat), .A2(G148gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT3), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT2), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G141gat), .A2(G148gat), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n259_), .B(new_n260_), .C1(new_n261_), .C2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n254_), .B1(new_n256_), .B2(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n253_), .B1(KEYINPUT1), .B2(new_n251_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n265_), .B1(KEYINPUT1), .B2(new_n251_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n257_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n266_), .A2(new_n262_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT29), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n264_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT86), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n270_), .A2(KEYINPUT86), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n250_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n273_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n275_), .A2(new_n249_), .A3(new_n271_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT87), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT87), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n274_), .A2(new_n276_), .A3(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(G211gat), .B(G218gat), .Z(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT21), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT88), .ZN(new_n283_));
  INV_X1    g082(.A(G204gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n283_), .B1(new_n284_), .B2(G197gat), .ZN(new_n285_));
  INV_X1    g084(.A(G197gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n286_), .A2(KEYINPUT88), .A3(G204gat), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n285_), .B(new_n287_), .C1(new_n286_), .C2(G204gat), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n282_), .B1(KEYINPUT89), .B2(new_n288_), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n288_), .A2(KEYINPUT89), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n288_), .A2(KEYINPUT21), .ZN(new_n292_));
  XOR2_X1   g091(.A(G197gat), .B(G204gat), .Z(new_n293_));
  AOI21_X1  g092(.A(new_n281_), .B1(new_n293_), .B2(KEYINPUT21), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n291_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n264_), .A2(new_n268_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT29), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT90), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n299_), .A2(G228gat), .A3(G233gat), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n296_), .A2(new_n298_), .A3(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G228gat), .A2(G233gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT90), .ZN(new_n303_));
  AOI22_X1  g102(.A1(new_n296_), .A2(new_n298_), .B1(new_n303_), .B2(new_n300_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G78gat), .B(G106gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT91), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  OR3_X1    g106(.A1(new_n301_), .A2(new_n304_), .A3(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n307_), .B1(new_n301_), .B2(new_n304_), .ZN(new_n309_));
  AOI22_X1  g108(.A1(new_n278_), .A2(new_n280_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n305_), .B1(new_n301_), .B2(new_n304_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n308_), .A2(new_n277_), .A3(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n246_), .B1(new_n310_), .B2(new_n313_), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n278_), .A2(new_n280_), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n308_), .A2(new_n309_), .ZN(new_n316_));
  OAI211_X1 g115(.A(KEYINPUT92), .B(new_n312_), .C1(new_n315_), .C2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n314_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n237_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n297_), .A2(new_n320_), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n321_), .A2(KEYINPUT4), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G225gat), .A2(G233gat), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n237_), .A2(new_n264_), .A3(new_n268_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n321_), .A2(KEYINPUT4), .A3(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n322_), .A2(new_n323_), .A3(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT99), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G1gat), .B(G29gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(G85gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT0), .B(G57gat), .ZN(new_n330_));
  XOR2_X1   g129(.A(new_n329_), .B(new_n330_), .Z(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n323_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n321_), .A2(new_n333_), .A3(new_n324_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n327_), .A2(new_n332_), .A3(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n323_), .B1(new_n322_), .B2(new_n325_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n333_), .B1(new_n321_), .B2(new_n324_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n331_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT33), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT33), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n340_), .B(new_n331_), .C1(new_n336_), .C2(new_n337_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n335_), .A2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT20), .B1(new_n296_), .B2(new_n222_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT93), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n219_), .A2(KEYINPUT24), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n346_), .A2(KEYINPUT94), .B1(new_n210_), .B2(new_n211_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n347_), .B1(KEYINPUT94), .B2(new_n346_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT95), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n214_), .A2(new_n349_), .ZN(new_n350_));
  AND3_X1   g149(.A1(new_n203_), .A2(new_n213_), .A3(new_n349_), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n217_), .B(new_n348_), .C1(new_n350_), .C2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n207_), .B(KEYINPUT96), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(new_n206_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n205_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n352_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n296_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT93), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n358_), .B(KEYINPUT20), .C1(new_n296_), .C2(new_n222_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n345_), .A2(new_n357_), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT19), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n296_), .A2(new_n222_), .ZN(new_n364_));
  OAI211_X1 g163(.A(KEYINPUT20), .B(new_n364_), .C1(new_n356_), .C2(new_n296_), .ZN(new_n365_));
  OR2_X1    g164(.A1(new_n365_), .A2(new_n362_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n363_), .A2(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(G8gat), .B(G36gat), .Z(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G64gat), .B(G92gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n367_), .A2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n363_), .A2(new_n366_), .A3(new_n372_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n374_), .A2(KEYINPUT98), .A3(new_n375_), .ZN(new_n376_));
  OR3_X1    g175(.A1(new_n367_), .A2(KEYINPUT98), .A3(new_n373_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n343_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  OR3_X1    g177(.A1(new_n336_), .A2(new_n331_), .A3(new_n337_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(new_n338_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n372_), .A2(KEYINPUT32), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n380_), .B1(new_n367_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n365_), .A2(new_n362_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n384_), .B1(new_n360_), .B2(new_n362_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT100), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n386_), .A3(new_n382_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n382_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT100), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n383_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n319_), .B1(new_n378_), .B2(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n380_), .B1(new_n314_), .B2(new_n317_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT27), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n376_), .A2(new_n377_), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n385_), .A2(new_n373_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n395_), .A2(new_n375_), .A3(KEYINPUT27), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n392_), .A2(new_n394_), .A3(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n245_), .B1(new_n391_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n394_), .A2(new_n396_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n241_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n380_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NOR3_X1   g201(.A1(new_n399_), .A2(new_n402_), .A3(new_n318_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n398_), .A2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G190gat), .B(G218gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G134gat), .B(G162gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT36), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G232gat), .A2(G233gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT34), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT35), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(KEYINPUT35), .ZN(new_n412_));
  INV_X1    g211(.A(G106gat), .ZN(new_n413_));
  OR2_X1    g212(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT64), .ZN(new_n415_));
  NAND2_X1  g214(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n414_), .A2(new_n415_), .A3(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n415_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n413_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  XOR2_X1   g218(.A(G85gat), .B(G92gat), .Z(new_n420_));
  NAND2_X1  g219(.A1(G99gat), .A2(G106gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT6), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT6), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n423_), .A2(G99gat), .A3(G106gat), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n420_), .A2(KEYINPUT9), .B1(new_n422_), .B2(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(KEYINPUT65), .B(G85gat), .Z(new_n426_));
  INV_X1    g225(.A(KEYINPUT9), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n426_), .A2(new_n427_), .A3(G92gat), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n419_), .A2(new_n425_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT66), .ZN(new_n430_));
  INV_X1    g229(.A(G99gat), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n430_), .A2(new_n431_), .A3(new_n413_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT7), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n422_), .A2(new_n424_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT7), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n430_), .A2(new_n435_), .A3(new_n431_), .A4(new_n413_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n433_), .A2(new_n434_), .A3(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT8), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n437_), .A2(new_n438_), .A3(new_n420_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n438_), .B1(new_n437_), .B2(new_n420_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n429_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT67), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT67), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n429_), .B(new_n443_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G29gat), .B(G36gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G43gat), .B(G50gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n412_), .B1(new_n445_), .B2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n411_), .B1(new_n449_), .B2(KEYINPUT73), .ZN(new_n450_));
  NOR3_X1   g249(.A1(new_n439_), .A2(new_n440_), .A3(KEYINPUT69), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT69), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n437_), .A2(new_n420_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT8), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n437_), .A2(new_n438_), .A3(new_n420_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n452_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n429_), .B1(new_n451_), .B2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n448_), .B(KEYINPUT15), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n449_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n450_), .A2(new_n460_), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n449_), .B(new_n459_), .C1(KEYINPUT73), .C2(new_n411_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n407_), .A2(KEYINPUT36), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n461_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n463_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n408_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT37), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n468_), .B1(new_n464_), .B2(KEYINPUT74), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n467_), .B(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G57gat), .B(G64gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT11), .ZN(new_n473_));
  XOR2_X1   g272(.A(G71gat), .B(G78gat), .Z(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n472_), .A2(KEYINPUT11), .ZN(new_n476_));
  OR2_X1    g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n473_), .A2(new_n474_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G231gat), .A2(G233gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(KEYINPUT75), .B(G8gat), .ZN(new_n482_));
  INV_X1    g281(.A(G1gat), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT14), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G15gat), .B(G22gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G1gat), .B(G8gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n484_), .A2(new_n485_), .A3(new_n487_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n481_), .B(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT77), .ZN(new_n493_));
  XOR2_X1   g292(.A(G127gat), .B(G155gat), .Z(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G183gat), .B(G211gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT17), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n493_), .B(new_n500_), .ZN(new_n501_));
  OR3_X1    g300(.A1(new_n492_), .A2(KEYINPUT17), .A3(new_n499_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n471_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G113gat), .B(G141gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G169gat), .B(G197gat), .ZN(new_n506_));
  XOR2_X1   g305(.A(new_n505_), .B(new_n506_), .Z(new_n507_));
  NAND2_X1  g306(.A1(new_n491_), .A2(new_n448_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT78), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n491_), .A2(new_n448_), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G229gat), .A2(G233gat), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n458_), .A2(new_n490_), .A3(new_n489_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n509_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n512_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n514_), .A2(KEYINPUT79), .A3(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT80), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT80), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n514_), .A2(KEYINPUT79), .A3(new_n520_), .A4(new_n517_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n507_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n519_), .A2(new_n521_), .A3(new_n507_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT13), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n527_), .A2(KEYINPUT72), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT72), .B(KEYINPUT13), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n454_), .A2(new_n455_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n443_), .B1(new_n530_), .B2(new_n429_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n444_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n479_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n479_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n442_), .A2(new_n534_), .A3(new_n444_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n533_), .A2(KEYINPUT68), .A3(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G230gat), .A2(G233gat), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n536_), .B(new_n538_), .C1(KEYINPUT68), .C2(new_n535_), .ZN(new_n539_));
  XOR2_X1   g338(.A(KEYINPUT70), .B(KEYINPUT12), .Z(new_n540_));
  NAND2_X1  g339(.A1(new_n535_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n477_), .A2(KEYINPUT12), .A3(new_n478_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n457_), .A2(new_n543_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n541_), .A2(new_n537_), .A3(new_n544_), .A4(new_n533_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n539_), .A2(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(G120gat), .B(G148gat), .Z(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G176gat), .B(G204gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n546_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n551_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n539_), .A2(new_n545_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  MUX2_X1   g354(.A(new_n528_), .B(new_n529_), .S(new_n555_), .Z(new_n556_));
  NOR4_X1   g355(.A1(new_n404_), .A2(new_n504_), .A3(new_n526_), .A4(new_n556_), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n557_), .A2(KEYINPUT101), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(KEYINPUT101), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n558_), .A2(new_n483_), .A3(new_n380_), .A4(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT38), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n404_), .A2(new_n467_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n556_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n563_), .A2(new_n525_), .A3(new_n564_), .A4(new_n503_), .ZN(new_n565_));
  OAI21_X1  g364(.A(G1gat), .B1(new_n565_), .B2(new_n401_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n560_), .A2(new_n561_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n562_), .A2(new_n566_), .A3(new_n567_), .ZN(G1324gat));
  NAND4_X1  g367(.A1(new_n558_), .A2(new_n399_), .A3(new_n482_), .A4(new_n559_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT102), .ZN(new_n570_));
  INV_X1    g369(.A(new_n399_), .ZN(new_n571_));
  OAI21_X1  g370(.A(G8gat), .B1(new_n565_), .B2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT39), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT40), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n570_), .A2(KEYINPUT40), .A3(new_n573_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(G1325gat));
  INV_X1    g377(.A(new_n245_), .ZN(new_n579_));
  OAI21_X1  g378(.A(G15gat), .B1(new_n565_), .B2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n580_), .B(KEYINPUT103), .Z(new_n581_));
  OR2_X1    g380(.A1(new_n581_), .A2(KEYINPUT41), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(KEYINPUT41), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n558_), .A2(new_n559_), .ZN(new_n584_));
  OR3_X1    g383(.A1(new_n584_), .A2(G15gat), .A3(new_n579_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n582_), .A2(new_n583_), .A3(new_n585_), .ZN(G1326gat));
  OAI21_X1  g385(.A(G22gat), .B1(new_n565_), .B2(new_n319_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT42), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n319_), .A2(G22gat), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n588_), .B1(new_n584_), .B2(new_n589_), .ZN(G1327gat));
  NAND2_X1  g389(.A1(new_n391_), .A2(new_n397_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(new_n579_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n403_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT43), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n594_), .A2(KEYINPUT104), .A3(new_n595_), .A4(new_n470_), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n595_), .B(new_n470_), .C1(new_n398_), .C2(new_n403_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT104), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(KEYINPUT43), .B1(new_n404_), .B2(new_n471_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n596_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  NOR3_X1   g400(.A1(new_n556_), .A2(new_n526_), .A3(new_n503_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT44), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(G29gat), .B1(new_n605_), .B2(new_n401_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n503_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(new_n467_), .ZN(new_n608_));
  OR4_X1    g407(.A1(new_n404_), .A2(new_n526_), .A3(new_n556_), .A4(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n401_), .A2(G29gat), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT105), .Z(new_n611_));
  OAI21_X1  g410(.A(new_n606_), .B1(new_n609_), .B2(new_n611_), .ZN(G1328gat));
  OAI21_X1  g411(.A(G36gat), .B1(new_n605_), .B2(new_n571_), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n609_), .A2(G36gat), .A3(new_n571_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n614_), .B(KEYINPUT45), .Z(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT46), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n613_), .A2(KEYINPUT46), .A3(new_n615_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(G1329gat));
  NAND2_X1  g419(.A1(new_n400_), .A2(G43gat), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n609_), .A2(new_n579_), .ZN(new_n622_));
  OAI22_X1  g421(.A1(new_n605_), .A2(new_n621_), .B1(G43gat), .B2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g423(.A(KEYINPUT106), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n603_), .B(KEYINPUT44), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(new_n318_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n625_), .B1(new_n627_), .B2(G50gat), .ZN(new_n628_));
  AOI211_X1 g427(.A(KEYINPUT106), .B(new_n248_), .C1(new_n626_), .C2(new_n318_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n318_), .A2(new_n248_), .ZN(new_n630_));
  OAI22_X1  g429(.A1(new_n628_), .A2(new_n629_), .B1(new_n609_), .B2(new_n630_), .ZN(G1331gat));
  NAND4_X1  g430(.A1(new_n563_), .A2(new_n526_), .A3(new_n556_), .A4(new_n503_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G57gat), .B1(new_n632_), .B2(new_n401_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n594_), .A2(new_n526_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n634_), .A2(new_n564_), .A3(new_n504_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT107), .Z(new_n636_));
  OR2_X1    g435(.A1(new_n401_), .A2(G57gat), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n633_), .B1(new_n636_), .B2(new_n637_), .ZN(G1332gat));
  OAI21_X1  g437(.A(G64gat), .B1(new_n632_), .B2(new_n571_), .ZN(new_n639_));
  XOR2_X1   g438(.A(KEYINPUT108), .B(KEYINPUT48), .Z(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n571_), .A2(G64gat), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n641_), .B1(new_n636_), .B2(new_n642_), .ZN(G1333gat));
  OAI21_X1  g442(.A(G71gat), .B1(new_n632_), .B2(new_n579_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT49), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n579_), .A2(G71gat), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n645_), .B1(new_n636_), .B2(new_n646_), .ZN(G1334gat));
  OAI21_X1  g446(.A(G78gat), .B1(new_n632_), .B2(new_n319_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT50), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n319_), .A2(G78gat), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n649_), .B1(new_n636_), .B2(new_n650_), .ZN(G1335gat));
  OR3_X1    g450(.A1(new_n634_), .A2(new_n564_), .A3(new_n608_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(G85gat), .B1(new_n653_), .B2(new_n380_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n564_), .A2(new_n525_), .A3(new_n503_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n601_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n426_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n656_), .A2(new_n401_), .A3(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n654_), .A2(new_n658_), .ZN(G1336gat));
  INV_X1    g458(.A(G92gat), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n660_), .B1(new_n652_), .B2(new_n571_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT109), .Z(new_n662_));
  NOR3_X1   g461(.A1(new_n656_), .A2(new_n660_), .A3(new_n571_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1337gat));
  OAI21_X1  g463(.A(G99gat), .B1(new_n656_), .B2(new_n579_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n400_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n665_), .B(KEYINPUT110), .C1(new_n652_), .C2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g467(.A1(new_n653_), .A2(new_n413_), .A3(new_n318_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT52), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n601_), .A2(KEYINPUT111), .A3(new_n318_), .A4(new_n655_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n671_), .A2(G106gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n601_), .A2(new_n318_), .A3(new_n655_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT111), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n670_), .B1(new_n672_), .B2(new_n675_), .ZN(new_n676_));
  AND4_X1   g475(.A1(new_n670_), .A2(new_n675_), .A3(G106gat), .A4(new_n671_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n669_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT53), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT53), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n680_), .B(new_n669_), .C1(new_n676_), .C2(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(G1339gat));
  NAND4_X1  g481(.A1(new_n571_), .A2(new_n319_), .A3(new_n380_), .A4(new_n400_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT118), .Z(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT114), .ZN(new_n686_));
  AOI22_X1  g485(.A1(new_n479_), .A2(new_n445_), .B1(new_n457_), .B2(new_n543_), .ZN(new_n687_));
  AOI211_X1 g486(.A(new_n686_), .B(new_n537_), .C1(new_n687_), .C2(new_n541_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n541_), .A2(new_n533_), .A3(new_n544_), .ZN(new_n689_));
  AOI21_X1  g488(.A(KEYINPUT114), .B1(new_n689_), .B2(new_n538_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n545_), .A2(KEYINPUT55), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT55), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n687_), .A2(new_n693_), .A3(new_n537_), .A4(new_n541_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n692_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT115), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n691_), .A2(new_n695_), .A3(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n689_), .A2(new_n538_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(new_n686_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n689_), .A2(KEYINPUT114), .A3(new_n538_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n692_), .A2(new_n694_), .ZN(new_n702_));
  AOI21_X1  g501(.A(KEYINPUT115), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  OAI211_X1 g502(.A(KEYINPUT56), .B(new_n551_), .C1(new_n697_), .C2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT117), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n696_), .B1(new_n691_), .B2(new_n695_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n701_), .A2(KEYINPUT115), .A3(new_n702_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n709_), .A2(KEYINPUT117), .A3(KEYINPUT56), .A4(new_n551_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n551_), .B1(new_n697_), .B2(new_n703_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT56), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n706_), .A2(new_n710_), .A3(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n507_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n509_), .A2(new_n513_), .A3(new_n515_), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n715_), .B(new_n716_), .C1(new_n511_), .C2(new_n513_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT116), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n718_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n514_), .A2(new_n517_), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n719_), .B(new_n720_), .C1(new_n721_), .C2(new_n715_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n554_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n714_), .A2(KEYINPUT58), .A3(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(KEYINPUT58), .B1(new_n714_), .B2(new_n724_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n726_), .A2(new_n727_), .A3(new_n471_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n467_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n524_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n554_), .B1(new_n730_), .B2(new_n522_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n713_), .B2(new_n704_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n555_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n722_), .A2(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n729_), .B1(new_n732_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT57), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n723_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT56), .B1(new_n709_), .B2(new_n551_), .ZN(new_n739_));
  AOI211_X1 g538(.A(new_n712_), .B(new_n553_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n738_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n734_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n743_), .A2(KEYINPUT57), .A3(new_n729_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n737_), .A2(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n607_), .B1(new_n728_), .B2(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(KEYINPUT112), .B1(new_n525_), .B2(new_n607_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n523_), .A2(new_n748_), .A3(new_n524_), .A4(new_n503_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n471_), .A2(new_n564_), .A3(new_n747_), .A4(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT113), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT54), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT54), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n750_), .A2(new_n751_), .A3(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n750_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT113), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n685_), .B1(new_n746_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(G113gat), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(new_n761_), .A3(new_n525_), .ZN(new_n762_));
  AOI21_X1  g561(.A(KEYINPUT57), .B1(new_n743_), .B2(new_n729_), .ZN(new_n763_));
  AOI211_X1 g562(.A(new_n736_), .B(new_n467_), .C1(new_n741_), .C2(new_n742_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n714_), .A2(new_n724_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT58), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n768_), .A2(new_n470_), .A3(new_n725_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n503_), .B1(new_n765_), .B2(new_n769_), .ZN(new_n770_));
  AOI22_X1  g569(.A1(new_n753_), .A2(new_n755_), .B1(KEYINPUT113), .B2(new_n757_), .ZN(new_n771_));
  OAI211_X1 g570(.A(KEYINPUT119), .B(new_n684_), .C1(new_n770_), .C2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT59), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n746_), .A2(new_n759_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n775_), .A2(KEYINPUT119), .A3(KEYINPUT59), .A4(new_n684_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n526_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n762_), .B1(new_n777_), .B2(new_n761_), .ZN(G1340gat));
  AOI21_X1  g577(.A(new_n564_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n779_));
  INV_X1    g578(.A(G120gat), .ZN(new_n780_));
  INV_X1    g579(.A(new_n760_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n780_), .B1(new_n564_), .B2(KEYINPUT60), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n780_), .A2(KEYINPUT60), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n782_), .B1(KEYINPUT120), .B2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n784_), .B1(KEYINPUT120), .B2(new_n782_), .ZN(new_n785_));
  OAI22_X1  g584(.A1(new_n779_), .A2(new_n780_), .B1(new_n781_), .B2(new_n785_), .ZN(G1341gat));
  INV_X1    g585(.A(G127gat), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n787_), .B1(new_n781_), .B2(new_n607_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT121), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT121), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n790_), .B(new_n787_), .C1(new_n781_), .C2(new_n607_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n774_), .A2(new_n776_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n607_), .A2(new_n787_), .ZN(new_n793_));
  AOI22_X1  g592(.A1(new_n789_), .A2(new_n791_), .B1(new_n792_), .B2(new_n793_), .ZN(G1342gat));
  INV_X1    g593(.A(G134gat), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n471_), .A2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT59), .B1(new_n760_), .B2(KEYINPUT119), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n772_), .A2(new_n773_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n796_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(G134gat), .B1(new_n760_), .B2(new_n467_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n799_), .A2(KEYINPUT122), .A3(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT122), .ZN(new_n803_));
  INV_X1    g602(.A(new_n796_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n803_), .B1(new_n805_), .B2(new_n800_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n802_), .A2(new_n806_), .ZN(G1343gat));
  NOR2_X1   g606(.A1(new_n770_), .A2(new_n771_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n579_), .A2(new_n318_), .A3(new_n380_), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n808_), .A2(new_n399_), .A3(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n525_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n556_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g613(.A1(new_n810_), .A2(new_n503_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(KEYINPUT61), .B(G155gat), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n815_), .B(new_n816_), .ZN(G1346gat));
  INV_X1    g616(.A(G162gat), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n810_), .A2(new_n818_), .A3(new_n467_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n810_), .A2(new_n470_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n819_), .B1(new_n820_), .B2(new_n818_), .ZN(G1347gat));
  NOR4_X1   g620(.A1(new_n579_), .A2(new_n571_), .A3(new_n318_), .A4(new_n380_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n525_), .B(new_n822_), .C1(new_n770_), .C2(new_n771_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n823_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n775_), .A2(new_n353_), .A3(new_n525_), .A4(new_n822_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT62), .B1(new_n823_), .B2(G169gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT123), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n827_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT123), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n829_), .A2(new_n830_), .A3(new_n825_), .A4(new_n824_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n828_), .A2(new_n831_), .ZN(G1348gat));
  NAND2_X1  g631(.A1(new_n775_), .A2(new_n822_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n556_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n835_), .A2(new_n211_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n836_), .B1(new_n206_), .B2(new_n835_), .ZN(G1349gat));
  INV_X1    g636(.A(G183gat), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT124), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n834_), .A2(new_n215_), .A3(new_n503_), .A4(new_n839_), .ZN(new_n840_));
  OAI22_X1  g639(.A1(new_n833_), .A2(new_n607_), .B1(KEYINPUT124), .B2(G183gat), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(G1350gat));
  OAI21_X1  g641(.A(G190gat), .B1(new_n833_), .B2(new_n471_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n467_), .A2(new_n216_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n833_), .B2(new_n844_), .ZN(G1351gat));
  NAND3_X1  g644(.A1(new_n579_), .A2(new_n392_), .A3(new_n399_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n808_), .A2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n525_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n556_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g650(.A(KEYINPUT63), .ZN(new_n852_));
  INV_X1    g651(.A(G211gat), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n503_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  XOR2_X1   g653(.A(new_n854_), .B(KEYINPUT125), .Z(new_n855_));
  NAND2_X1  g654(.A1(new_n847_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n852_), .A2(new_n853_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n856_), .B(new_n857_), .ZN(G1354gat));
  NOR3_X1   g657(.A1(new_n808_), .A2(new_n729_), .A3(new_n846_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT126), .ZN(new_n860_));
  OR2_X1    g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(G218gat), .B1(new_n859_), .B2(new_n860_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n470_), .A2(G218gat), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(KEYINPUT127), .ZN(new_n864_));
  AOI22_X1  g663(.A1(new_n861_), .A2(new_n862_), .B1(new_n847_), .B2(new_n864_), .ZN(G1355gat));
endmodule


