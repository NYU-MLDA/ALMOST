//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 0 1 1 0 0 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 0 0 1 0 0 1 1 0 0 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n887_, new_n889_,
    new_n890_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT87), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT87), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n207_), .B1(G169gat), .B2(G176gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209_));
  NAND4_X1  g008(.A1(new_n206_), .A2(KEYINPUT24), .A3(new_n208_), .A4(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT25), .B(G183gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT26), .B(G190gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  AND2_X1   g012(.A1(new_n206_), .A2(new_n208_), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n210_), .B(new_n213_), .C1(new_n214_), .C2(KEYINPUT24), .ZN(new_n215_));
  INV_X1    g014(.A(G183gat), .ZN(new_n216_));
  INV_X1    g015(.A(G190gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT23), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT23), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n220_), .A2(G183gat), .A3(G190gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT88), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n222_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n219_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(G169gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n228_), .B1(new_n218_), .B2(new_n221_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n227_), .B1(new_n229_), .B2(KEYINPUT89), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT89), .ZN(new_n231_));
  AOI211_X1 g030(.A(new_n231_), .B(new_n228_), .C1(new_n218_), .C2(new_n221_), .ZN(new_n232_));
  OAI22_X1  g031(.A1(new_n215_), .A2(new_n225_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT90), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  OAI221_X1 g034(.A(KEYINPUT90), .B1(new_n230_), .B2(new_n232_), .C1(new_n225_), .C2(new_n215_), .ZN(new_n236_));
  OR2_X1    g035(.A1(G197gat), .A2(G204gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G197gat), .A2(G204gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT21), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n237_), .A2(KEYINPUT21), .A3(new_n238_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G211gat), .B(G218gat), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n242_), .A2(new_n243_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n235_), .A2(new_n236_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT20), .ZN(new_n249_));
  INV_X1    g048(.A(G176gat), .ZN(new_n250_));
  INV_X1    g049(.A(G169gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT22), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT22), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(G169gat), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n252_), .A2(new_n254_), .A3(KEYINPUT102), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT102), .B1(new_n252_), .B2(new_n254_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n250_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n257_), .B(new_n209_), .C1(new_n225_), .C2(new_n228_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT24), .ZN(new_n259_));
  AOI22_X1  g058(.A1(new_n218_), .A2(new_n221_), .B1(new_n259_), .B2(new_n205_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n209_), .A2(KEYINPUT24), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT101), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n214_), .A2(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n261_), .A2(KEYINPUT101), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n213_), .B(new_n260_), .C1(new_n263_), .C2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n258_), .A2(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n249_), .B1(new_n266_), .B2(new_n246_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n204_), .B1(new_n248_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G8gat), .B(G36gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT18), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G64gat), .B(G92gat), .ZN(new_n272_));
  XOR2_X1   g071(.A(new_n271_), .B(new_n272_), .Z(new_n273_));
  NAND3_X1  g072(.A1(new_n258_), .A2(new_n247_), .A3(new_n265_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT103), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n258_), .A2(new_n247_), .A3(KEYINPUT103), .A4(new_n265_), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n276_), .A2(new_n204_), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n235_), .A2(new_n236_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n249_), .B1(new_n279_), .B2(new_n246_), .ZN(new_n280_));
  AND3_X1   g079(.A1(new_n278_), .A2(KEYINPUT104), .A3(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(KEYINPUT104), .B1(new_n278_), .B2(new_n280_), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n269_), .B(new_n273_), .C1(new_n281_), .C2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT27), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n248_), .A2(new_n267_), .A3(new_n204_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n247_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n274_), .ZN(new_n287_));
  NOR3_X1   g086(.A1(new_n286_), .A2(new_n249_), .A3(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n285_), .B1(new_n288_), .B2(new_n204_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n273_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n284_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n283_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT108), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT108), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n283_), .A2(new_n291_), .A3(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n269_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(new_n290_), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n297_), .A2(new_n283_), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n293_), .B(new_n295_), .C1(new_n298_), .C2(KEYINPUT27), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G227gat), .A2(G233gat), .ZN(new_n300_));
  INV_X1    g099(.A(G15gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(G71gat), .ZN(new_n303_));
  INV_X1    g102(.A(G99gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT91), .B(G43gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT30), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n279_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n235_), .A2(new_n236_), .A3(KEYINPUT30), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n307_), .A2(KEYINPUT92), .A3(new_n309_), .A4(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n305_), .B(new_n306_), .Z(new_n312_));
  NAND3_X1  g111(.A1(new_n309_), .A2(KEYINPUT92), .A3(new_n310_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(KEYINPUT92), .B1(new_n309_), .B2(new_n310_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n311_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT93), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G127gat), .B(G134gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G113gat), .B(G120gat), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n319_), .B(new_n320_), .Z(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT31), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n318_), .A2(new_n322_), .ZN(new_n323_));
  XOR2_X1   g122(.A(G141gat), .B(G148gat), .Z(new_n324_));
  NOR2_X1   g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT1), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G155gat), .A2(G162gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT94), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT94), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n329_), .A2(G155gat), .A3(G162gat), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n326_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT95), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n325_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n328_), .A2(new_n330_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT1), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT95), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n333_), .A2(new_n336_), .A3(KEYINPUT96), .ZN(new_n337_));
  INV_X1    g136(.A(new_n334_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(new_n326_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(KEYINPUT96), .B1(new_n333_), .B2(new_n336_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n324_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT106), .ZN(new_n343_));
  INV_X1    g142(.A(G141gat), .ZN(new_n344_));
  INV_X1    g143(.A(G148gat), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT98), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n346_), .B(KEYINPUT2), .Z(new_n347_));
  NAND3_X1  g146(.A1(new_n344_), .A2(new_n345_), .A3(KEYINPUT97), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n348_), .B(KEYINPUT3), .Z(new_n349_));
  AOI211_X1 g148(.A(new_n338_), .B(new_n325_), .C1(new_n347_), .C2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n342_), .A2(new_n343_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n321_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n352_), .A2(KEYINPUT105), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT105), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n333_), .A2(new_n336_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT96), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n358_), .A2(new_n339_), .A3(new_n337_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n350_), .B1(new_n359_), .B2(new_n324_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n355_), .B1(new_n360_), .B2(new_n343_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n342_), .A2(new_n355_), .A3(new_n351_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(new_n321_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n354_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G225gat), .A2(G233gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G1gat), .B(G29gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(G85gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT0), .B(G57gat), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n368_), .B(new_n369_), .Z(new_n370_));
  INV_X1    g169(.A(KEYINPUT4), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n352_), .A2(KEYINPUT105), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n372_), .A2(new_n362_), .A3(new_n321_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n371_), .B1(new_n373_), .B2(new_n354_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n342_), .A2(new_n351_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n375_), .A2(new_n371_), .A3(new_n321_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n365_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n366_), .B(new_n370_), .C1(new_n374_), .C2(new_n378_), .ZN(new_n379_));
  OAI211_X1 g178(.A(KEYINPUT93), .B(new_n311_), .C1(new_n314_), .C2(new_n315_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n318_), .A2(new_n380_), .A3(new_n322_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n370_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n378_), .B1(new_n364_), .B2(KEYINPUT4), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n377_), .B1(new_n373_), .B2(new_n354_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n382_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n323_), .A2(new_n379_), .A3(new_n381_), .A4(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n360_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G22gat), .B(G50gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT28), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n388_), .B(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G228gat), .A2(G233gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(KEYINPUT99), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n246_), .B(new_n393_), .C1(new_n360_), .C2(new_n387_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G78gat), .B(G106gat), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n247_), .B1(new_n375_), .B2(KEYINPUT29), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n392_), .A2(KEYINPUT99), .ZN(new_n398_));
  OAI211_X1 g197(.A(new_n394_), .B(new_n396_), .C1(new_n397_), .C2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n391_), .B1(new_n400_), .B2(KEYINPUT100), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n394_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n395_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(new_n399_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n401_), .A2(new_n404_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n403_), .A2(KEYINPUT100), .A3(new_n399_), .A4(new_n391_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NOR3_X1   g206(.A1(new_n299_), .A2(new_n386_), .A3(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(KEYINPUT27), .B1(new_n297_), .B2(new_n283_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n295_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n385_), .A2(new_n379_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n411_), .A2(new_n413_), .A3(new_n407_), .A4(new_n293_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n273_), .A2(KEYINPUT32), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n289_), .A2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n417_), .B1(new_n296_), .B2(new_n416_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n418_), .B1(new_n385_), .B2(new_n379_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n370_), .A2(KEYINPUT33), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n366_), .B(new_n420_), .C1(new_n374_), .C2(new_n378_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n370_), .B1(new_n364_), .B2(new_n377_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n376_), .A2(new_n365_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n422_), .B1(new_n374_), .B2(new_n423_), .ZN(new_n424_));
  AND4_X1   g223(.A1(new_n421_), .A2(new_n424_), .A3(new_n283_), .A4(new_n297_), .ZN(new_n425_));
  XOR2_X1   g224(.A(KEYINPUT107), .B(KEYINPUT33), .Z(new_n426_));
  NAND2_X1  g225(.A1(new_n379_), .A2(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n419_), .B1(new_n425_), .B2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n414_), .B1(new_n428_), .B2(new_n407_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n323_), .A2(new_n381_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n408_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT86), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT15), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G43gat), .B(G50gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G29gat), .B(G36gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  XOR2_X1   g236(.A(G29gat), .B(G36gat), .Z(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n434_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n437_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n440_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n433_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n437_), .A2(new_n439_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n440_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(KEYINPUT15), .A3(new_n441_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n444_), .A2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G1gat), .B(G8gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT81), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G15gat), .B(G22gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G1gat), .A2(G8gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT14), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n451_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT81), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n450_), .B(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n455_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n456_), .A2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n432_), .B1(new_n449_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G229gat), .A2(G233gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n447_), .A2(new_n441_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT85), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n447_), .A2(KEYINPUT85), .A3(new_n441_), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n467_), .B(new_n468_), .C1(new_n456_), .C2(new_n460_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n449_), .A2(new_n432_), .A3(new_n461_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n463_), .A2(new_n464_), .A3(new_n469_), .A4(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n467_), .A2(new_n468_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(new_n461_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(new_n469_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n464_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n471_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G113gat), .B(G141gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G169gat), .B(G197gat), .ZN(new_n479_));
  XOR2_X1   g278(.A(new_n478_), .B(new_n479_), .Z(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n477_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n471_), .A2(new_n476_), .A3(new_n480_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n431_), .A2(new_n485_), .ZN(new_n486_));
  OAI211_X1 g285(.A(G231gat), .B(G233gat), .C1(new_n456_), .C2(new_n460_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G57gat), .B(G64gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT11), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT68), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT68), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n488_), .A2(new_n491_), .A3(KEYINPUT11), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n488_), .A2(KEYINPUT11), .ZN(new_n494_));
  XOR2_X1   g293(.A(G71gat), .B(G78gat), .Z(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n490_), .A2(new_n494_), .A3(new_n495_), .A4(new_n492_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n458_), .A2(new_n459_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n451_), .A2(new_n455_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G231gat), .A2(G233gat), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n501_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n487_), .A2(new_n500_), .A3(new_n504_), .ZN(new_n505_));
  AND3_X1   g304(.A1(new_n501_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n503_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n499_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT69), .B1(new_n505_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT82), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n505_), .A2(new_n508_), .A3(KEYINPUT69), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n512_), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT82), .B1(new_n514_), .B2(new_n509_), .ZN(new_n515_));
  XOR2_X1   g314(.A(G127gat), .B(G155gat), .Z(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT16), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G183gat), .B(G211gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT17), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n513_), .A2(new_n515_), .A3(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n519_), .B(KEYINPUT17), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n505_), .A2(new_n508_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT83), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n522_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT84), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n522_), .A2(KEYINPUT84), .A3(new_n526_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G190gat), .B(G218gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G134gat), .B(G162gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n534_), .B(KEYINPUT36), .Z(new_n535_));
  NAND2_X1  g334(.A1(G232gat), .A2(G233gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT34), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT35), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G99gat), .A2(G106gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT6), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT6), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n541_), .A2(G99gat), .A3(G106gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G85gat), .A2(G92gat), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n543_), .B1(KEYINPUT9), .B2(new_n544_), .ZN(new_n545_));
  OR2_X1    g344(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n546_));
  INV_X1    g345(.A(G106gat), .ZN(new_n547_));
  NAND2_X1  g346(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n546_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  OR2_X1    g348(.A1(G85gat), .A2(G92gat), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n550_), .A2(KEYINPUT9), .A3(new_n544_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(KEYINPUT65), .B1(new_n545_), .B2(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n544_), .A2(KEYINPUT9), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n554_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT65), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n555_), .A2(new_n556_), .A3(new_n549_), .A4(new_n551_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n553_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT8), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT67), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n541_), .B1(G99gat), .B2(G106gat), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n539_), .A2(KEYINPUT6), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n560_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n540_), .A2(new_n542_), .A3(KEYINPUT67), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n304_), .A2(new_n547_), .A3(KEYINPUT66), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(KEYINPUT7), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT7), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n567_), .A2(new_n304_), .A3(new_n547_), .A4(KEYINPUT66), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n563_), .A2(new_n564_), .A3(new_n566_), .A4(new_n568_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n550_), .A2(new_n544_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n559_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n566_), .A2(new_n543_), .A3(new_n568_), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n572_), .A2(new_n559_), .A3(new_n570_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n558_), .B1(new_n571_), .B2(new_n573_), .ZN(new_n574_));
  OAI22_X1  g373(.A1(new_n574_), .A2(new_n465_), .B1(KEYINPUT35), .B2(new_n537_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n449_), .A2(new_n574_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n575_), .B1(KEYINPUT77), .B2(new_n576_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n576_), .A2(KEYINPUT77), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n538_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n538_), .B(KEYINPUT78), .Z(new_n580_));
  NAND2_X1  g379(.A1(new_n576_), .A2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n581_), .A2(new_n575_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n535_), .B1(new_n579_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT79), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  OAI211_X1 g384(.A(KEYINPUT79), .B(new_n535_), .C1(new_n579_), .C2(new_n582_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n534_), .A2(KEYINPUT36), .ZN(new_n587_));
  OR3_X1    g386(.A1(new_n579_), .A2(new_n582_), .A3(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n585_), .A2(new_n586_), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT37), .ZN(new_n590_));
  XNOR2_X1  g389(.A(KEYINPUT80), .B(KEYINPUT37), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n588_), .A2(new_n583_), .A3(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n531_), .B1(new_n590_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT13), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n574_), .A2(new_n500_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n574_), .A2(KEYINPUT69), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(new_n597_), .A3(KEYINPUT12), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT12), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n574_), .B(new_n500_), .C1(KEYINPUT69), .C2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n499_), .B(new_n558_), .C1(new_n571_), .C2(new_n573_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G230gat), .A2(G233gat), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n603_), .B(KEYINPUT64), .Z(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n601_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT70), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n604_), .B1(new_n596_), .B2(new_n602_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n607_), .A2(new_n608_), .A3(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G176gat), .B(G204gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT72), .ZN(new_n613_));
  XNOR2_X1  g412(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G120gat), .B(G148gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n605_), .B1(new_n598_), .B2(new_n600_), .ZN(new_n618_));
  OAI21_X1  g417(.A(KEYINPUT70), .B1(new_n618_), .B2(new_n609_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n611_), .A2(new_n617_), .A3(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT74), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n609_), .B1(new_n601_), .B2(new_n606_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n617_), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT73), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT73), .ZN(new_n625_));
  NOR4_X1   g424(.A1(new_n618_), .A2(new_n625_), .A3(new_n609_), .A4(new_n617_), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n620_), .B(new_n621_), .C1(new_n624_), .C2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n607_), .A2(new_n610_), .A3(new_n623_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(new_n625_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n622_), .A2(KEYINPUT73), .A3(new_n623_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n621_), .B1(new_n632_), .B2(new_n620_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n595_), .B1(new_n628_), .B2(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n624_), .A2(new_n626_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n611_), .A2(new_n617_), .A3(new_n619_), .ZN(new_n636_));
  OAI21_X1  g435(.A(KEYINPUT74), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n637_), .A2(KEYINPUT13), .A3(new_n627_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n634_), .A2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n594_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n486_), .A2(new_n640_), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n641_), .A2(G1gat), .A3(new_n413_), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n642_), .A2(KEYINPUT38), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(KEYINPUT38), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n588_), .A2(new_n583_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n431_), .A2(new_n646_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n639_), .A2(new_n485_), .A3(new_n527_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(G1gat), .B1(new_n649_), .B2(new_n413_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n643_), .A2(new_n644_), .A3(new_n650_), .ZN(G1324gat));
  XNOR2_X1  g450(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n647_), .A2(new_n299_), .A3(new_n648_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n653_), .A2(new_n654_), .A3(G8gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n654_), .B1(new_n653_), .B2(G8gat), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n299_), .ZN(new_n658_));
  OR3_X1    g457(.A1(new_n641_), .A2(G8gat), .A3(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n652_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n659_), .B(new_n652_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n660_), .A2(new_n662_), .ZN(G1325gat));
  INV_X1    g462(.A(new_n430_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n647_), .A2(new_n664_), .A3(new_n648_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(G15gat), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n666_), .A2(KEYINPUT110), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(KEYINPUT110), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n667_), .A2(KEYINPUT41), .A3(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n641_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n670_), .A2(new_n301_), .A3(new_n664_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT41), .B1(new_n667_), .B2(new_n668_), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1326gat));
  INV_X1    g473(.A(new_n407_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G22gat), .B1(new_n649_), .B2(new_n675_), .ZN(new_n676_));
  XOR2_X1   g475(.A(new_n676_), .B(KEYINPUT42), .Z(new_n677_));
  NOR3_X1   g476(.A1(new_n641_), .A2(G22gat), .A3(new_n675_), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1327gat));
  INV_X1    g478(.A(new_n531_), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n639_), .A2(new_n680_), .A3(new_n645_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n486_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(G29gat), .B1(new_n683_), .B2(new_n412_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n590_), .A2(new_n592_), .ZN(new_n685_));
  OAI21_X1  g484(.A(KEYINPUT43), .B1(new_n431_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n687_));
  INV_X1    g486(.A(new_n685_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n298_), .A2(new_n427_), .A3(new_n421_), .A4(new_n424_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n419_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(new_n675_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n664_), .B1(new_n692_), .B2(new_n414_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n687_), .B(new_n688_), .C1(new_n693_), .C2(new_n408_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n686_), .A2(new_n694_), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n639_), .A2(new_n485_), .A3(new_n680_), .ZN(new_n696_));
  AOI21_X1  g495(.A(KEYINPUT44), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698_));
  INV_X1    g497(.A(new_n696_), .ZN(new_n699_));
  AOI211_X1 g498(.A(new_n698_), .B(new_n699_), .C1(new_n686_), .C2(new_n694_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n697_), .A2(new_n700_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n412_), .A2(G29gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n684_), .B1(new_n701_), .B2(new_n702_), .ZN(G1328gat));
  INV_X1    g502(.A(KEYINPUT46), .ZN(new_n704_));
  INV_X1    g503(.A(G36gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(new_n701_), .B2(new_n299_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n658_), .A2(G36gat), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  OR3_X1    g507(.A1(new_n682_), .A2(KEYINPUT45), .A3(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(KEYINPUT45), .B1(new_n682_), .B2(new_n708_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n704_), .B1(new_n706_), .B2(new_n712_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n697_), .A2(new_n700_), .A3(new_n658_), .ZN(new_n714_));
  OAI211_X1 g513(.A(KEYINPUT46), .B(new_n711_), .C1(new_n714_), .C2(new_n705_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1329gat));
  NAND2_X1  g515(.A1(new_n664_), .A2(G43gat), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n701_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(G43gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n720_), .B1(new_n682_), .B2(new_n430_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT47), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT47), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n719_), .A2(new_n724_), .A3(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1330gat));
  AOI21_X1  g525(.A(G50gat), .B1(new_n683_), .B2(new_n407_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n407_), .A2(G50gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n701_), .B2(new_n728_), .ZN(G1331gat));
  NAND2_X1  g528(.A1(new_n639_), .A2(new_n485_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n730_), .A2(new_n531_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n647_), .A2(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(G57gat), .B1(new_n732_), .B2(new_n413_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n431_), .A2(new_n484_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(new_n639_), .A3(new_n593_), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n413_), .A2(G57gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n733_), .B1(new_n735_), .B2(new_n736_), .ZN(G1332gat));
  OR3_X1    g536(.A1(new_n735_), .A2(G64gat), .A3(new_n658_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n732_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n299_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(KEYINPUT111), .B(KEYINPUT48), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n740_), .A2(G64gat), .A3(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n740_), .B2(G64gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n738_), .B1(new_n742_), .B2(new_n743_), .ZN(G1333gat));
  OR3_X1    g543(.A1(new_n735_), .A2(G71gat), .A3(new_n430_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G71gat), .B1(new_n732_), .B2(new_n430_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n746_), .A2(KEYINPUT49), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n746_), .A2(KEYINPUT49), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n745_), .B1(new_n747_), .B2(new_n748_), .ZN(G1334gat));
  OR3_X1    g548(.A1(new_n735_), .A2(G78gat), .A3(new_n675_), .ZN(new_n750_));
  OAI21_X1  g549(.A(G78gat), .B1(new_n732_), .B2(new_n675_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n751_), .A2(KEYINPUT50), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n751_), .A2(KEYINPUT50), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n750_), .B1(new_n752_), .B2(new_n753_), .ZN(G1335gat));
  INV_X1    g553(.A(new_n639_), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n755_), .A2(new_n680_), .A3(new_n645_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n734_), .A2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(G85gat), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n758_), .A2(new_n759_), .A3(new_n412_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n730_), .A2(new_n680_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n695_), .A2(new_n761_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n762_), .A2(new_n413_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n760_), .B1(new_n763_), .B2(new_n759_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT112), .ZN(G1336gat));
  OAI21_X1  g564(.A(G92gat), .B1(new_n762_), .B2(new_n658_), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n658_), .A2(G92gat), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n766_), .B1(new_n757_), .B2(new_n767_), .ZN(G1337gat));
  NOR2_X1   g567(.A1(new_n762_), .A2(new_n430_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n769_), .A2(new_n304_), .ZN(new_n770_));
  AND4_X1   g569(.A1(new_n664_), .A2(new_n758_), .A3(new_n546_), .A4(new_n548_), .ZN(new_n771_));
  OR3_X1    g570(.A1(new_n770_), .A2(KEYINPUT51), .A3(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT51), .B1(new_n770_), .B2(new_n771_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(G1338gat));
  NAND3_X1  g573(.A1(new_n758_), .A2(new_n547_), .A3(new_n407_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n695_), .A2(new_n407_), .A3(new_n761_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT52), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n776_), .A2(new_n777_), .A3(G106gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n776_), .B2(G106gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT53), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n782_), .B(new_n775_), .C1(new_n778_), .C2(new_n779_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n781_), .A2(new_n783_), .ZN(G1339gat));
  AOI21_X1  g583(.A(new_n480_), .B1(new_n474_), .B2(new_n464_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n470_), .A2(new_n469_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n786_), .B1(new_n787_), .B2(new_n462_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n475_), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n787_), .A2(new_n786_), .A3(new_n462_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n785_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n483_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n602_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n793_), .B1(new_n598_), .B2(new_n600_), .ZN(new_n794_));
  OAI22_X1  g593(.A1(KEYINPUT55), .A2(new_n618_), .B1(new_n794_), .B2(new_n604_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n618_), .A2(KEYINPUT55), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n617_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT56), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  OAI211_X1 g598(.A(KEYINPUT56), .B(new_n617_), .C1(new_n795_), .C2(new_n796_), .ZN(new_n800_));
  AOI211_X1 g599(.A(new_n635_), .B(new_n792_), .C1(new_n799_), .C2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n802_));
  OAI21_X1  g601(.A(KEYINPUT58), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT58), .ZN(new_n804_));
  INV_X1    g603(.A(new_n799_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n800_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n792_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n632_), .ZN(new_n809_));
  OAI211_X1 g608(.A(KEYINPUT116), .B(new_n804_), .C1(new_n807_), .C2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n803_), .A2(new_n810_), .A3(new_n688_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n812_), .A2(KEYINPUT57), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n808_), .B1(new_n628_), .B2(new_n633_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n484_), .B(new_n632_), .C1(new_n805_), .C2(new_n806_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n813_), .B1(new_n816_), .B2(new_n645_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n792_), .B1(new_n637_), .B2(new_n627_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n632_), .A2(new_n484_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n819_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n645_), .B(new_n813_), .C1(new_n818_), .C2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n811_), .B1(new_n817_), .B2(new_n822_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n593_), .A2(new_n634_), .A3(new_n485_), .A4(new_n638_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n828_), .A2(KEYINPUT113), .ZN(new_n829_));
  OR2_X1    g628(.A1(new_n824_), .A2(new_n829_), .ZN(new_n830_));
  AOI22_X1  g629(.A1(new_n823_), .A2(new_n527_), .B1(new_n827_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n658_), .A2(new_n675_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n664_), .A2(new_n412_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n831_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT59), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n645_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n839_), .B1(new_n812_), .B2(KEYINPUT57), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n821_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n680_), .B1(new_n841_), .B2(new_n811_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n824_), .A2(new_n829_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n843_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n842_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n834_), .A2(new_n837_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n838_), .A2(new_n847_), .A3(new_n485_), .ZN(new_n848_));
  INV_X1    g647(.A(G113gat), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT117), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n850_), .B1(new_n831_), .B2(new_n835_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n527_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(new_n841_), .B2(new_n811_), .ZN(new_n853_));
  OAI211_X1 g652(.A(KEYINPUT117), .B(new_n834_), .C1(new_n853_), .C2(new_n844_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n851_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n484_), .A2(new_n849_), .ZN(new_n856_));
  OAI22_X1  g655(.A1(new_n848_), .A2(new_n849_), .B1(new_n855_), .B2(new_n856_), .ZN(G1340gat));
  XNOR2_X1  g656(.A(KEYINPUT118), .B(G120gat), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n639_), .A2(new_n858_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n851_), .B(new_n854_), .C1(KEYINPUT60), .C2(new_n859_), .ZN(new_n860_));
  OR2_X1    g659(.A1(new_n860_), .A2(KEYINPUT60), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n838_), .A2(new_n847_), .A3(new_n755_), .ZN(new_n862_));
  AOI22_X1  g661(.A1(new_n861_), .A2(new_n858_), .B1(new_n862_), .B2(new_n860_), .ZN(G1341gat));
  NOR2_X1   g662(.A1(new_n838_), .A2(new_n847_), .ZN(new_n864_));
  XOR2_X1   g663(.A(KEYINPUT119), .B(G127gat), .Z(new_n865_));
  NAND2_X1  g664(.A1(new_n852_), .A2(new_n865_), .ZN(new_n866_));
  XOR2_X1   g665(.A(new_n866_), .B(KEYINPUT120), .Z(new_n867_));
  INV_X1    g666(.A(G127gat), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n851_), .A2(new_n680_), .A3(new_n854_), .ZN(new_n869_));
  AOI22_X1  g668(.A1(new_n864_), .A2(new_n867_), .B1(new_n868_), .B2(new_n869_), .ZN(G1342gat));
  NAND3_X1  g669(.A1(new_n851_), .A2(new_n646_), .A3(new_n854_), .ZN(new_n871_));
  INV_X1    g670(.A(G134gat), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  XOR2_X1   g672(.A(KEYINPUT121), .B(G134gat), .Z(new_n874_));
  NOR2_X1   g673(.A1(new_n685_), .A2(new_n874_), .ZN(new_n875_));
  OAI221_X1 g674(.A(new_n875_), .B1(new_n845_), .B2(new_n846_), .C1(new_n836_), .C2(new_n837_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n873_), .A2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT122), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n873_), .A2(KEYINPUT122), .A3(new_n876_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1343gat));
  INV_X1    g680(.A(new_n831_), .ZN(new_n882_));
  NOR4_X1   g681(.A1(new_n664_), .A2(new_n299_), .A3(new_n675_), .A4(new_n413_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n485_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(new_n344_), .ZN(G1344gat));
  NOR2_X1   g685(.A1(new_n884_), .A2(new_n755_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(new_n345_), .ZN(G1345gat));
  NOR2_X1   g687(.A1(new_n884_), .A2(new_n531_), .ZN(new_n889_));
  XOR2_X1   g688(.A(KEYINPUT61), .B(G155gat), .Z(new_n890_));
  XNOR2_X1  g689(.A(new_n889_), .B(new_n890_), .ZN(G1346gat));
  INV_X1    g690(.A(G162gat), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n884_), .A2(new_n892_), .A3(new_n685_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n884_), .B2(new_n645_), .ZN(new_n894_));
  OR2_X1    g693(.A1(new_n894_), .A2(KEYINPUT123), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(KEYINPUT123), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n893_), .B1(new_n895_), .B2(new_n896_), .ZN(G1347gat));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n658_), .A2(new_n386_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n845_), .A2(new_n407_), .A3(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n484_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n898_), .B1(new_n902_), .B2(G169gat), .ZN(new_n903_));
  AOI211_X1 g702(.A(KEYINPUT62), .B(new_n251_), .C1(new_n901_), .C2(new_n484_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n901_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n484_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n906_));
  XOR2_X1   g705(.A(new_n906_), .B(KEYINPUT124), .Z(new_n907_));
  OAI22_X1  g706(.A1(new_n903_), .A2(new_n904_), .B1(new_n905_), .B2(new_n907_), .ZN(G1348gat));
  OAI21_X1  g707(.A(new_n675_), .B1(new_n853_), .B2(new_n844_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT125), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n900_), .B1(new_n909_), .B2(new_n910_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n882_), .A2(KEYINPUT125), .A3(new_n675_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n755_), .A2(new_n250_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n911_), .A2(new_n912_), .A3(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT126), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n250_), .B1(new_n905_), .B2(new_n755_), .ZN(new_n917_));
  NAND4_X1  g716(.A1(new_n911_), .A2(KEYINPUT126), .A3(new_n912_), .A4(new_n913_), .ZN(new_n918_));
  AND3_X1   g717(.A1(new_n916_), .A2(new_n917_), .A3(new_n918_), .ZN(G1349gat));
  NOR3_X1   g718(.A1(new_n905_), .A2(new_n211_), .A3(new_n527_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n911_), .A2(new_n680_), .A3(new_n912_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n920_), .B1(new_n216_), .B2(new_n921_), .ZN(G1350gat));
  OAI21_X1  g721(.A(G190gat), .B1(new_n905_), .B2(new_n685_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n901_), .A2(new_n212_), .A3(new_n646_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1351gat));
  NOR4_X1   g724(.A1(new_n658_), .A2(new_n664_), .A3(new_n412_), .A4(new_n675_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n882_), .A2(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(new_n484_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g729(.A1(new_n928_), .A2(new_n639_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g731(.A(KEYINPUT63), .B(G211gat), .C1(new_n928_), .C2(new_n852_), .ZN(new_n933_));
  XOR2_X1   g732(.A(KEYINPUT63), .B(G211gat), .Z(new_n934_));
  NAND4_X1  g733(.A1(new_n882_), .A2(new_n852_), .A3(new_n926_), .A4(new_n934_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n935_), .A2(KEYINPUT127), .ZN(new_n936_));
  AND2_X1   g735(.A1(new_n935_), .A2(KEYINPUT127), .ZN(new_n937_));
  NOR3_X1   g736(.A1(new_n933_), .A2(new_n936_), .A3(new_n937_), .ZN(G1354gat));
  OAI21_X1  g737(.A(G218gat), .B1(new_n927_), .B2(new_n685_), .ZN(new_n939_));
  OR2_X1    g738(.A1(new_n645_), .A2(G218gat), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n939_), .B1(new_n927_), .B2(new_n940_), .ZN(G1355gat));
endmodule


