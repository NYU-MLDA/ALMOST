//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 1 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n912_;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G169gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(KEYINPUT80), .A2(G176gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(KEYINPUT80), .A2(G176gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n202_), .A2(new_n203_), .A3(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT81), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n208_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n212_));
  AOI22_X1  g011(.A1(new_n211_), .A2(new_n212_), .B1(G169gat), .B2(G176gat), .ZN(new_n213_));
  AND2_X1   g012(.A1(new_n203_), .A2(new_n204_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(KEYINPUT81), .A3(new_n202_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n207_), .A2(new_n213_), .A3(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G183gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT25), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT25), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(G183gat), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G190gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT26), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT26), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(G190gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n221_), .A2(new_n223_), .A3(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n210_), .B(new_n209_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(G169gat), .ZN(new_n229_));
  INV_X1    g028(.A(G176gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G169gat), .A2(G176gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(KEYINPUT24), .A3(new_n232_), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n231_), .A2(KEYINPUT24), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n226_), .A2(new_n228_), .A3(new_n233_), .A4(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n216_), .A2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G71gat), .B(G99gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(G43gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n236_), .B(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G227gat), .A2(G233gat), .ZN(new_n240_));
  INV_X1    g039(.A(G15gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT30), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n239_), .A2(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n239_), .A2(new_n243_), .ZN(new_n245_));
  OR3_X1    g044(.A1(new_n244_), .A2(new_n245_), .A3(KEYINPUT83), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(KEYINPUT84), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT83), .B1(new_n244_), .B2(new_n245_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G127gat), .B(G134gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G113gat), .B(G120gat), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT82), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n249_), .A2(new_n250_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n249_), .A2(new_n250_), .A3(KEYINPUT82), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT31), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n248_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n247_), .A2(new_n259_), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n246_), .A2(KEYINPUT84), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n246_), .A2(KEYINPUT84), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n261_), .A2(new_n248_), .A3(new_n258_), .A4(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n260_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT102), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT20), .ZN(new_n266_));
  INV_X1    g065(.A(G204gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(G197gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT88), .ZN(new_n269_));
  INV_X1    g068(.A(G197gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(G204gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n268_), .A2(KEYINPUT88), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT21), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT90), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n271_), .A2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n270_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n268_), .A2(KEYINPUT89), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT21), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n268_), .A2(KEYINPUT89), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n278_), .A2(new_n279_), .A3(new_n280_), .A4(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G211gat), .B(G218gat), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n274_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n278_), .A2(new_n281_), .A3(new_n279_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n283_), .A2(new_n280_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n284_), .A2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n266_), .B1(new_n288_), .B2(new_n236_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT94), .B(KEYINPUT24), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n291_), .A2(new_n231_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n292_), .A2(new_n227_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n224_), .A2(G190gat), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n222_), .A2(KEYINPUT26), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT93), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT93), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n223_), .A2(new_n225_), .A3(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(new_n221_), .A3(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n291_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n299_), .A2(KEYINPUT95), .A3(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(KEYINPUT95), .B1(new_n299_), .B2(new_n300_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n293_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n213_), .A2(new_n205_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT101), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n288_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n303_), .A2(KEYINPUT101), .A3(new_n304_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n290_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G226gat), .A2(G233gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT19), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n265_), .B1(new_n309_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n293_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT95), .ZN(new_n315_));
  AND3_X1   g114(.A1(new_n223_), .A2(new_n225_), .A3(new_n297_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n297_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n218_), .A2(new_n220_), .ZN(new_n318_));
  NOR3_X1   g117(.A1(new_n316_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n300_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n315_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n299_), .A2(KEYINPUT95), .A3(new_n300_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n314_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n304_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n306_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  AND2_X1   g124(.A1(new_n284_), .A2(new_n287_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n325_), .A2(new_n326_), .A3(new_n308_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(new_n289_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n328_), .A2(KEYINPUT102), .A3(new_n311_), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT20), .B1(new_n288_), .B2(new_n236_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n330_), .B1(new_n305_), .B2(new_n288_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n311_), .B(KEYINPUT92), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n313_), .A2(new_n329_), .A3(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(G8gat), .B(G36gat), .Z(new_n335_));
  XNOR2_X1  g134(.A(G64gat), .B(G92gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT32), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n334_), .A2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(G155gat), .A2(G162gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT85), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G155gat), .A2(G162gat), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT86), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G141gat), .A2(G148gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT2), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n352_));
  NOR2_X1   g151(.A1(G141gat), .A2(G148gat), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n351_), .B(new_n352_), .C1(new_n354_), .C2(KEYINPUT3), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n345_), .B(new_n346_), .C1(new_n348_), .C2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n343_), .B(KEYINPUT85), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n346_), .B(KEYINPUT1), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n354_), .B(new_n349_), .C1(new_n357_), .C2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n356_), .A2(new_n359_), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n257_), .A2(new_n360_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n252_), .A2(new_n254_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT4), .B1(new_n361_), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G225gat), .A2(G233gat), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n257_), .A2(new_n360_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT4), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n364_), .A2(new_n366_), .A3(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n367_), .B1(new_n360_), .B2(new_n362_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n365_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  XOR2_X1   g172(.A(G1gat), .B(G29gat), .Z(new_n374_));
  XNOR2_X1  g173(.A(G57gat), .B(G85gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT98), .B(KEYINPUT0), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n373_), .A2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n370_), .A2(new_n378_), .A3(new_n372_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n312_), .B(new_n289_), .C1(new_n305_), .C2(new_n288_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n383_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n384_));
  OR3_X1    g183(.A1(new_n384_), .A2(KEYINPUT100), .A3(new_n341_), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT100), .B1(new_n384_), .B2(new_n341_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n342_), .A2(new_n382_), .A3(new_n385_), .A4(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n339_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n303_), .A2(new_n326_), .A3(new_n304_), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n389_), .A2(new_n312_), .A3(new_n289_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n288_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n236_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n266_), .B1(new_n326_), .B2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n332_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n388_), .B1(new_n390_), .B2(new_n394_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n383_), .B(new_n339_), .C1(new_n331_), .C2(new_n332_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n395_), .A2(KEYINPUT97), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT97), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n384_), .A2(new_n398_), .A3(new_n388_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n366_), .B1(new_n364_), .B2(new_n369_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n378_), .B1(new_n371_), .B2(new_n365_), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT99), .ZN(new_n404_));
  AOI21_X1  g203(.A(KEYINPUT33), .B1(new_n380_), .B2(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n378_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT33), .ZN(new_n407_));
  NOR3_X1   g206(.A1(new_n406_), .A2(KEYINPUT99), .A3(new_n407_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n400_), .B(new_n403_), .C1(new_n405_), .C2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n387_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT91), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n326_), .B1(KEYINPUT29), .B2(new_n360_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n415_));
  OAI21_X1  g214(.A(G228gat), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  OR2_X1    g215(.A1(new_n412_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n412_), .A2(new_n416_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G78gat), .B(G106gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n420_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n417_), .A2(new_n418_), .A3(new_n422_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n360_), .A2(KEYINPUT29), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G22gat), .B(G50gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT28), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n424_), .B(new_n426_), .ZN(new_n427_));
  AND4_X1   g226(.A1(new_n411_), .A2(new_n421_), .A3(new_n423_), .A4(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n423_), .A2(KEYINPUT91), .ZN(new_n429_));
  AOI22_X1  g228(.A1(new_n429_), .A2(new_n427_), .B1(new_n421_), .B2(new_n423_), .ZN(new_n430_));
  OR2_X1    g229(.A1(new_n428_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n410_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n396_), .A2(KEYINPUT27), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n433_), .B1(new_n334_), .B2(new_n388_), .ZN(new_n434_));
  XOR2_X1   g233(.A(KEYINPUT103), .B(KEYINPUT27), .Z(new_n435_));
  AND3_X1   g234(.A1(new_n397_), .A2(new_n399_), .A3(new_n435_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n382_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n428_), .A2(new_n430_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n437_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n264_), .B1(new_n432_), .B2(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT104), .B1(new_n434_), .B2(new_n436_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT104), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n397_), .A2(new_n399_), .A3(new_n435_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n333_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n328_), .A2(new_n311_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n445_), .B1(new_n446_), .B2(new_n265_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n339_), .B1(new_n447_), .B2(new_n329_), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n443_), .B(new_n444_), .C1(new_n448_), .C2(new_n433_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n442_), .A2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n382_), .B1(new_n260_), .B2(new_n263_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n450_), .A2(new_n431_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT105), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n439_), .B1(new_n442_), .B2(new_n449_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n455_), .A2(KEYINPUT105), .A3(new_n451_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n441_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G1gat), .B(G8gat), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n458_), .A2(KEYINPUT71), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(KEYINPUT71), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G15gat), .B(G22gat), .ZN(new_n462_));
  INV_X1    g261(.A(G1gat), .ZN(new_n463_));
  INV_X1    g262(.A(G8gat), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT14), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n462_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n461_), .A2(new_n466_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n459_), .A2(new_n465_), .A3(new_n462_), .A4(new_n460_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G29gat), .B(G36gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G43gat), .B(G50gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n469_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n467_), .A2(new_n472_), .A3(new_n468_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT77), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G229gat), .A2(G233gat), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n474_), .A2(KEYINPUT77), .A3(new_n475_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n478_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(KEYINPUT68), .B(KEYINPUT15), .Z(new_n483_));
  XNOR2_X1  g282(.A(new_n472_), .B(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n469_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n485_), .A2(new_n479_), .A3(new_n475_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT78), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT78), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n485_), .A2(new_n488_), .A3(new_n479_), .A4(new_n475_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n482_), .A2(new_n487_), .A3(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT79), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G113gat), .B(G141gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G169gat), .B(G197gat), .ZN(new_n493_));
  XOR2_X1   g292(.A(new_n492_), .B(new_n493_), .Z(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n491_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n490_), .A2(KEYINPUT79), .A3(new_n494_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT106), .B1(new_n457_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n264_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n440_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n439_), .B1(new_n387_), .B2(new_n409_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n500_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  AND4_X1   g302(.A1(KEYINPUT105), .A2(new_n450_), .A3(new_n431_), .A4(new_n451_), .ZN(new_n504_));
  AOI21_X1  g303(.A(KEYINPUT105), .B1(new_n455_), .B2(new_n451_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n503_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT106), .ZN(new_n507_));
  INV_X1    g306(.A(new_n498_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n506_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n499_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G99gat), .A2(G106gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT6), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT9), .ZN(new_n513_));
  INV_X1    g312(.A(G85gat), .ZN(new_n514_));
  INV_X1    g313(.A(G92gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G85gat), .A2(G92gat), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT65), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n513_), .B(new_n516_), .C1(new_n518_), .C2(new_n519_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n516_), .A2(KEYINPUT65), .A3(KEYINPUT9), .A4(new_n517_), .ZN(new_n521_));
  OR2_X1    g320(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n522_));
  INV_X1    g321(.A(G106gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n522_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n512_), .A2(new_n520_), .A3(new_n521_), .A4(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n516_), .A2(new_n517_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT6), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n511_), .B(new_n529_), .ZN(new_n530_));
  OR3_X1    g329(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n528_), .B1(new_n530_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT8), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT8), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n536_), .B(new_n528_), .C1(new_n530_), .C2(new_n533_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n527_), .B1(new_n535_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(new_n484_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT69), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G232gat), .A2(G233gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT34), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n541_), .A2(KEYINPUT35), .A3(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n538_), .A2(new_n472_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n540_), .A2(new_n545_), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n540_), .B(new_n545_), .C1(KEYINPUT35), .C2(new_n543_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n544_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G190gat), .B(G218gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G134gat), .B(G162gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n553_), .A2(KEYINPUT36), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n550_), .A2(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n553_), .B(KEYINPUT36), .Z(new_n556_));
  NAND3_X1  g355(.A1(new_n547_), .A2(new_n549_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT37), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT70), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n559_), .B1(new_n557_), .B2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n558_), .B(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(G183gat), .B(G211gat), .Z(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT73), .ZN(new_n564_));
  XNOR2_X1  g363(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT74), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n564_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G127gat), .B(G155gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT17), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G231gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n469_), .B(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(G64gat), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(G57gat), .ZN(new_n575_));
  INV_X1    g374(.A(G57gat), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(G64gat), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n575_), .A2(new_n577_), .A3(KEYINPUT11), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(KEYINPUT66), .B(G71gat), .ZN(new_n580_));
  INV_X1    g379(.A(G78gat), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n580_), .A2(new_n581_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n579_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(KEYINPUT66), .B(G71gat), .Z(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(G78gat), .ZN(new_n587_));
  AOI21_X1  g386(.A(KEYINPUT11), .B1(new_n575_), .B2(new_n577_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n587_), .B(new_n582_), .C1(new_n588_), .C2(new_n578_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n585_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n573_), .B(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n571_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT75), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n592_), .B1(new_n570_), .B2(new_n569_), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n594_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n595_), .B1(new_n594_), .B2(new_n596_), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n562_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT67), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n601_), .B1(new_n538_), .B2(new_n590_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT12), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G230gat), .A2(G233gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT64), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n538_), .A2(new_n590_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT12), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n601_), .B(new_n608_), .C1(new_n538_), .C2(new_n590_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n603_), .A2(new_n606_), .A3(new_n607_), .A4(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n607_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n538_), .A2(new_n590_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n605_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n610_), .A2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G120gat), .B(G148gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT5), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G176gat), .B(G204gat), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n616_), .B(new_n617_), .Z(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n614_), .B(new_n619_), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n620_), .A2(KEYINPUT13), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(KEYINPUT13), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n600_), .A2(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n624_), .B(KEYINPUT76), .Z(new_n625_));
  NOR2_X1   g424(.A1(new_n510_), .A2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n626_), .A2(new_n463_), .A3(new_n382_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT38), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n627_), .A2(new_n628_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n623_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n631_), .A2(new_n599_), .A3(new_n508_), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n632_), .B(KEYINPUT107), .Z(new_n633_));
  INV_X1    g432(.A(KEYINPUT109), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT108), .ZN(new_n635_));
  INV_X1    g434(.A(new_n557_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n554_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n637_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n635_), .B1(new_n636_), .B2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n555_), .A2(KEYINPUT108), .A3(new_n557_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n634_), .B1(new_n506_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n506_), .A2(new_n634_), .A3(new_n641_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n633_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n463_), .B1(new_n645_), .B2(new_n382_), .ZN(new_n646_));
  OR3_X1    g445(.A1(new_n629_), .A2(new_n630_), .A3(new_n646_), .ZN(G1324gat));
  INV_X1    g446(.A(new_n450_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n626_), .A2(new_n464_), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n633_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n644_), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n648_), .B(new_n650_), .C1(new_n651_), .C2(new_n642_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT39), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n652_), .A2(new_n653_), .A3(G8gat), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n653_), .B1(new_n652_), .B2(G8gat), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n649_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT40), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n649_), .B(KEYINPUT40), .C1(new_n654_), .C2(new_n655_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1325gat));
  NAND3_X1  g459(.A1(new_n626_), .A2(new_n241_), .A3(new_n264_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n645_), .A2(new_n264_), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n662_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(KEYINPUT41), .B1(new_n662_), .B2(G15gat), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n661_), .B1(new_n663_), .B2(new_n664_), .ZN(G1326gat));
  INV_X1    g464(.A(G22gat), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n626_), .A2(new_n666_), .A3(new_n439_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n645_), .ZN(new_n668_));
  OAI21_X1  g467(.A(G22gat), .B1(new_n668_), .B2(new_n431_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n669_), .A2(KEYINPUT42), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(KEYINPUT42), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n667_), .B1(new_n670_), .B2(new_n671_), .ZN(G1327gat));
  NOR2_X1   g471(.A1(new_n641_), .A2(new_n599_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(new_n631_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n674_), .B1(new_n499_), .B2(new_n509_), .ZN(new_n675_));
  AOI21_X1  g474(.A(G29gat), .B1(new_n675_), .B2(new_n382_), .ZN(new_n676_));
  OAI21_X1  g475(.A(KEYINPUT43), .B1(new_n562_), .B2(KEYINPUT111), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n678_), .B1(new_n457_), .B2(new_n562_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n558_), .B(new_n561_), .Z(new_n680_));
  NAND3_X1  g479(.A1(new_n506_), .A2(new_n680_), .A3(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n599_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n631_), .A2(new_n683_), .A3(new_n508_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT110), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(KEYINPUT44), .B1(new_n682_), .B2(new_n686_), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n457_), .A2(new_n562_), .A3(new_n678_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n677_), .B1(new_n506_), .B2(new_n680_), .ZN(new_n689_));
  OAI211_X1 g488(.A(KEYINPUT44), .B(new_n686_), .C1(new_n688_), .C2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT112), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n685_), .B1(new_n679_), .B2(new_n681_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT112), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n692_), .A2(new_n693_), .A3(KEYINPUT44), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n687_), .B1(new_n691_), .B2(new_n694_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n382_), .A2(G29gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n676_), .B1(new_n695_), .B2(new_n696_), .ZN(G1328gat));
  INV_X1    g496(.A(KEYINPUT46), .ZN(new_n698_));
  INV_X1    g497(.A(G36gat), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n691_), .A2(new_n694_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n648_), .B1(new_n692_), .B2(KEYINPUT44), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n699_), .B1(new_n700_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT45), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n450_), .A2(G36gat), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n675_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n704_), .B1(new_n675_), .B2(new_n705_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n698_), .B1(new_n703_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n708_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n706_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n701_), .B1(new_n691_), .B2(new_n694_), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n712_), .B(KEYINPUT46), .C1(new_n713_), .C2(new_n699_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n710_), .A2(new_n714_), .ZN(G1329gat));
  NAND2_X1  g514(.A1(new_n264_), .A2(G43gat), .ZN(new_n716_));
  AOI211_X1 g515(.A(new_n716_), .B(new_n687_), .C1(new_n691_), .C2(new_n694_), .ZN(new_n717_));
  AOI21_X1  g516(.A(G43gat), .B1(new_n675_), .B2(new_n264_), .ZN(new_n718_));
  OAI21_X1  g517(.A(KEYINPUT47), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n716_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n695_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n718_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT47), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n721_), .A2(new_n722_), .A3(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n719_), .A2(new_n724_), .ZN(G1330gat));
  AOI21_X1  g524(.A(G50gat), .B1(new_n675_), .B2(new_n439_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n439_), .A2(G50gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n695_), .B2(new_n727_), .ZN(G1331gat));
  NOR4_X1   g527(.A1(new_n457_), .A2(new_n508_), .A3(new_n631_), .A4(new_n600_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n729_), .A2(new_n576_), .A3(new_n382_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n623_), .A2(new_n599_), .A3(new_n498_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n732_), .A2(new_n382_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n730_), .B1(new_n733_), .B2(new_n576_), .ZN(G1332gat));
  NAND3_X1  g533(.A1(new_n729_), .A2(new_n574_), .A3(new_n648_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n574_), .B1(new_n732_), .B2(new_n648_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT48), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n736_), .A2(new_n737_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n738_), .B2(new_n739_), .ZN(G1333gat));
  INV_X1    g539(.A(G71gat), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n729_), .A2(new_n741_), .A3(new_n264_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n732_), .B2(new_n264_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(KEYINPUT113), .B(KEYINPUT49), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n743_), .A2(new_n744_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n742_), .B1(new_n745_), .B2(new_n746_), .ZN(G1334gat));
  NAND3_X1  g546(.A1(new_n729_), .A2(new_n581_), .A3(new_n439_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n581_), .B1(new_n732_), .B2(new_n439_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT50), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n749_), .A2(new_n750_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(G1335gat));
  NAND3_X1  g552(.A1(new_n683_), .A2(new_n498_), .A3(new_n623_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n754_), .B1(new_n679_), .B2(new_n681_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n755_), .A2(G85gat), .A3(new_n382_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT114), .ZN(new_n757_));
  AND4_X1   g556(.A1(new_n506_), .A2(new_n498_), .A3(new_n623_), .A4(new_n673_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n382_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n757_), .B1(new_n759_), .B2(new_n514_), .ZN(new_n760_));
  AOI211_X1 g559(.A(KEYINPUT114), .B(G85gat), .C1(new_n758_), .C2(new_n382_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n756_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT115), .ZN(G1336gat));
  NAND3_X1  g562(.A1(new_n758_), .A2(new_n515_), .A3(new_n648_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n755_), .A2(new_n648_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(new_n515_), .ZN(G1337gat));
  NAND4_X1  g565(.A1(new_n758_), .A2(new_n264_), .A3(new_n522_), .A4(new_n524_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT116), .ZN(new_n768_));
  INV_X1    g567(.A(G99gat), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n755_), .A2(new_n264_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n768_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n772_), .A2(KEYINPUT117), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n771_), .A2(new_n773_), .ZN(new_n774_));
  OAI221_X1 g573(.A(new_n768_), .B1(KEYINPUT117), .B2(new_n772_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1338gat));
  NAND3_X1  g575(.A1(new_n758_), .A2(new_n523_), .A3(new_n439_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n755_), .A2(new_n439_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n779_), .B2(G106gat), .ZN(new_n780_));
  AOI211_X1 g579(.A(KEYINPUT52), .B(new_n523_), .C1(new_n755_), .C2(new_n439_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n777_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT53), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT53), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n784_), .B(new_n777_), .C1(new_n780_), .C2(new_n781_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(G1339gat));
  NAND4_X1  g585(.A1(new_n562_), .A2(new_n631_), .A3(new_n599_), .A4(new_n498_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT54), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n787_), .B(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n610_), .A2(new_n613_), .A3(new_n619_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n496_), .A2(new_n497_), .A3(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT56), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT118), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n610_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(new_n610_), .B2(new_n793_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n611_), .B1(KEYINPUT12), .B2(new_n602_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n606_), .B1(new_n797_), .B2(new_n609_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n795_), .A2(new_n796_), .A3(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n792_), .B1(new_n799_), .B2(new_n619_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n610_), .A2(new_n793_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT55), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n610_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n798_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n802_), .A2(new_n803_), .A3(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(KEYINPUT56), .A3(new_n618_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n791_), .B1(new_n800_), .B2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n480_), .B1(new_n478_), .B2(new_n481_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n479_), .B1(new_n485_), .B2(new_n475_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n495_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n482_), .A2(new_n487_), .A3(new_n489_), .A4(new_n494_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n620_), .A2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n641_), .B1(new_n807_), .B2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n641_), .B(KEYINPUT57), .C1(new_n813_), .C2(new_n807_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT119), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n800_), .A2(new_n818_), .A3(new_n806_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n810_), .A2(new_n790_), .A3(new_n811_), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT56), .B1(new_n805_), .B2(new_n618_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n820_), .B1(new_n821_), .B2(KEYINPUT119), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT120), .B1(new_n819_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT58), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n680_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  AOI211_X1 g624(.A(KEYINPUT120), .B(KEYINPUT58), .C1(new_n819_), .C2(new_n822_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n816_), .B(new_n817_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n789_), .B1(new_n683_), .B2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n455_), .A2(new_n382_), .A3(new_n264_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(G113gat), .B1(new_n830_), .B2(new_n508_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT121), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n831_), .B(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(KEYINPUT59), .B1(new_n828_), .B2(new_n829_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n827_), .A2(new_n683_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT122), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n827_), .A2(KEYINPUT122), .A3(new_n683_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n789_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  OR2_X1    g638(.A1(new_n829_), .A2(KEYINPUT59), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n834_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT123), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n834_), .B(KEYINPUT123), .C1(new_n839_), .C2(new_n840_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n508_), .A2(G113gat), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n833_), .B1(new_n845_), .B2(new_n846_), .ZN(G1340gat));
  OAI21_X1  g646(.A(G120gat), .B1(new_n841_), .B2(new_n631_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT60), .ZN(new_n849_));
  AOI21_X1  g648(.A(G120gat), .B1(new_n623_), .B2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(KEYINPUT124), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT124), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(new_n849_), .B2(G120gat), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n830_), .B(new_n851_), .C1(new_n850_), .C2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n848_), .A2(new_n854_), .ZN(G1341gat));
  AOI21_X1  g654(.A(G127gat), .B1(new_n830_), .B2(new_n599_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n683_), .A2(KEYINPUT125), .ZN(new_n857_));
  MUX2_X1   g656(.A(KEYINPUT125), .B(new_n857_), .S(G127gat), .Z(new_n858_));
  AOI21_X1  g657(.A(new_n856_), .B1(new_n845_), .B2(new_n858_), .ZN(G1342gat));
  NAND3_X1  g658(.A1(new_n843_), .A2(new_n680_), .A3(new_n844_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(G134gat), .ZN(new_n861_));
  INV_X1    g660(.A(G134gat), .ZN(new_n862_));
  INV_X1    g661(.A(new_n641_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n830_), .A2(new_n862_), .A3(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n861_), .A2(new_n864_), .ZN(G1343gat));
  NOR2_X1   g664(.A1(new_n828_), .A2(new_n264_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n866_), .A2(new_n382_), .A3(new_n439_), .A4(new_n450_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n867_), .A2(new_n498_), .ZN(new_n868_));
  XOR2_X1   g667(.A(new_n868_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g668(.A1(new_n867_), .A2(new_n631_), .ZN(new_n870_));
  XOR2_X1   g669(.A(new_n870_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g670(.A1(new_n867_), .A2(new_n683_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT61), .B(G155gat), .ZN(new_n873_));
  XOR2_X1   g672(.A(new_n872_), .B(new_n873_), .Z(G1346gat));
  OAI21_X1  g673(.A(G162gat), .B1(new_n867_), .B2(new_n562_), .ZN(new_n875_));
  OR2_X1    g674(.A1(new_n641_), .A2(G162gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n867_), .B2(new_n876_), .ZN(G1347gat));
  NAND3_X1  g676(.A1(new_n648_), .A2(new_n431_), .A3(new_n451_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n839_), .A2(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n229_), .B1(new_n879_), .B2(new_n508_), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n880_), .A2(KEYINPUT62), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n879_), .A2(new_n202_), .A3(new_n508_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(KEYINPUT62), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n881_), .A2(new_n882_), .A3(new_n883_), .ZN(G1348gat));
  NAND2_X1  g683(.A1(new_n879_), .A2(new_n623_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n828_), .A2(new_n439_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n648_), .A2(new_n451_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n887_), .A2(new_n230_), .A3(new_n631_), .ZN(new_n888_));
  AOI22_X1  g687(.A1(new_n885_), .A2(new_n214_), .B1(new_n886_), .B2(new_n888_), .ZN(G1349gat));
  NOR2_X1   g688(.A1(new_n887_), .A2(new_n683_), .ZN(new_n890_));
  AOI21_X1  g689(.A(G183gat), .B1(new_n886_), .B2(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n683_), .A2(new_n221_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n879_), .B2(new_n892_), .ZN(G1350gat));
  NAND4_X1  g692(.A1(new_n879_), .A2(new_n296_), .A3(new_n298_), .A4(new_n863_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n839_), .A2(new_n562_), .A3(new_n878_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n222_), .B2(new_n895_), .ZN(G1351gat));
  NOR3_X1   g695(.A1(new_n450_), .A2(new_n382_), .A3(new_n431_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n866_), .A2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n498_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(new_n270_), .ZN(G1352gat));
  INV_X1    g699(.A(new_n898_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n623_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(KEYINPUT126), .B(G204gat), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n902_), .B(new_n903_), .ZN(G1353gat));
  AOI21_X1  g703(.A(new_n683_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n901_), .A2(new_n905_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n907_));
  XOR2_X1   g706(.A(new_n906_), .B(new_n907_), .Z(G1354gat));
  AND3_X1   g707(.A1(new_n901_), .A2(G218gat), .A3(new_n680_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n898_), .A2(new_n641_), .ZN(new_n910_));
  OR2_X1    g709(.A1(new_n910_), .A2(KEYINPUT127), .ZN(new_n911_));
  AOI21_X1  g710(.A(G218gat), .B1(new_n910_), .B2(KEYINPUT127), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n909_), .B1(new_n911_), .B2(new_n912_), .ZN(G1355gat));
endmodule


