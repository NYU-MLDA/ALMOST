//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 1 1 1 0 0 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n785_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n921_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n960_,
    new_n961_, new_n962_, new_n964_, new_n966_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n973_, new_n974_, new_n975_;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203_));
  INV_X1    g002(.A(G1gat), .ZN(new_n204_));
  INV_X1    g003(.A(G8gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n203_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G1gat), .B(G8gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G57gat), .B(G64gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT11), .ZN(new_n211_));
  XOR2_X1   g010(.A(G71gat), .B(G78gat), .Z(new_n212_));
  OR2_X1    g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n210_), .A2(KEYINPUT11), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(new_n212_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n213_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G231gat), .ZN(new_n217_));
  INV_X1    g016(.A(G233gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n216_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT69), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n213_), .B(new_n219_), .C1(new_n214_), .C2(new_n215_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n222_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n209_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n226_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n209_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(new_n229_), .A3(new_n224_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n227_), .A2(new_n230_), .A3(KEYINPUT70), .ZN(new_n231_));
  XOR2_X1   g030(.A(G127gat), .B(G155gat), .Z(new_n232_));
  XNOR2_X1  g031(.A(G183gat), .B(G211gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT71), .B(KEYINPUT16), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT17), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n231_), .A2(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(KEYINPUT70), .B1(new_n227_), .B2(new_n230_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n202_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n240_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n242_), .A2(KEYINPUT72), .A3(new_n238_), .A4(new_n231_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n236_), .B(KEYINPUT17), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n230_), .A2(new_n227_), .A3(new_n245_), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n244_), .A2(new_n246_), .A3(KEYINPUT73), .ZN(new_n247_));
  AOI21_X1  g046(.A(KEYINPUT73), .B1(new_n244_), .B2(new_n246_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT68), .B(KEYINPUT37), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G232gat), .A2(G233gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT67), .ZN(new_n254_));
  XOR2_X1   g053(.A(KEYINPUT66), .B(KEYINPUT34), .Z(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G29gat), .B(G36gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G43gat), .B(G50gat), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n258_), .B(new_n259_), .Z(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT15), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n258_), .B(new_n259_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT15), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  XOR2_X1   g063(.A(KEYINPUT10), .B(G99gat), .Z(new_n265_));
  INV_X1    g064(.A(G106gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  XOR2_X1   g066(.A(G85gat), .B(G92gat), .Z(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT9), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G99gat), .A2(G106gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT6), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT9), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n272_), .A2(G85gat), .A3(G92gat), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n267_), .A2(new_n269_), .A3(new_n271_), .A4(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n268_), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n276_));
  AND2_X1   g075(.A1(new_n271_), .A2(new_n276_), .ZN(new_n277_));
  NOR3_X1   g076(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT64), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n275_), .B1(new_n277_), .B2(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n274_), .B1(new_n281_), .B2(KEYINPUT8), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT8), .ZN(new_n283_));
  AOI211_X1 g082(.A(new_n283_), .B(new_n275_), .C1(new_n277_), .C2(new_n280_), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n261_), .B(new_n264_), .C1(new_n282_), .C2(new_n284_), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n257_), .A2(KEYINPUT35), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n280_), .A2(new_n271_), .A3(new_n276_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n268_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(new_n283_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n281_), .A2(KEYINPUT8), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n290_), .A2(new_n291_), .A3(new_n274_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n292_), .A2(new_n260_), .ZN(new_n293_));
  OAI211_X1 g092(.A(KEYINPUT35), .B(new_n257_), .C1(new_n287_), .C2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G190gat), .B(G218gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G134gat), .B(G162gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n297_), .A2(KEYINPUT36), .ZN(new_n298_));
  INV_X1    g097(.A(new_n292_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(new_n262_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n257_), .A2(KEYINPUT35), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n300_), .A2(new_n285_), .A3(new_n301_), .A4(new_n286_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n294_), .A2(new_n298_), .A3(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  XOR2_X1   g103(.A(new_n297_), .B(KEYINPUT36), .Z(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n306_), .B1(new_n294_), .B2(new_n302_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n252_), .B1(new_n304_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n307_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n309_), .A2(new_n303_), .A3(new_n251_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n250_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n216_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n313_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n290_), .A2(new_n291_), .A3(new_n274_), .A4(new_n216_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(KEYINPUT12), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT12), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n292_), .A2(new_n317_), .A3(new_n313_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G230gat), .A2(G233gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n314_), .A2(new_n315_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n320_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n321_), .A2(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(G120gat), .B(G148gat), .Z(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT65), .B(KEYINPUT5), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G176gat), .B(G204gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n325_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n330_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n321_), .A2(new_n324_), .A3(new_n332_), .ZN(new_n333_));
  AND3_X1   g132(.A1(new_n331_), .A2(KEYINPUT13), .A3(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(KEYINPUT13), .B1(new_n331_), .B2(new_n333_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n209_), .B(new_n260_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G229gat), .A2(G233gat), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n261_), .A2(new_n264_), .A3(new_n209_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n229_), .A2(new_n262_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n341_), .A2(new_n338_), .A3(new_n342_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n340_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G113gat), .B(G141gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G169gat), .B(G197gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n345_), .B(new_n346_), .Z(new_n347_));
  OR2_X1    g146(.A1(new_n347_), .A2(KEYINPUT74), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n344_), .B(new_n348_), .Z(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n336_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G226gat), .A2(G233gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT19), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT95), .ZN(new_n354_));
  INV_X1    g153(.A(G211gat), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n355_), .A2(G218gat), .ZN(new_n356_));
  INV_X1    g155(.A(G218gat), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n357_), .A2(G211gat), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT21), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G197gat), .A2(G204gat), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(G197gat), .A2(G204gat), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n360_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  OR2_X1    g163(.A1(G197gat), .A2(G204gat), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(KEYINPUT21), .A3(new_n361_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n359_), .A2(new_n364_), .A3(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT84), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n357_), .A2(G211gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n355_), .A2(G218gat), .ZN(new_n370_));
  AOI21_X1  g169(.A(KEYINPUT83), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n371_), .A2(new_n366_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n369_), .A2(new_n370_), .A3(KEYINPUT83), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n368_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT83), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n375_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n376_));
  NOR3_X1   g175(.A1(new_n362_), .A2(new_n363_), .A3(new_n360_), .ZN(new_n377_));
  AND4_X1   g176(.A1(new_n368_), .A2(new_n376_), .A3(new_n373_), .A4(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n367_), .B1(new_n374_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G183gat), .A2(G190gat), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT23), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n383_));
  INV_X1    g182(.A(G169gat), .ZN(new_n384_));
  INV_X1    g183(.A(G176gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n382_), .B(new_n383_), .C1(new_n386_), .C2(KEYINPUT24), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT26), .B(G190gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT25), .B(G183gat), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n387_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G169gat), .A2(G176gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT24), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT86), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n392_), .A2(new_n393_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n394_), .B1(new_n393_), .B2(new_n392_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n390_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n385_), .A2(KEYINPUT76), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT76), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(G176gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n384_), .A2(KEYINPUT22), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT22), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(G169gat), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n397_), .A2(new_n399_), .A3(new_n400_), .A4(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(G183gat), .ZN(new_n404_));
  INV_X1    g203(.A(G190gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n382_), .A2(new_n383_), .A3(new_n406_), .ZN(new_n407_));
  AND3_X1   g206(.A1(KEYINPUT87), .A2(G169gat), .A3(G176gat), .ZN(new_n408_));
  AOI21_X1  g207(.A(KEYINPUT87), .B1(G169gat), .B2(G176gat), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n403_), .A2(new_n407_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n396_), .A2(new_n411_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n354_), .B(KEYINPUT20), .C1(new_n379_), .C2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT89), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT75), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n415_), .B1(new_n405_), .B2(KEYINPUT26), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n416_), .B(new_n389_), .C1(new_n388_), .C2(new_n415_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n387_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n386_), .A2(KEYINPUT24), .A3(new_n391_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n417_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n391_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT76), .B(G176gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT22), .B(G169gat), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n421_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT77), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n407_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  AOI211_X1 g225(.A(KEYINPUT77), .B(new_n421_), .C1(new_n422_), .C2(new_n423_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n420_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n379_), .A2(new_n414_), .A3(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n414_), .B1(new_n379_), .B2(new_n428_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n413_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n367_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n376_), .A2(new_n377_), .A3(new_n373_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT84), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n372_), .A2(new_n368_), .A3(new_n373_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n432_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(new_n396_), .A3(new_n411_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n354_), .B1(new_n437_), .B2(KEYINPUT20), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n353_), .B1(new_n431_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT88), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n411_), .A2(new_n440_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n403_), .A2(new_n407_), .A3(KEYINPUT88), .A4(new_n410_), .ZN(new_n442_));
  AOI22_X1  g241(.A1(new_n441_), .A2(new_n442_), .B1(new_n390_), .B2(new_n395_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT20), .B1(new_n443_), .B2(new_n436_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n379_), .A2(new_n428_), .ZN(new_n445_));
  NOR3_X1   g244(.A1(new_n444_), .A2(new_n445_), .A3(new_n353_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n353_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n450_), .B1(new_n443_), .B2(new_n436_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n451_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n353_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT94), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n439_), .A2(new_n447_), .A3(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(G8gat), .B(G36gat), .Z(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT18), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G64gat), .B(G92gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT32), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n456_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT96), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G1gat), .B(G29gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G57gat), .B(G85gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT92), .B(KEYINPUT0), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(G127gat), .B(G134gat), .Z(new_n470_));
  XOR2_X1   g269(.A(G113gat), .B(G120gat), .Z(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G127gat), .B(G134gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G113gat), .B(G120gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n472_), .A2(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(G155gat), .A2(G162gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G155gat), .A2(G162gat), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n477_), .B1(KEYINPUT1), .B2(new_n478_), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n478_), .A2(KEYINPUT1), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G141gat), .A2(G148gat), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(G141gat), .A2(G148gat), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n481_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT3), .ZN(new_n487_));
  INV_X1    g286(.A(G141gat), .ZN(new_n488_));
  INV_X1    g287(.A(G148gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT2), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n482_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n490_), .A2(new_n492_), .A3(new_n493_), .A4(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT81), .ZN(new_n496_));
  XOR2_X1   g295(.A(G155gat), .B(G162gat), .Z(new_n497_));
  AND3_X1   g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n496_), .B1(new_n495_), .B2(new_n497_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n476_), .B(new_n486_), .C1(new_n498_), .C2(new_n499_), .ZN(new_n500_));
  AOI211_X1 g299(.A(new_n483_), .B(new_n484_), .C1(new_n479_), .C2(new_n480_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n495_), .A2(new_n497_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT81), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n501_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT79), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n473_), .A2(new_n474_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n473_), .A2(new_n474_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n506_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n506_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n500_), .B(KEYINPUT4), .C1(new_n505_), .C2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G225gat), .A2(G233gat), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n486_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n510_), .B1(new_n476_), .B2(new_n506_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT90), .B(KEYINPUT4), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n516_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n513_), .A2(KEYINPUT91), .A3(new_n515_), .A4(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n516_), .A2(new_n517_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n521_), .A2(new_n500_), .A3(new_n514_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n519_), .A2(new_n515_), .ZN(new_n524_));
  AOI21_X1  g323(.A(KEYINPUT91), .B1(new_n524_), .B2(new_n513_), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n464_), .B(new_n469_), .C1(new_n523_), .C2(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n469_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT91), .ZN(new_n528_));
  INV_X1    g327(.A(new_n513_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n519_), .A2(new_n515_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n528_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n469_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n531_), .A2(new_n532_), .A3(new_n522_), .A4(new_n520_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n527_), .A2(KEYINPUT96), .A3(new_n533_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n452_), .A2(new_n453_), .A3(KEYINPUT94), .A4(new_n461_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n463_), .A2(new_n526_), .A3(new_n534_), .A4(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT33), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n533_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n460_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n441_), .A2(new_n442_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n396_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n449_), .B1(new_n541_), .B2(new_n379_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n379_), .A2(new_n428_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT89), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n379_), .A2(new_n414_), .A3(new_n428_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n542_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n353_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n448_), .B1(new_n541_), .B2(new_n379_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n403_), .A2(new_n391_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT77), .ZN(new_n550_));
  INV_X1    g349(.A(new_n427_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(new_n551_), .A3(new_n407_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n436_), .A2(new_n552_), .A3(new_n420_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n547_), .B1(new_n548_), .B2(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n539_), .B1(new_n546_), .B2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n452_), .A2(new_n453_), .A3(new_n460_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n521_), .A2(new_n500_), .A3(new_n515_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n559_), .A2(new_n469_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n513_), .A2(new_n514_), .A3(new_n519_), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n560_), .A2(KEYINPUT93), .A3(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(KEYINPUT93), .B1(new_n560_), .B2(new_n561_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n533_), .A2(new_n537_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n538_), .A2(new_n558_), .A3(new_n564_), .A4(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n536_), .A2(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(KEYINPUT79), .B1(new_n472_), .B2(new_n475_), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT31), .B1(new_n568_), .B2(new_n510_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT31), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n509_), .A2(new_n570_), .A3(new_n511_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G71gat), .B(G99gat), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n573_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n569_), .A2(new_n571_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G227gat), .A2(G233gat), .ZN(new_n578_));
  INV_X1    g377(.A(G15gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT30), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n428_), .A2(new_n582_), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n581_), .B(new_n420_), .C1(new_n426_), .C2(new_n427_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(KEYINPUT78), .B(G43gat), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n583_), .A2(new_n584_), .A3(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n586_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n577_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n569_), .A2(new_n575_), .A3(new_n571_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n575_), .B1(new_n569_), .B2(new_n571_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n583_), .A2(new_n584_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(new_n585_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n593_), .A2(new_n595_), .A3(new_n587_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n590_), .A2(new_n596_), .A3(KEYINPUT80), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(KEYINPUT80), .B1(new_n590_), .B2(new_n596_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(G22gat), .B(G50gat), .Z(new_n601_));
  OAI21_X1  g400(.A(new_n601_), .B1(new_n516_), .B2(KEYINPUT29), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT29), .ZN(new_n603_));
  INV_X1    g402(.A(new_n601_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n505_), .A2(new_n603_), .A3(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(KEYINPUT82), .B(KEYINPUT28), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n602_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n606_), .B1(new_n602_), .B2(new_n605_), .ZN(new_n608_));
  OAI21_X1  g407(.A(KEYINPUT85), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n602_), .A2(new_n605_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n606_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT85), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n602_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n612_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n436_), .B1(KEYINPUT29), .B2(new_n516_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G228gat), .A2(G233gat), .ZN(new_n617_));
  INV_X1    g416(.A(G78gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(new_n266_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n616_), .B(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n609_), .A2(new_n615_), .A3(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n379_), .B1(new_n505_), .B2(new_n603_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(new_n620_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n624_), .A2(new_n613_), .A3(new_n614_), .A4(new_n612_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n622_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n600_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n567_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n590_), .A2(new_n596_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT80), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n632_), .A2(new_n625_), .A3(new_n597_), .A4(new_n622_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n626_), .A2(new_n630_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT27), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n546_), .A2(new_n554_), .A3(new_n539_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n460_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n636_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT97), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n557_), .A2(KEYINPUT97), .A3(new_n636_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n534_), .A2(new_n526_), .ZN(new_n644_));
  OAI21_X1  g443(.A(KEYINPUT20), .B1(new_n379_), .B2(new_n412_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT95), .ZN(new_n646_));
  OAI211_X1 g445(.A(new_n646_), .B(new_n413_), .C1(new_n430_), .C2(new_n429_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n446_), .B1(new_n647_), .B2(new_n353_), .ZN(new_n648_));
  OAI211_X1 g447(.A(KEYINPUT27), .B(new_n556_), .C1(new_n648_), .C2(new_n460_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n635_), .A2(new_n643_), .A3(new_n644_), .A4(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n351_), .B1(new_n629_), .B2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n312_), .A2(new_n651_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n652_), .A2(G1gat), .A3(new_n644_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT38), .Z(new_n654_));
  NAND2_X1  g453(.A1(new_n629_), .A2(new_n650_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n304_), .A2(new_n307_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT98), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n244_), .A2(new_n246_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n351_), .A2(new_n660_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n659_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G1gat), .B1(new_n663_), .B2(new_n644_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n654_), .A2(new_n664_), .ZN(G1324gat));
  NAND2_X1  g464(.A1(new_n643_), .A2(new_n649_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n659_), .A2(new_n666_), .A3(new_n661_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT39), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n667_), .A2(new_n668_), .A3(G8gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n667_), .B2(G8gat), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n666_), .A2(new_n205_), .ZN(new_n671_));
  OAI22_X1  g470(.A1(new_n669_), .A2(new_n670_), .B1(new_n652_), .B2(new_n671_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g472(.A(G15gat), .B1(new_n663_), .B2(new_n600_), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n674_), .A2(KEYINPUT41), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(KEYINPUT41), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n652_), .A2(G15gat), .A3(new_n600_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT99), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n675_), .A2(new_n676_), .A3(new_n678_), .ZN(G1326gat));
  OAI21_X1  g478(.A(G22gat), .B1(new_n663_), .B2(new_n626_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n680_), .A2(KEYINPUT42), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n680_), .A2(KEYINPUT42), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n626_), .A2(G22gat), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT100), .Z(new_n684_));
  OAI22_X1  g483(.A1(new_n681_), .A2(new_n682_), .B1(new_n652_), .B2(new_n684_), .ZN(G1327gat));
  NOR2_X1   g484(.A1(new_n249_), .A2(new_n657_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n651_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n644_), .ZN(new_n689_));
  AOI21_X1  g488(.A(G29gat), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n308_), .A2(new_n310_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n691_), .B1(new_n629_), .B2(new_n650_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT101), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(KEYINPUT97), .B1(new_n557_), .B2(new_n636_), .ZN(new_n695_));
  AOI211_X1 g494(.A(new_n640_), .B(KEYINPUT27), .C1(new_n555_), .C2(new_n556_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n644_), .B(new_n649_), .C1(new_n695_), .C2(new_n696_), .ZN(new_n697_));
  AOI22_X1  g496(.A1(new_n622_), .A2(new_n625_), .B1(new_n596_), .B2(new_n590_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n626_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n600_), .B2(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n697_), .A2(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n627_), .B1(new_n536_), .B2(new_n566_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n311_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT101), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n703_), .A2(new_n704_), .A3(KEYINPUT43), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n694_), .A2(new_n705_), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n693_), .B(new_n311_), .C1(new_n701_), .C2(new_n702_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT102), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT102), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n655_), .A2(new_n709_), .A3(new_n693_), .A4(new_n311_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n706_), .A2(new_n711_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n249_), .A2(new_n351_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT44), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n712_), .A2(KEYINPUT44), .A3(new_n713_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n689_), .A2(G29gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n690_), .B1(new_n718_), .B2(new_n719_), .ZN(G1328gat));
  NAND3_X1  g519(.A1(new_n716_), .A2(new_n666_), .A3(new_n717_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(G36gat), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n666_), .A2(KEYINPUT103), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n666_), .A2(KEYINPUT103), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n687_), .A2(G36gat), .A3(new_n726_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT45), .Z(new_n728_));
  NAND2_X1  g527(.A1(new_n722_), .A2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT46), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n722_), .A2(KEYINPUT46), .A3(new_n728_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1329gat));
  NAND4_X1  g532(.A1(new_n716_), .A2(G43gat), .A3(new_n630_), .A4(new_n717_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n687_), .A2(new_n600_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(G43gat), .B2(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g536(.A(G50gat), .B1(new_n688_), .B2(new_n699_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n699_), .A2(G50gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n718_), .B2(new_n739_), .ZN(G1331gat));
  NOR3_X1   g539(.A1(new_n250_), .A2(new_n350_), .A3(new_n336_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n659_), .A2(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n742_), .A2(G57gat), .A3(new_n689_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n743_), .A2(KEYINPUT105), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n743_), .A2(KEYINPUT105), .ZN(new_n745_));
  INV_X1    g544(.A(G57gat), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n336_), .A2(new_n350_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n747_), .A2(new_n655_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n312_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  OR2_X1    g549(.A1(new_n750_), .A2(KEYINPUT104), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(KEYINPUT104), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(new_n689_), .A3(new_n752_), .ZN(new_n753_));
  AOI211_X1 g552(.A(new_n744_), .B(new_n745_), .C1(new_n746_), .C2(new_n753_), .ZN(G1332gat));
  OR3_X1    g553(.A1(new_n749_), .A2(G64gat), .A3(new_n726_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n659_), .A2(new_n725_), .A3(new_n741_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT48), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n756_), .A2(new_n757_), .A3(G64gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n756_), .B2(G64gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n755_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT106), .ZN(G1333gat));
  OR3_X1    g560(.A1(new_n749_), .A2(G71gat), .A3(new_n600_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n600_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n659_), .A2(new_n763_), .A3(new_n741_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT49), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n764_), .A2(new_n765_), .A3(G71gat), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n764_), .B2(G71gat), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n762_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  XOR2_X1   g567(.A(new_n768_), .B(KEYINPUT107), .Z(G1334gat));
  NAND3_X1  g568(.A1(new_n750_), .A2(new_n618_), .A3(new_n699_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n742_), .A2(new_n699_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n771_), .A2(G78gat), .A3(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n771_), .B2(G78gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n770_), .B1(new_n773_), .B2(new_n774_), .ZN(G1335gat));
  INV_X1    g574(.A(G85gat), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n250_), .A2(new_n747_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n777_), .B1(new_n706_), .B2(new_n711_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n776_), .B1(new_n778_), .B2(new_n689_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n748_), .A2(new_n686_), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n780_), .A2(new_n776_), .A3(new_n689_), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1336gat));
  AOI21_X1  g581(.A(G92gat), .B1(new_n780_), .B2(new_n666_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n725_), .A2(G92gat), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT109), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n783_), .B1(new_n778_), .B2(new_n785_), .ZN(G1337gat));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n630_), .A2(new_n265_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n780_), .A2(new_n788_), .ZN(new_n789_));
  AOI211_X1 g588(.A(new_n600_), .B(new_n777_), .C1(new_n706_), .C2(new_n711_), .ZN(new_n790_));
  INV_X1    g589(.A(G99gat), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n787_), .B(new_n789_), .C1(new_n790_), .C2(new_n791_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(KEYINPUT112), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n789_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT110), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n787_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  OAI211_X1 g595(.A(KEYINPUT110), .B(new_n789_), .C1(new_n790_), .C2(new_n791_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT111), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n791_), .B1(new_n778_), .B2(new_n763_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n789_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n795_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  AND4_X1   g600(.A1(KEYINPUT111), .A2(new_n801_), .A3(KEYINPUT51), .A4(new_n797_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n793_), .B1(new_n798_), .B2(new_n802_), .ZN(G1338gat));
  NAND3_X1  g602(.A1(new_n780_), .A2(new_n266_), .A3(new_n699_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n778_), .A2(new_n699_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(G106gat), .ZN(new_n807_));
  AOI211_X1 g606(.A(KEYINPUT52), .B(new_n266_), .C1(new_n778_), .C2(new_n699_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n804_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g609(.A1(new_n689_), .A2(new_n698_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n666_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n316_), .A2(new_n323_), .A3(new_n318_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n321_), .A2(KEYINPUT55), .A3(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n323_), .B1(new_n316_), .B2(new_n318_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n332_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n815_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT56), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n815_), .A2(KEYINPUT56), .A3(new_n818_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n333_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n824_), .A2(new_n349_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n331_), .A2(new_n333_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n341_), .A2(new_n342_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n341_), .A2(KEYINPUT116), .A3(new_n342_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n339_), .A3(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n347_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  AOI22_X1  g632(.A1(new_n833_), .A2(KEYINPUT117), .B1(new_n347_), .B2(new_n344_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n831_), .A2(new_n835_), .A3(new_n832_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n823_), .A2(new_n825_), .B1(new_n826_), .B2(new_n838_), .ZN(new_n839_));
  OAI211_X1 g638(.A(KEYINPUT118), .B(KEYINPUT57), .C1(new_n839_), .C2(new_n656_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n815_), .A2(KEYINPUT56), .A3(new_n818_), .ZN(new_n842_));
  AOI21_X1  g641(.A(KEYINPUT56), .B1(new_n815_), .B2(new_n818_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n825_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n826_), .A2(new_n838_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n656_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n841_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n840_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n822_), .A2(KEYINPUT120), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT120), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n815_), .A2(new_n818_), .A3(new_n851_), .A4(KEYINPUT56), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n850_), .A2(new_n821_), .A3(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(KEYINPUT119), .B1(new_n837_), .B2(new_n824_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n333_), .A2(new_n834_), .A3(new_n855_), .A4(new_n836_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n853_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT58), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n691_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n853_), .A2(new_n857_), .A3(KEYINPUT58), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(KEYINPUT121), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT121), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n853_), .A2(new_n857_), .A3(new_n863_), .A4(KEYINPUT58), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n860_), .A2(new_n862_), .A3(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n849_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT122), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n849_), .A2(new_n865_), .A3(KEYINPUT122), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n868_), .A2(new_n660_), .A3(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT73), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n660_), .A2(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n244_), .A2(new_n246_), .A3(KEYINPUT73), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n872_), .A2(new_n349_), .A3(new_n336_), .A4(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT113), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n311_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n249_), .A2(KEYINPUT113), .A3(new_n349_), .A4(new_n336_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n879_));
  XOR2_X1   g678(.A(new_n879_), .B(KEYINPUT115), .Z(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n878_), .A2(new_n881_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n879_), .A2(KEYINPUT115), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n878_), .B2(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n813_), .B1(new_n870_), .B2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(G113gat), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n885_), .A2(new_n886_), .A3(new_n350_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n878_), .A2(new_n883_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n880_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n866_), .A2(new_n250_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n888_), .B(new_n812_), .C1(new_n891_), .C2(new_n893_), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n894_), .B(new_n350_), .C1(new_n885_), .C2(new_n888_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n887_), .B1(new_n896_), .B2(new_n886_), .ZN(G1340gat));
  INV_X1    g696(.A(G120gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n898_), .B1(new_n336_), .B2(KEYINPUT60), .ZN(new_n899_));
  OAI211_X1 g698(.A(new_n885_), .B(new_n899_), .C1(KEYINPUT60), .C2(new_n898_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n336_), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n894_), .B(new_n901_), .C1(new_n885_), .C2(new_n888_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n900_), .B1(new_n903_), .B2(new_n898_), .ZN(G1341gat));
  INV_X1    g703(.A(G127gat), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n885_), .A2(new_n905_), .A3(new_n249_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n660_), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n894_), .B(new_n907_), .C1(new_n885_), .C2(new_n888_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n906_), .B1(new_n909_), .B2(new_n905_), .ZN(G1342gat));
  INV_X1    g709(.A(G134gat), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n885_), .A2(new_n911_), .A3(new_n656_), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n894_), .B(new_n311_), .C1(new_n885_), .C2(new_n888_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n912_), .B1(new_n914_), .B2(new_n911_), .ZN(G1343gat));
  NAND2_X1  g714(.A1(new_n870_), .A2(new_n884_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n633_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n725_), .A2(new_n644_), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n916_), .A2(new_n917_), .A3(new_n350_), .A4(new_n918_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G141gat), .ZN(G1344gat));
  NAND4_X1  g719(.A1(new_n916_), .A2(new_n917_), .A3(new_n901_), .A4(new_n918_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g721(.A1(new_n916_), .A2(new_n917_), .A3(new_n249_), .A4(new_n918_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(KEYINPUT61), .B(G155gat), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n923_), .B(new_n924_), .ZN(G1346gat));
  NAND2_X1  g724(.A1(new_n916_), .A2(new_n917_), .ZN(new_n926_));
  NOR3_X1   g725(.A1(new_n926_), .A2(new_n644_), .A3(new_n725_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n311_), .A2(G162gat), .ZN(new_n928_));
  XOR2_X1   g727(.A(new_n928_), .B(KEYINPUT123), .Z(new_n929_));
  INV_X1    g728(.A(G162gat), .ZN(new_n930_));
  NAND4_X1  g729(.A1(new_n916_), .A2(new_n917_), .A3(new_n656_), .A4(new_n918_), .ZN(new_n931_));
  AOI22_X1  g730(.A1(new_n927_), .A2(new_n929_), .B1(new_n930_), .B2(new_n931_), .ZN(G1347gat));
  NOR2_X1   g731(.A1(new_n726_), .A2(new_n689_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(new_n763_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n934_), .A2(new_n699_), .ZN(new_n935_));
  OAI211_X1 g734(.A(new_n350_), .B(new_n935_), .C1(new_n891_), .C2(new_n893_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n384_), .B1(new_n937_), .B2(KEYINPUT62), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n936_), .A2(new_n938_), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT62), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n939_), .A2(KEYINPUT124), .A3(new_n940_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n935_), .B1(new_n891_), .B2(new_n893_), .ZN(new_n942_));
  INV_X1    g741(.A(new_n942_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n943_), .A2(new_n423_), .A3(new_n350_), .ZN(new_n944_));
  OAI211_X1 g743(.A(new_n936_), .B(new_n938_), .C1(new_n937_), .C2(KEYINPUT62), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n941_), .A2(new_n944_), .A3(new_n945_), .ZN(G1348gat));
  INV_X1    g745(.A(new_n422_), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n947_), .B1(new_n943_), .B2(new_n901_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n699_), .B1(new_n870_), .B2(new_n884_), .ZN(new_n949_));
  INV_X1    g748(.A(KEYINPUT125), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n949_), .B(new_n950_), .ZN(new_n951_));
  NOR3_X1   g750(.A1(new_n934_), .A2(new_n385_), .A3(new_n336_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n948_), .B1(new_n951_), .B2(new_n952_), .ZN(G1349gat));
  NOR3_X1   g752(.A1(new_n942_), .A2(new_n389_), .A3(new_n660_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n934_), .A2(new_n250_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n950_), .B1(new_n916_), .B2(new_n626_), .ZN(new_n956_));
  AOI211_X1 g755(.A(KEYINPUT125), .B(new_n699_), .C1(new_n870_), .C2(new_n884_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n955_), .B1(new_n956_), .B2(new_n957_), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n954_), .B1(new_n958_), .B2(new_n404_), .ZN(G1350gat));
  OAI21_X1  g758(.A(G190gat), .B1(new_n942_), .B2(new_n691_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n656_), .A2(new_n388_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n961_), .B(KEYINPUT126), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n960_), .B1(new_n942_), .B2(new_n962_), .ZN(G1351gat));
  NAND4_X1  g762(.A1(new_n916_), .A2(new_n917_), .A3(new_n350_), .A4(new_n933_), .ZN(new_n964_));
  XNOR2_X1  g763(.A(new_n964_), .B(G197gat), .ZN(G1352gat));
  NAND4_X1  g764(.A1(new_n916_), .A2(new_n917_), .A3(new_n901_), .A4(new_n933_), .ZN(new_n966_));
  XNOR2_X1  g765(.A(new_n966_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g766(.A(new_n660_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n968_));
  NAND4_X1  g767(.A1(new_n916_), .A2(new_n917_), .A3(new_n933_), .A4(new_n968_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n970_));
  XOR2_X1   g769(.A(new_n970_), .B(KEYINPUT127), .Z(new_n971_));
  XNOR2_X1  g770(.A(new_n969_), .B(new_n971_), .ZN(G1354gat));
  NOR2_X1   g771(.A1(new_n657_), .A2(G218gat), .ZN(new_n973_));
  NAND4_X1  g772(.A1(new_n916_), .A2(new_n917_), .A3(new_n933_), .A4(new_n973_), .ZN(new_n974_));
  NOR4_X1   g773(.A1(new_n926_), .A2(new_n689_), .A3(new_n691_), .A4(new_n726_), .ZN(new_n975_));
  OAI21_X1  g774(.A(new_n974_), .B1(new_n975_), .B2(new_n357_), .ZN(G1355gat));
endmodule


