//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 0 0 1 1 1 0 0 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n619_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n800_, new_n801_,
    new_n802_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n819_, new_n820_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n856_, new_n857_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n883_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XOR2_X1   g006(.A(new_n206_), .B(new_n207_), .Z(new_n208_));
  XOR2_X1   g007(.A(G29gat), .B(G36gat), .Z(new_n209_));
  XOR2_X1   g008(.A(G43gat), .B(G50gat), .Z(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n208_), .B(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT72), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G229gat), .A2(G233gat), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n211_), .B(KEYINPUT15), .ZN(new_n217_));
  INV_X1    g016(.A(new_n208_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n216_), .B1(new_n208_), .B2(new_n211_), .ZN(new_n220_));
  AOI22_X1  g019(.A1(new_n214_), .A2(new_n216_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  XOR2_X1   g020(.A(G113gat), .B(G141gat), .Z(new_n222_));
  XNOR2_X1  g021(.A(G169gat), .B(G197gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n221_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n221_), .A2(new_n224_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G57gat), .B(G64gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT11), .ZN(new_n230_));
  XOR2_X1   g029(.A(G71gat), .B(G78gat), .Z(new_n231_));
  NOR2_X1   g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n230_), .A2(new_n231_), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n229_), .A2(KEYINPUT11), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n232_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  OR2_X1    g035(.A1(G85gat), .A2(G92gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G85gat), .A2(G92gat), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(G99gat), .A2(G106gat), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT7), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G99gat), .A2(G106gat), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT6), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n239_), .B1(new_n242_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT8), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n247_), .A2(KEYINPUT66), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n246_), .B(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT10), .B(G99gat), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT64), .B(G106gat), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n245_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT9), .ZN(new_n254_));
  AND3_X1   g053(.A1(new_n238_), .A2(KEYINPUT65), .A3(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT65), .B1(new_n238_), .B2(new_n254_), .ZN(new_n256_));
  OAI221_X1 g055(.A(new_n237_), .B1(new_n254_), .B2(new_n238_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n253_), .A2(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n236_), .B1(new_n249_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT12), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n260_), .B(KEYINPUT67), .Z(new_n261_));
  NAND3_X1  g060(.A1(new_n249_), .A2(new_n258_), .A3(new_n236_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n262_), .B1(new_n259_), .B2(KEYINPUT12), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G230gat), .A2(G233gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n262_), .ZN(new_n267_));
  OAI211_X1 g066(.A(G230gat), .B(G233gat), .C1(new_n267_), .C2(new_n259_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G120gat), .B(G148gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT5), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G176gat), .B(G204gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT68), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n269_), .A2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n266_), .A2(new_n268_), .A3(new_n273_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n278_), .A2(KEYINPUT13), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(KEYINPUT13), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n279_), .A2(KEYINPUT69), .A3(new_n280_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n228_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G226gat), .A2(G233gat), .ZN(new_n286_));
  XOR2_X1   g085(.A(new_n286_), .B(KEYINPUT19), .Z(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT20), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT25), .B(G183gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT26), .B(G190gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT23), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(G169gat), .ZN(new_n297_));
  INV_X1    g096(.A(G176gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n299_), .A2(KEYINPUT24), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G169gat), .A2(G176gat), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n299_), .A2(KEYINPUT24), .A3(new_n301_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n291_), .A2(new_n296_), .A3(new_n300_), .A4(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(G183gat), .ZN(new_n304_));
  INV_X1    g103(.A(G190gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n294_), .A2(new_n295_), .A3(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT74), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(G176gat), .B1(KEYINPUT73), .B2(KEYINPUT22), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(G169gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n307_), .A2(new_n308_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n303_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(G204gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(G197gat), .ZN(new_n316_));
  INV_X1    g115(.A(G197gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(G204gat), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT21), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G211gat), .B(G218gat), .ZN(new_n321_));
  OR3_X1    g120(.A1(new_n319_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n316_), .A2(new_n318_), .A3(new_n320_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT84), .ZN(new_n324_));
  AND3_X1   g123(.A1(new_n316_), .A2(new_n318_), .A3(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(KEYINPUT21), .B1(new_n316_), .B2(new_n324_), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n323_), .B(new_n321_), .C1(new_n325_), .C2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n322_), .A2(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n288_), .B1(new_n314_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n297_), .A2(KEYINPUT22), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT22), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(G169gat), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n330_), .A2(new_n332_), .A3(new_n298_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT87), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n333_), .A2(new_n334_), .A3(new_n301_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n334_), .B1(new_n333_), .B2(new_n301_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n307_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT88), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT88), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n339_), .B(new_n307_), .C1(new_n335_), .C2(new_n336_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n338_), .A2(new_n340_), .A3(new_n303_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n329_), .B1(new_n341_), .B2(new_n328_), .ZN(new_n342_));
  XOR2_X1   g141(.A(G8gat), .B(G36gat), .Z(new_n343_));
  XNOR2_X1  g142(.A(G64gat), .B(G92gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT20), .B1(new_n314_), .B2(new_n328_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n348_), .B1(new_n341_), .B2(new_n328_), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n342_), .B(new_n347_), .C1(new_n349_), .C2(new_n287_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT101), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n322_), .A2(new_n327_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n353_), .A2(new_n337_), .A3(new_n303_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n314_), .A2(new_n328_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT98), .B(KEYINPUT20), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n287_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n359_), .A2(KEYINPUT99), .ZN(new_n360_));
  INV_X1    g159(.A(new_n303_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n361_), .B1(new_n337_), .B2(KEYINPUT88), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n353_), .B1(new_n362_), .B2(new_n340_), .ZN(new_n363_));
  NOR3_X1   g162(.A1(new_n363_), .A2(new_n358_), .A3(new_n348_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n359_), .A2(KEYINPUT99), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n360_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n352_), .B1(new_n366_), .B2(new_n347_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n350_), .A2(new_n351_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT27), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT90), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n350_), .A2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n358_), .B1(new_n363_), .B2(new_n348_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n372_), .A2(KEYINPUT90), .A3(new_n342_), .A4(new_n347_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n342_), .B1(new_n349_), .B2(new_n287_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n347_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n371_), .A2(new_n373_), .A3(new_n376_), .ZN(new_n377_));
  OR2_X1    g176(.A1(new_n377_), .A2(KEYINPUT27), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n369_), .A2(new_n378_), .ZN(new_n379_));
  XOR2_X1   g178(.A(KEYINPUT82), .B(KEYINPUT28), .Z(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G22gat), .B(G50gat), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT78), .ZN(new_n383_));
  INV_X1    g182(.A(G155gat), .ZN(new_n384_));
  INV_X1    g183(.A(G162gat), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n383_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G155gat), .A2(G162gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT1), .ZN(new_n388_));
  OAI21_X1  g187(.A(KEYINPUT78), .B1(G155gat), .B2(G162gat), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n386_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT79), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT80), .B1(new_n387_), .B2(KEYINPUT1), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT80), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT1), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n393_), .A2(new_n394_), .A3(G155gat), .A4(G162gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n392_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT79), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n386_), .A2(new_n388_), .A3(new_n398_), .A4(new_n389_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n391_), .A2(new_n397_), .A3(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G141gat), .A2(G148gat), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(G141gat), .A2(G148gat), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n400_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n386_), .A2(new_n389_), .A3(new_n387_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(G141gat), .ZN(new_n408_));
  INV_X1    g207(.A(G148gat), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(new_n409_), .A3(KEYINPUT3), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT3), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n411_), .B1(G141gat), .B2(G148gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  AND3_X1   g212(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n414_));
  AOI21_X1  g213(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT81), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n413_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n417_), .B1(new_n413_), .B2(new_n416_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n407_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n405_), .A2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n382_), .B1(new_n421_), .B2(KEYINPUT29), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NOR3_X1   g222(.A1(new_n421_), .A2(KEYINPUT29), .A3(new_n382_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n381_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n424_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n426_), .A2(new_n380_), .A3(new_n422_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n353_), .B1(new_n421_), .B2(KEYINPUT29), .ZN(new_n430_));
  INV_X1    g229(.A(G228gat), .ZN(new_n431_));
  INV_X1    g230(.A(G233gat), .ZN(new_n432_));
  OR2_X1    g231(.A1(new_n432_), .A2(KEYINPUT83), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(KEYINPUT83), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n431_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT85), .ZN(new_n436_));
  OR2_X1    g235(.A1(new_n430_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G78gat), .B(G106gat), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT85), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n435_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n430_), .A2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n437_), .A2(new_n439_), .A3(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT86), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n429_), .A2(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n439_), .B1(new_n437_), .B2(new_n442_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n443_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n446_), .A2(new_n449_), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n429_), .A2(new_n445_), .B1(new_n448_), .B2(new_n443_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n379_), .A2(new_n453_), .ZN(new_n454_));
  XOR2_X1   g253(.A(G127gat), .B(G134gat), .Z(new_n455_));
  XOR2_X1   g254(.A(G113gat), .B(G120gat), .Z(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n404_), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n386_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n396_), .B1(new_n460_), .B2(new_n398_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n459_), .B1(new_n461_), .B2(new_n391_), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n410_), .A2(new_n412_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n415_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT81), .B1(new_n463_), .B2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n413_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n406_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n458_), .B1(new_n462_), .B2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n405_), .A2(new_n420_), .A3(new_n457_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(KEYINPUT4), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G225gat), .A2(G233gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT92), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n457_), .B1(new_n405_), .B2(new_n420_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT93), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT4), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n475_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n476_), .B1(new_n475_), .B2(new_n477_), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n472_), .B(new_n474_), .C1(new_n478_), .C2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n470_), .A2(new_n471_), .A3(new_n473_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT94), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT94), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n470_), .A2(new_n483_), .A3(new_n471_), .A4(new_n473_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n482_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n480_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G1gat), .B(G29gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(G85gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT0), .B(G57gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n486_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n490_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n480_), .A2(new_n485_), .A3(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G227gat), .A2(G233gat), .ZN(new_n496_));
  INV_X1    g295(.A(G71gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(G99gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n314_), .B(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G15gat), .B(G43gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT75), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n502_), .B(KEYINPUT30), .Z(new_n503_));
  XNOR2_X1  g302(.A(new_n500_), .B(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT77), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n457_), .B(KEYINPUT31), .Z(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT76), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT77), .B1(new_n504_), .B2(new_n508_), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n506_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n454_), .A2(new_n495_), .A3(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n495_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n516_), .B1(new_n378_), .B2(new_n369_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n371_), .A2(new_n376_), .A3(KEYINPUT91), .A4(new_n373_), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n493_), .A2(KEYINPUT95), .A3(KEYINPUT33), .ZN(new_n519_));
  AOI21_X1  g318(.A(KEYINPUT33), .B1(new_n493_), .B2(KEYINPUT95), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n518_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT91), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n377_), .A2(new_n522_), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n472_), .B(new_n473_), .C1(new_n478_), .C2(new_n479_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n470_), .A2(new_n471_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n492_), .B1(new_n525_), .B2(new_n474_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n523_), .A2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT96), .B1(new_n521_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n493_), .A2(KEYINPUT95), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT33), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n493_), .A2(KEYINPUT95), .A3(KEYINPUT33), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT96), .ZN(new_n535_));
  AOI22_X1  g334(.A1(new_n377_), .A2(new_n522_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n534_), .A2(new_n535_), .A3(new_n536_), .A4(new_n518_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT100), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n347_), .A2(KEYINPUT32), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n538_), .B1(new_n366_), .B2(new_n539_), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n365_), .A2(new_n364_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n539_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n541_), .A2(KEYINPUT100), .A3(new_n360_), .A4(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n372_), .A2(new_n342_), .A3(new_n539_), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n545_), .B(KEYINPUT97), .Z(new_n546_));
  NAND3_X1  g345(.A1(new_n544_), .A2(new_n494_), .A3(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n529_), .A2(new_n537_), .A3(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n517_), .B1(new_n548_), .B2(new_n452_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n515_), .B1(new_n549_), .B2(new_n514_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n249_), .A2(new_n258_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT35), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G232gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT34), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  AOI22_X1  g354(.A1(new_n551_), .A2(new_n217_), .B1(new_n552_), .B2(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n556_), .B1(new_n551_), .B2(new_n212_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n555_), .A2(new_n552_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n557_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G190gat), .B(G218gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G134gat), .B(G162gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n563_), .A2(KEYINPUT36), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n560_), .A2(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n563_), .B(KEYINPUT36), .Z(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n565_), .B1(new_n560_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT70), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT37), .ZN(new_n570_));
  NOR3_X1   g369(.A1(new_n568_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n570_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G127gat), .B(G155gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT16), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G183gat), .B(G211gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n208_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(new_n235_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT71), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n578_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT17), .B1(new_n581_), .B2(new_n578_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  OAI211_X1 g384(.A(KEYINPUT17), .B(new_n578_), .C1(new_n581_), .C2(new_n582_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n574_), .A2(new_n588_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n285_), .A2(new_n550_), .A3(new_n589_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n494_), .A2(KEYINPUT102), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n494_), .A2(KEYINPUT102), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n590_), .A2(new_n203_), .A3(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n595_), .B(KEYINPUT38), .Z(new_n596_));
  NAND2_X1  g395(.A1(new_n550_), .A2(new_n568_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT103), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n598_), .A2(new_n285_), .A3(new_n587_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n203_), .B1(new_n599_), .B2(new_n494_), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n596_), .A2(new_n600_), .ZN(G1324gat));
  NAND3_X1  g400(.A1(new_n590_), .A2(new_n204_), .A3(new_n379_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT39), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n599_), .A2(new_n379_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n603_), .B1(new_n604_), .B2(G8gat), .ZN(new_n605_));
  AOI211_X1 g404(.A(KEYINPUT39), .B(new_n204_), .C1(new_n599_), .C2(new_n379_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n602_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n607_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g407(.A(G15gat), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n609_), .B1(new_n599_), .B2(new_n514_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT41), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n590_), .A2(new_n609_), .A3(new_n514_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(G1326gat));
  INV_X1    g412(.A(G22gat), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n614_), .B1(new_n599_), .B2(new_n453_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT42), .Z(new_n616_));
  NAND2_X1  g415(.A1(new_n453_), .A2(new_n614_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT104), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n590_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n616_), .A2(new_n619_), .ZN(G1327gat));
  INV_X1    g419(.A(G29gat), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT105), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n550_), .A2(new_n622_), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n515_), .B(KEYINPUT105), .C1(new_n549_), .C2(new_n514_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n573_), .ZN(new_n625_));
  OAI21_X1  g424(.A(KEYINPUT106), .B1(new_n625_), .B2(new_n571_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT106), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n572_), .A2(new_n627_), .A3(new_n573_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n623_), .A2(new_n624_), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(KEYINPUT43), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT43), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n550_), .A2(new_n633_), .A3(new_n574_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT109), .ZN(new_n636_));
  AOI211_X1 g435(.A(new_n228_), .B(new_n587_), .C1(new_n283_), .C2(new_n284_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n635_), .A2(new_n636_), .A3(KEYINPUT44), .A4(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n629_), .B1(new_n550_), .B2(new_n622_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n633_), .B1(new_n639_), .B2(new_n624_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n634_), .ZN(new_n641_));
  OAI211_X1 g440(.A(KEYINPUT44), .B(new_n637_), .C1(new_n640_), .C2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT109), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n638_), .A2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n641_), .B1(new_n631_), .B2(KEYINPUT43), .ZN(new_n645_));
  INV_X1    g444(.A(new_n637_), .ZN(new_n646_));
  OAI21_X1  g445(.A(KEYINPUT107), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT107), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n648_), .B(new_n637_), .C1(new_n640_), .C2(new_n641_), .ZN(new_n649_));
  XOR2_X1   g448(.A(KEYINPUT108), .B(KEYINPUT44), .Z(new_n650_));
  NAND3_X1  g449(.A1(new_n647_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n644_), .A2(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n621_), .B1(new_n652_), .B2(new_n594_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n568_), .A2(new_n587_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n285_), .A2(new_n550_), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT110), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n285_), .A2(KEYINPUT110), .A3(new_n550_), .A4(new_n654_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n659_), .A2(G29gat), .A3(new_n495_), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n653_), .A2(new_n660_), .ZN(G1328gat));
  INV_X1    g460(.A(new_n379_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(G36gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n657_), .A2(new_n658_), .A3(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT112), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT112), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n657_), .A2(new_n666_), .A3(new_n658_), .A4(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT45), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n644_), .A2(new_n379_), .A3(new_n651_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n670_), .A2(KEYINPUT111), .A3(G36gat), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT111), .B1(new_n670_), .B2(G36gat), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n669_), .B(KEYINPUT46), .C1(new_n672_), .C2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT45), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n668_), .B(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n673_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n677_), .B2(new_n671_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(KEYINPUT113), .B(KEYINPUT46), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n674_), .B1(new_n678_), .B2(new_n679_), .ZN(G1329gat));
  INV_X1    g479(.A(G43gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n681_), .B1(new_n652_), .B2(new_n514_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT47), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n659_), .A2(G43gat), .A3(new_n513_), .ZN(new_n684_));
  OR3_X1    g483(.A1(new_n682_), .A2(new_n683_), .A3(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n683_), .B1(new_n682_), .B2(new_n684_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1330gat));
  OR3_X1    g486(.A1(new_n659_), .A2(G50gat), .A3(new_n452_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n644_), .A2(new_n453_), .A3(new_n651_), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n689_), .A2(KEYINPUT114), .A3(G50gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT114), .B1(new_n689_), .B2(G50gat), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n688_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT115), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT115), .ZN(new_n694_));
  OAI211_X1 g493(.A(new_n694_), .B(new_n688_), .C1(new_n690_), .C2(new_n691_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(G1331gat));
  INV_X1    g495(.A(G57gat), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n283_), .A2(new_n284_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n228_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n701_), .A2(new_n588_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n702_), .A2(new_n598_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n697_), .B1(new_n703_), .B2(new_n494_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n700_), .A2(new_n550_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n705_), .A2(new_n588_), .A3(new_n574_), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n706_), .A2(new_n697_), .A3(new_n594_), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n704_), .A2(new_n707_), .ZN(G1332gat));
  INV_X1    g507(.A(G64gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n703_), .B2(new_n379_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT48), .Z(new_n711_));
  NAND3_X1  g510(.A1(new_n706_), .A2(new_n709_), .A3(new_n379_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1333gat));
  AOI21_X1  g512(.A(new_n497_), .B1(new_n703_), .B2(new_n514_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT49), .Z(new_n715_));
  NOR2_X1   g514(.A1(new_n513_), .A2(G71gat), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT116), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n706_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n715_), .A2(new_n718_), .ZN(G1334gat));
  INV_X1    g518(.A(G78gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n720_), .B1(new_n703_), .B2(new_n453_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT50), .Z(new_n722_));
  NAND3_X1  g521(.A1(new_n706_), .A2(new_n720_), .A3(new_n453_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1335gat));
  NOR3_X1   g523(.A1(new_n645_), .A2(new_n701_), .A3(new_n587_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT117), .ZN(new_n726_));
  OAI21_X1  g525(.A(G85gat), .B1(new_n726_), .B2(new_n495_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n705_), .A2(new_n568_), .A3(new_n587_), .ZN(new_n728_));
  INV_X1    g527(.A(G85gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n728_), .A2(new_n729_), .A3(new_n594_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n727_), .A2(new_n730_), .ZN(G1336gat));
  AOI21_X1  g530(.A(G92gat), .B1(new_n728_), .B2(new_n379_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n726_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n379_), .A2(G92gat), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT118), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n732_), .B1(new_n733_), .B2(new_n735_), .ZN(G1337gat));
  NAND2_X1  g535(.A1(new_n725_), .A2(new_n514_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(G99gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n728_), .A2(new_n251_), .A3(new_n514_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g540(.A1(new_n728_), .A2(new_n252_), .A3(new_n453_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n725_), .A2(new_n453_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(G106gat), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n744_), .A2(KEYINPUT52), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n744_), .A2(KEYINPUT52), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n742_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g547(.A1(new_n281_), .A2(new_n589_), .A3(new_n228_), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT54), .Z(new_n750_));
  OAI21_X1  g549(.A(KEYINPUT55), .B1(new_n264_), .B2(new_n265_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(new_n266_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n264_), .A2(KEYINPUT55), .A3(new_n265_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n274_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT56), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n277_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT119), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n699_), .B1(new_n754_), .B2(new_n757_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n756_), .A2(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n754_), .A2(new_n757_), .A3(new_n755_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n214_), .A2(new_n215_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n215_), .B1(new_n208_), .B2(new_n211_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n224_), .B1(new_n219_), .B2(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n226_), .B1(new_n761_), .B2(new_n763_), .ZN(new_n764_));
  AOI22_X1  g563(.A1(new_n759_), .A2(new_n760_), .B1(new_n278_), .B2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT57), .ZN(new_n766_));
  INV_X1    g565(.A(new_n568_), .ZN(new_n767_));
  OR3_X1    g566(.A1(new_n765_), .A2(new_n766_), .A3(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n766_), .B1(new_n765_), .B2(new_n767_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n754_), .A2(new_n755_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n764_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n771_), .A2(new_n756_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT58), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT120), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n574_), .B1(new_n772_), .B2(KEYINPUT58), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n768_), .B(new_n769_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n750_), .B1(new_n776_), .B2(new_n588_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n777_), .A2(KEYINPUT121), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT121), .ZN(new_n779_));
  AOI211_X1 g578(.A(new_n779_), .B(new_n750_), .C1(new_n776_), .C2(new_n588_), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n454_), .A2(new_n514_), .A3(new_n594_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n781_), .A2(new_n699_), .A3(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(G113gat), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n777_), .A2(KEYINPUT59), .A3(new_n782_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n783_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n787_), .B2(KEYINPUT59), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n228_), .A2(new_n785_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT122), .ZN(new_n790_));
  AOI22_X1  g589(.A1(new_n784_), .A2(new_n785_), .B1(new_n788_), .B2(new_n790_), .ZN(G1340gat));
  INV_X1    g590(.A(new_n698_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT60), .ZN(new_n793_));
  AOI21_X1  g592(.A(G120gat), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n794_), .B1(new_n793_), .B2(G120gat), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n781_), .A2(new_n783_), .A3(new_n795_), .ZN(new_n796_));
  AOI211_X1 g595(.A(new_n698_), .B(new_n786_), .C1(new_n787_), .C2(KEYINPUT59), .ZN(new_n797_));
  INV_X1    g596(.A(G120gat), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n796_), .B1(new_n797_), .B2(new_n798_), .ZN(G1341gat));
  AOI211_X1 g598(.A(new_n588_), .B(new_n786_), .C1(new_n787_), .C2(KEYINPUT59), .ZN(new_n800_));
  INV_X1    g599(.A(G127gat), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n587_), .A2(new_n801_), .ZN(new_n802_));
  OAI22_X1  g601(.A1(new_n800_), .A2(new_n801_), .B1(new_n787_), .B2(new_n802_), .ZN(G1342gat));
  OAI211_X1 g602(.A(new_n767_), .B(new_n783_), .C1(new_n778_), .C2(new_n780_), .ZN(new_n804_));
  INV_X1    g603(.A(G134gat), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT123), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT123), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n804_), .A2(new_n808_), .A3(new_n805_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n574_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n810_), .A2(new_n805_), .ZN(new_n811_));
  AOI22_X1  g610(.A1(new_n807_), .A2(new_n809_), .B1(new_n788_), .B2(new_n811_), .ZN(G1343gat));
  NOR4_X1   g611(.A1(new_n379_), .A2(new_n593_), .A3(new_n514_), .A4(new_n452_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n781_), .A2(new_n699_), .A3(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(G141gat), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n781_), .A2(new_n408_), .A3(new_n699_), .A4(new_n813_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(G1344gat));
  NAND3_X1  g616(.A1(new_n781_), .A2(new_n792_), .A3(new_n813_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(G148gat), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n781_), .A2(new_n409_), .A3(new_n792_), .A4(new_n813_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(G1345gat));
  NAND3_X1  g620(.A1(new_n781_), .A2(new_n587_), .A3(new_n813_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(KEYINPUT61), .B(G155gat), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n823_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n781_), .A2(new_n587_), .A3(new_n813_), .A4(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(G1346gat));
  AND2_X1   g626(.A1(new_n781_), .A2(new_n813_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n629_), .A2(new_n385_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n781_), .A2(new_n767_), .A3(new_n813_), .ZN(new_n830_));
  AOI22_X1  g629(.A1(new_n828_), .A2(new_n829_), .B1(new_n830_), .B2(new_n385_), .ZN(G1347gat));
  INV_X1    g630(.A(new_n777_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n662_), .A2(new_n513_), .A3(new_n594_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n832_), .A2(new_n452_), .A3(new_n699_), .A4(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(G169gat), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT124), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n834_), .A2(KEYINPUT124), .A3(G169gat), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(KEYINPUT62), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n330_), .A2(new_n332_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n834_), .A2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT124), .B1(new_n834_), .B2(G169gat), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT62), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n841_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n839_), .A2(new_n844_), .ZN(G1348gat));
  NAND2_X1  g644(.A1(new_n832_), .A2(new_n452_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n833_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(G176gat), .B1(new_n848_), .B2(new_n792_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n781_), .A2(new_n452_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n698_), .A2(new_n298_), .A3(new_n847_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n849_), .B1(new_n850_), .B2(new_n851_), .ZN(G1349gat));
  NOR4_X1   g651(.A1(new_n846_), .A2(new_n289_), .A3(new_n588_), .A4(new_n847_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n781_), .A2(new_n452_), .A3(new_n587_), .A4(new_n833_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n853_), .B1(new_n854_), .B2(new_n304_), .ZN(G1350gat));
  NAND3_X1  g654(.A1(new_n848_), .A2(new_n767_), .A3(new_n290_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n846_), .A2(new_n810_), .A3(new_n847_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(new_n305_), .ZN(G1351gat));
  NOR3_X1   g657(.A1(new_n662_), .A2(new_n516_), .A3(new_n514_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n781_), .A2(new_n699_), .A3(new_n859_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT125), .B(G197gat), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n781_), .A2(new_n699_), .A3(new_n859_), .A4(new_n861_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(G1352gat));
  NAND3_X1  g664(.A1(new_n781_), .A2(new_n792_), .A3(new_n859_), .ZN(new_n866_));
  XOR2_X1   g665(.A(KEYINPUT126), .B(G204gat), .Z(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n315_), .A2(KEYINPUT126), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n866_), .B2(new_n869_), .ZN(G1353gat));
  OAI211_X1 g669(.A(new_n587_), .B(new_n859_), .C1(new_n778_), .C2(new_n780_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n872_));
  AND2_X1   g671(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n871_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n871_), .A2(new_n872_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT127), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n871_), .A2(KEYINPUT127), .A3(new_n872_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n874_), .B1(new_n877_), .B2(new_n878_), .ZN(G1354gat));
  NAND3_X1  g678(.A1(new_n781_), .A2(new_n574_), .A3(new_n859_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(G218gat), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n568_), .A2(G218gat), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n781_), .A2(new_n859_), .A3(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n883_), .ZN(G1355gat));
endmodule


