//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 1 0 0 1 0 0 1 0 0 1 1 0 1 1 1 0 0 0 1 1 1 0 1 0 0 1 1 0 1 0 0 0 1 1 1 1 1 0 0 1 1 0 0 0 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n633_, new_n634_, new_n635_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n830_, new_n831_, new_n832_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n847_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n893_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_;
  XNOR2_X1  g000(.A(KEYINPUT73), .B(G15gat), .ZN(new_n202_));
  INV_X1    g001(.A(G22gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G1gat), .ZN(new_n205_));
  INV_X1    g004(.A(G8gat), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT14), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G1gat), .B(G8gat), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n209_), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G29gat), .B(G36gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G43gat), .B(G50gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n210_), .A2(new_n211_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n215_), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT76), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT76), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n212_), .A2(new_n220_), .A3(new_n215_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n216_), .B1(new_n219_), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G229gat), .A2(G233gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n215_), .B(KEYINPUT15), .ZN(new_n226_));
  AOI22_X1  g025(.A1(new_n221_), .A2(new_n219_), .B1(new_n217_), .B2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n225_), .B1(new_n224_), .B2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G113gat), .B(G141gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G169gat), .B(G197gat), .ZN(new_n230_));
  XOR2_X1   g029(.A(new_n229_), .B(new_n230_), .Z(new_n231_));
  NAND2_X1  g030(.A1(new_n228_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n231_), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n225_), .B(new_n233_), .C1(new_n224_), .C2(new_n227_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G120gat), .B(G148gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT5), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G176gat), .B(G204gat), .ZN(new_n238_));
  XOR2_X1   g037(.A(new_n237_), .B(new_n238_), .Z(new_n239_));
  XNOR2_X1  g038(.A(G57gat), .B(G64gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n240_), .A2(KEYINPUT11), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(KEYINPUT11), .ZN(new_n243_));
  XOR2_X1   g042(.A(G71gat), .B(G78gat), .Z(new_n244_));
  NAND3_X1  g043(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n245_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G99gat), .A2(G106gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT6), .ZN(new_n248_));
  INV_X1    g047(.A(G99gat), .ZN(new_n249_));
  INV_X1    g048(.A(G106gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(new_n250_), .A3(KEYINPUT65), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT7), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT7), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n253_), .A2(new_n249_), .A3(new_n250_), .A4(KEYINPUT65), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n248_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n255_));
  OR2_X1    g054(.A1(G85gat), .A2(G92gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G85gat), .A2(G92gat), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n255_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT8), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT9), .ZN(new_n262_));
  AND3_X1   g061(.A1(new_n257_), .A2(KEYINPUT64), .A3(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(KEYINPUT64), .B1(new_n257_), .B2(new_n262_), .ZN(new_n264_));
  OAI221_X1 g063(.A(new_n256_), .B1(new_n262_), .B2(new_n257_), .C1(new_n263_), .C2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT10), .B(G99gat), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n265_), .B(new_n248_), .C1(G106gat), .C2(new_n266_), .ZN(new_n267_));
  AND2_X1   g066(.A1(new_n261_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n255_), .A2(KEYINPUT8), .A3(new_n258_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n246_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(KEYINPUT66), .A2(KEYINPUT12), .ZN(new_n271_));
  AND2_X1   g070(.A1(KEYINPUT66), .A2(KEYINPUT12), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n270_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n273_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n246_), .A2(new_n269_), .A3(new_n267_), .A4(new_n261_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G230gat), .A2(G233gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT67), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT68), .B1(new_n274_), .B2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n277_), .B(KEYINPUT67), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT68), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n270_), .A2(new_n272_), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n281_), .A2(new_n282_), .A3(new_n273_), .A4(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n280_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n270_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n276_), .B1(new_n286_), .B2(new_n275_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n239_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n287_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n239_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n280_), .A2(new_n284_), .A3(new_n289_), .A4(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n288_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT13), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n292_), .A2(new_n293_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n297_), .A2(KEYINPUT69), .ZN(new_n298_));
  INV_X1    g097(.A(new_n296_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(new_n294_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT69), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n235_), .B1(new_n298_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(G169gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT22), .ZN(new_n305_));
  AOI21_X1  g104(.A(G176gat), .B1(new_n305_), .B2(KEYINPUT78), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT22), .B(G169gat), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n306_), .B1(KEYINPUT78), .B2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT79), .ZN(new_n309_));
  INV_X1    g108(.A(G183gat), .ZN(new_n310_));
  INV_X1    g109(.A(G190gat), .ZN(new_n311_));
  OR3_X1    g110(.A1(new_n310_), .A2(new_n311_), .A3(KEYINPUT23), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT23), .B1(new_n310_), .B2(new_n311_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(G183gat), .A2(G190gat), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  AOI22_X1  g115(.A1(new_n314_), .A2(new_n316_), .B1(G169gat), .B2(G176gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n309_), .A2(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(new_n313_), .B(KEYINPUT77), .Z(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n312_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT25), .B(G183gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT26), .B(G190gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT24), .ZN(new_n323_));
  NOR2_X1   g122(.A1(G169gat), .A2(G176gat), .ZN(new_n324_));
  AOI22_X1  g123(.A1(new_n321_), .A2(new_n322_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G169gat), .A2(G176gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT24), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n327_), .A2(new_n324_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n320_), .A2(new_n325_), .A3(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n318_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G197gat), .B(G204gat), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT21), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  OR2_X1    g132(.A1(G197gat), .A2(G204gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G197gat), .A2(G204gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(KEYINPUT21), .A3(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G211gat), .B(G218gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n333_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n336_), .A2(new_n337_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n330_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT20), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(G176gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n307_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(new_n326_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n346_), .B1(new_n320_), .B2(new_n316_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT93), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n324_), .B1(new_n327_), .B2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n349_), .B1(new_n348_), .B2(new_n327_), .ZN(new_n350_));
  AND3_X1   g149(.A1(new_n350_), .A2(new_n314_), .A3(new_n325_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n340_), .B1(new_n347_), .B2(new_n351_), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n352_), .A2(KEYINPUT94), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(KEYINPUT94), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n343_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G226gat), .A2(G233gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  XOR2_X1   g157(.A(new_n358_), .B(KEYINPUT92), .Z(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n342_), .B1(new_n330_), .B2(new_n340_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n347_), .A2(new_n351_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT88), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n340_), .B(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n361_), .A2(new_n365_), .ZN(new_n366_));
  OAI22_X1  g165(.A1(new_n355_), .A2(new_n360_), .B1(new_n358_), .B2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G8gat), .B(G36gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT18), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G64gat), .B(G92gat), .ZN(new_n370_));
  XOR2_X1   g169(.A(new_n369_), .B(new_n370_), .Z(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n367_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT27), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n352_), .B(KEYINPUT94), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n359_), .B1(new_n375_), .B2(new_n343_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n358_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n340_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n377_), .B1(new_n362_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(new_n361_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n376_), .A2(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n374_), .B1(new_n382_), .B2(new_n371_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n355_), .A2(new_n360_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(new_n371_), .A3(new_n380_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n372_), .B1(new_n376_), .B2(new_n381_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  AOI22_X1  g186(.A1(new_n373_), .A2(new_n383_), .B1(new_n387_), .B2(new_n374_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT4), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G155gat), .A2(G162gat), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT81), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(KEYINPUT81), .A2(G155gat), .A3(G162gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT1), .ZN(new_n395_));
  INV_X1    g194(.A(G155gat), .ZN(new_n396_));
  INV_X1    g195(.A(G162gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT1), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n392_), .A2(new_n399_), .A3(new_n393_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n395_), .A2(new_n398_), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(G141gat), .ZN(new_n402_));
  INV_X1    g201(.A(G148gat), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(G141gat), .A2(G148gat), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n401_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT83), .ZN(new_n408_));
  AND3_X1   g207(.A1(KEYINPUT81), .A2(G155gat), .A3(G162gat), .ZN(new_n409_));
  AOI21_X1  g208(.A(KEYINPUT81), .B1(G155gat), .B2(G162gat), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n398_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT82), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(KEYINPUT82), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n402_), .A2(new_n403_), .A3(KEYINPUT3), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT3), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n419_), .B1(G141gat), .B2(G148gat), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n417_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n421_));
  AOI211_X1 g220(.A(new_n408_), .B(new_n411_), .C1(new_n416_), .C2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n418_), .A2(new_n420_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n417_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n423_), .A2(new_n424_), .A3(new_n414_), .A4(new_n415_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n411_), .ZN(new_n426_));
  AOI21_X1  g225(.A(KEYINPUT83), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n407_), .B1(new_n422_), .B2(new_n427_), .ZN(new_n428_));
  XOR2_X1   g227(.A(G127gat), .B(G134gat), .Z(new_n429_));
  XNOR2_X1  g228(.A(G113gat), .B(G120gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n428_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n428_), .A2(new_n431_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(KEYINPUT95), .A3(new_n433_), .ZN(new_n434_));
  OR3_X1    g233(.A1(new_n428_), .A2(KEYINPUT95), .A3(new_n431_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n389_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n428_), .A2(new_n389_), .A3(new_n431_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G225gat), .A2(G233gat), .ZN(new_n438_));
  XOR2_X1   g237(.A(new_n438_), .B(KEYINPUT96), .Z(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  OR3_X1    g239(.A1(new_n436_), .A2(KEYINPUT97), .A3(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT97), .B1(new_n436_), .B2(new_n440_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n434_), .A2(new_n435_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n438_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n441_), .A2(new_n442_), .A3(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G1gat), .B(G29gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(G85gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(KEYINPUT0), .B(G57gat), .ZN(new_n448_));
  XOR2_X1   g247(.A(new_n447_), .B(new_n448_), .Z(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n445_), .A2(new_n450_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n441_), .A2(new_n449_), .A3(new_n442_), .A4(new_n444_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G71gat), .B(G99gat), .ZN(new_n453_));
  INV_X1    g252(.A(G43gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n330_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n455_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n318_), .A2(new_n329_), .A3(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G227gat), .A2(G233gat), .ZN(new_n459_));
  XOR2_X1   g258(.A(new_n459_), .B(G15gat), .Z(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT30), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT31), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n456_), .A2(new_n458_), .A3(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n462_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT80), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n456_), .A2(new_n458_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n462_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT80), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n469_), .A2(new_n470_), .A3(new_n463_), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n466_), .A2(new_n471_), .A3(new_n431_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n431_), .B1(new_n466_), .B2(new_n471_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n451_), .A2(new_n452_), .A3(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G78gat), .B(G106gat), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G228gat), .A2(G233gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n428_), .A2(KEYINPUT29), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n364_), .B1(new_n479_), .B2(KEYINPUT87), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT87), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n428_), .A2(new_n481_), .A3(KEYINPUT29), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n478_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT86), .ZN(new_n484_));
  INV_X1    g283(.A(new_n406_), .ZN(new_n485_));
  AOI22_X1  g284(.A1(new_n394_), .A2(KEYINPUT1), .B1(new_n396_), .B2(new_n397_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n485_), .B1(new_n486_), .B2(new_n400_), .ZN(new_n487_));
  NOR3_X1   g286(.A1(new_n419_), .A2(G141gat), .A3(G148gat), .ZN(new_n488_));
  AOI21_X1  g287(.A(KEYINPUT3), .B1(new_n402_), .B2(new_n403_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n424_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n414_), .A2(new_n415_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n426_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(new_n408_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n425_), .A2(KEYINPUT83), .A3(new_n426_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n487_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT29), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n484_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n428_), .A2(KEYINPUT86), .A3(KEYINPUT29), .ZN(new_n498_));
  INV_X1    g297(.A(new_n478_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n378_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n497_), .A2(new_n498_), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n477_), .B1(new_n483_), .B2(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT87), .B1(new_n495_), .B2(new_n496_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n364_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(new_n482_), .A3(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(new_n499_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n507_), .A2(new_n501_), .A3(new_n476_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n503_), .A2(KEYINPUT85), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT89), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n495_), .A2(new_n496_), .ZN(new_n511_));
  XOR2_X1   g310(.A(KEYINPUT84), .B(KEYINPUT28), .Z(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G22gat), .B(G50gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT89), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n503_), .A2(new_n516_), .A3(new_n508_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n510_), .A2(new_n515_), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT90), .ZN(new_n519_));
  INV_X1    g318(.A(new_n515_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n520_), .A2(new_n509_), .A3(KEYINPUT89), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n518_), .A2(new_n519_), .A3(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n519_), .B1(new_n518_), .B2(new_n521_), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n388_), .B(new_n475_), .C1(new_n522_), .C2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT100), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n509_), .A2(KEYINPUT89), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n517_), .A2(new_n515_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n521_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT90), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n518_), .A2(new_n519_), .A3(new_n521_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n532_), .A2(KEYINPUT100), .A3(new_n388_), .A4(new_n475_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n522_), .A2(new_n523_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n451_), .A2(new_n452_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(new_n388_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n474_), .B1(new_n534_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n436_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n437_), .A2(new_n438_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n449_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n443_), .B(KEYINPUT98), .Z(new_n542_));
  INV_X1    g341(.A(new_n439_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n541_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n387_), .B1(new_n544_), .B2(KEYINPUT99), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT33), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n452_), .A2(new_n546_), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n441_), .A2(new_n444_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n548_), .A2(KEYINPUT33), .A3(new_n449_), .A4(new_n442_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT99), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n550_), .B(new_n541_), .C1(new_n542_), .C2(new_n543_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n545_), .A2(new_n547_), .A3(new_n549_), .A4(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n367_), .A2(KEYINPUT32), .A3(new_n371_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n371_), .A2(KEYINPUT32), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n382_), .A2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n535_), .A2(new_n553_), .A3(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n532_), .A2(new_n552_), .A3(new_n556_), .ZN(new_n557_));
  AOI22_X1  g356(.A1(new_n526_), .A2(new_n533_), .B1(new_n538_), .B2(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n303_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n268_), .A2(new_n269_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(new_n226_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G232gat), .A2(G233gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT34), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n563_), .A2(KEYINPUT35), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n268_), .A2(new_n269_), .A3(new_n215_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n561_), .A2(new_n564_), .A3(new_n565_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n563_), .A2(KEYINPUT35), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G190gat), .B(G218gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT70), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT71), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G134gat), .B(G162gat), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n571_), .B(new_n573_), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n574_), .A2(KEYINPUT36), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n568_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT36), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n574_), .B(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n568_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n580_), .A2(KEYINPUT37), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT37), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n578_), .B(KEYINPUT72), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n568_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n582_), .B1(new_n584_), .B2(new_n576_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n581_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT74), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G231gat), .A2(G233gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n217_), .B(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(new_n246_), .ZN(new_n590_));
  XOR2_X1   g389(.A(G127gat), .B(G155gat), .Z(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT16), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G183gat), .B(G211gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT17), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n590_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n594_), .A2(new_n595_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n590_), .A2(new_n596_), .A3(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n587_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n599_), .A2(new_n587_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n586_), .A2(new_n603_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT75), .Z(new_n605_));
  NAND2_X1  g404(.A1(new_n559_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n607_), .A2(new_n205_), .A3(new_n535_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT38), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n303_), .A2(new_n603_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n580_), .B(KEYINPUT101), .Z(new_n612_));
  NOR2_X1   g411(.A1(new_n558_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(G1gat), .B1(new_n614_), .B2(new_n536_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n608_), .A2(new_n609_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n610_), .A2(new_n615_), .A3(new_n616_), .ZN(G1324gat));
  NAND2_X1  g416(.A1(new_n383_), .A2(new_n373_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n387_), .A2(new_n374_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n607_), .A2(new_n206_), .A3(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n611_), .A2(new_n613_), .A3(new_n620_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n622_), .A2(new_n623_), .A3(G8gat), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n623_), .B1(new_n622_), .B2(G8gat), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n621_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g426(.A(new_n474_), .ZN(new_n628_));
  OAI21_X1  g427(.A(G15gat), .B1(new_n614_), .B2(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT41), .ZN(new_n630_));
  NOR3_X1   g429(.A1(new_n606_), .A2(G15gat), .A3(new_n628_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n630_), .A2(new_n631_), .ZN(G1326gat));
  OAI21_X1  g431(.A(G22gat), .B1(new_n614_), .B2(new_n532_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT42), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n607_), .A2(new_n203_), .A3(new_n534_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(G1327gat));
  INV_X1    g435(.A(new_n580_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n603_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n559_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(G29gat), .B1(new_n641_), .B2(new_n535_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT44), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT43), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n526_), .A2(new_n533_), .ZN(new_n645_));
  OAI211_X1 g444(.A(new_n530_), .B(new_n531_), .C1(new_n620_), .C2(new_n535_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n557_), .A2(new_n646_), .A3(new_n628_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n644_), .B1(new_n648_), .B2(new_n586_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n586_), .ZN(new_n650_));
  AOI211_X1 g449(.A(KEYINPUT43), .B(new_n650_), .C1(new_n645_), .C2(new_n647_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n649_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n303_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(new_n603_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n643_), .B1(new_n652_), .B2(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(KEYINPUT43), .B1(new_n558_), .B2(new_n650_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n648_), .A2(new_n644_), .A3(new_n586_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n658_), .A2(KEYINPUT44), .A3(new_n603_), .A4(new_n653_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n655_), .A2(new_n659_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n535_), .A2(G29gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n642_), .B1(new_n660_), .B2(new_n661_), .ZN(G1328gat));
  NOR2_X1   g461(.A1(new_n388_), .A2(G36gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n559_), .A2(new_n639_), .A3(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT45), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n655_), .A2(new_n620_), .A3(new_n659_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n666_), .B1(new_n667_), .B2(G36gat), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT46), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n668_), .A2(KEYINPUT102), .A3(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n669_), .A2(KEYINPUT102), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n669_), .A2(KEYINPUT102), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n668_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n670_), .A2(new_n673_), .ZN(G1329gat));
  NOR2_X1   g473(.A1(new_n628_), .A2(new_n454_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n655_), .A2(new_n659_), .A3(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT103), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT103), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n655_), .A2(new_n659_), .A3(new_n678_), .A4(new_n675_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n454_), .B1(new_n640_), .B2(new_n628_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n677_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g481(.A(G50gat), .B1(new_n641_), .B2(new_n534_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n534_), .A2(G50gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n660_), .B2(new_n684_), .ZN(G1331gat));
  NOR3_X1   g484(.A1(new_n298_), .A2(new_n302_), .A3(new_n235_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n687_), .A2(new_n603_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n688_), .A2(new_n535_), .A3(new_n613_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(G57gat), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n687_), .A2(new_n558_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(new_n605_), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n536_), .A2(G57gat), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n690_), .B1(new_n692_), .B2(new_n693_), .ZN(G1332gat));
  OR3_X1    g493(.A1(new_n692_), .A2(G64gat), .A3(new_n388_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n688_), .A2(new_n620_), .A3(new_n613_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(G64gat), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n697_), .A2(KEYINPUT48), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n697_), .A2(KEYINPUT48), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n695_), .B1(new_n698_), .B2(new_n699_), .ZN(G1333gat));
  OR3_X1    g499(.A1(new_n692_), .A2(G71gat), .A3(new_n628_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n688_), .A2(new_n474_), .A3(new_n613_), .ZN(new_n702_));
  XOR2_X1   g501(.A(KEYINPUT104), .B(KEYINPUT49), .Z(new_n703_));
  AND3_X1   g502(.A1(new_n702_), .A2(G71gat), .A3(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n702_), .B2(G71gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n701_), .B1(new_n704_), .B2(new_n705_), .ZN(G1334gat));
  OR3_X1    g505(.A1(new_n692_), .A2(G78gat), .A3(new_n532_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n688_), .A2(new_n534_), .A3(new_n613_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(KEYINPUT105), .B(KEYINPUT50), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n708_), .A2(G78gat), .A3(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n708_), .B2(G78gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n710_), .B2(new_n711_), .ZN(G1335gat));
  NOR3_X1   g511(.A1(new_n687_), .A2(new_n558_), .A3(new_n638_), .ZN(new_n713_));
  AOI21_X1  g512(.A(G85gat), .B1(new_n713_), .B2(new_n535_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT106), .Z(new_n715_));
  NOR4_X1   g514(.A1(new_n298_), .A2(new_n302_), .A3(new_n602_), .A4(new_n235_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n658_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n658_), .A2(KEYINPUT107), .A3(new_n716_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(G85gat), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n536_), .A2(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n715_), .B1(new_n721_), .B2(new_n723_), .ZN(G1336gat));
  AOI21_X1  g523(.A(G92gat), .B1(new_n713_), .B2(new_n620_), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n725_), .A2(KEYINPUT108), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n719_), .A2(G92gat), .A3(new_n620_), .A4(new_n720_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(KEYINPUT108), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n726_), .A2(new_n727_), .A3(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT109), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n729_), .B(new_n730_), .ZN(G1337gat));
  OAI21_X1  g530(.A(G99gat), .B1(new_n717_), .B2(new_n628_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n713_), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n628_), .A2(new_n266_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n732_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g535(.A1(new_n713_), .A2(new_n250_), .A3(new_n534_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT111), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n738_), .A2(KEYINPUT52), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n534_), .B(new_n716_), .C1(new_n649_), .C2(new_n651_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT110), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n658_), .A2(new_n742_), .A3(new_n534_), .A4(new_n716_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n250_), .B1(new_n738_), .B2(KEYINPUT52), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n739_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n739_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n745_), .ZN(new_n748_));
  AOI211_X1 g547(.A(new_n747_), .B(new_n748_), .C1(new_n741_), .C2(new_n743_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n737_), .B1(new_n746_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT53), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT53), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n752_), .B(new_n737_), .C1(new_n746_), .C2(new_n749_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(G1339gat));
  NOR3_X1   g553(.A1(new_n586_), .A2(new_n603_), .A3(new_n235_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT54), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n755_), .A2(new_n756_), .A3(new_n297_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n755_), .B2(new_n297_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n222_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n231_), .B1(new_n760_), .B2(new_n223_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n227_), .A2(new_n224_), .ZN(new_n762_));
  AOI22_X1  g561(.A1(new_n228_), .A2(new_n231_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n763_), .A2(new_n291_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT56), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n274_), .A2(new_n279_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n276_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n283_), .A2(new_n275_), .A3(new_n273_), .ZN(new_n768_));
  AOI22_X1  g567(.A1(new_n766_), .A2(KEYINPUT55), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n280_), .A2(new_n284_), .A3(new_n770_), .ZN(new_n771_));
  AOI211_X1 g570(.A(new_n765_), .B(new_n290_), .C1(new_n769_), .C2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n769_), .A2(new_n771_), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT56), .B1(new_n773_), .B2(new_n239_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n764_), .B1(new_n772_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT58), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n764_), .B(KEYINPUT58), .C1(new_n772_), .C2(new_n774_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n777_), .A2(new_n586_), .A3(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT113), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT57), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n292_), .A2(new_n763_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n774_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n773_), .A2(KEYINPUT56), .A3(new_n239_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n783_), .A2(KEYINPUT112), .A3(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n235_), .A2(new_n291_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n772_), .B2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n782_), .B1(new_n785_), .B2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n781_), .B1(new_n789_), .B2(new_n637_), .ZN(new_n790_));
  NOR3_X1   g589(.A1(new_n774_), .A2(new_n772_), .A3(new_n787_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n235_), .B(new_n291_), .C1(new_n784_), .C2(KEYINPUT112), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  OAI211_X1 g592(.A(KEYINPUT57), .B(new_n580_), .C1(new_n793_), .C2(new_n782_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT113), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n777_), .A2(new_n795_), .A3(new_n586_), .A4(new_n778_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n780_), .A2(new_n790_), .A3(new_n794_), .A4(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n759_), .B1(new_n797_), .B2(new_n603_), .ZN(new_n798_));
  NOR4_X1   g597(.A1(new_n534_), .A2(new_n536_), .A3(new_n620_), .A4(new_n628_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n798_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(G113gat), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(new_n802_), .A3(new_n235_), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT59), .B1(new_n798_), .B2(new_n800_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n790_), .A2(new_n794_), .A3(new_n779_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n603_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n759_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT59), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(new_n809_), .A3(new_n799_), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n804_), .A2(KEYINPUT114), .A3(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT114), .B1(new_n804_), .B2(new_n810_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n235_), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n811_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n803_), .B1(new_n814_), .B2(new_n802_), .ZN(G1340gat));
  NOR2_X1   g614(.A1(new_n298_), .A2(new_n302_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n804_), .A2(new_n810_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(G120gat), .ZN(new_n818_));
  INV_X1    g617(.A(new_n801_), .ZN(new_n819_));
  INV_X1    g618(.A(G120gat), .ZN(new_n820_));
  INV_X1    g619(.A(new_n816_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n820_), .B1(new_n821_), .B2(KEYINPUT60), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n822_), .B1(KEYINPUT60), .B2(new_n820_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n818_), .B1(new_n819_), .B2(new_n823_), .ZN(G1341gat));
  AOI21_X1  g623(.A(G127gat), .B1(new_n801_), .B2(new_n602_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(KEYINPUT115), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n811_), .A2(new_n812_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n602_), .A2(G127gat), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n826_), .B1(new_n827_), .B2(new_n828_), .ZN(G1342gat));
  AOI21_X1  g628(.A(G134gat), .B1(new_n801_), .B2(new_n612_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n586_), .A2(G134gat), .ZN(new_n831_));
  XOR2_X1   g630(.A(new_n831_), .B(KEYINPUT116), .Z(new_n832_));
  AOI21_X1  g631(.A(new_n830_), .B1(new_n827_), .B2(new_n832_), .ZN(G1343gat));
  NAND2_X1  g632(.A1(new_n797_), .A2(new_n603_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n807_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n532_), .A2(new_n474_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n837_), .A2(new_n535_), .A3(new_n388_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n835_), .A2(new_n836_), .A3(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT117), .B1(new_n798_), .B2(new_n838_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n235_), .ZN(new_n843_));
  XOR2_X1   g642(.A(KEYINPUT118), .B(G141gat), .Z(new_n844_));
  XNOR2_X1  g643(.A(new_n843_), .B(new_n844_), .ZN(G1344gat));
  NAND2_X1  g644(.A1(new_n842_), .A2(new_n816_), .ZN(new_n846_));
  XOR2_X1   g645(.A(KEYINPUT119), .B(G148gat), .Z(new_n847_));
  XNOR2_X1  g646(.A(new_n846_), .B(new_n847_), .ZN(G1345gat));
  AOI21_X1  g647(.A(new_n836_), .B1(new_n835_), .B2(new_n839_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n798_), .A2(KEYINPUT117), .A3(new_n838_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n602_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(KEYINPUT120), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n842_), .A2(new_n853_), .A3(new_n602_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(KEYINPUT61), .B(G155gat), .ZN(new_n855_));
  AND3_X1   g654(.A1(new_n852_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n855_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(G1346gat));
  INV_X1    g657(.A(new_n842_), .ZN(new_n859_));
  OAI21_X1  g658(.A(G162gat), .B1(new_n859_), .B2(new_n650_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n842_), .A2(new_n397_), .A3(new_n612_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1347gat));
  AOI21_X1  g661(.A(new_n304_), .B1(KEYINPUT122), .B2(KEYINPUT62), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n534_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n536_), .A2(new_n620_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n628_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n865_), .A2(new_n235_), .A3(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n865_), .A2(KEYINPUT121), .A3(new_n235_), .A4(new_n867_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n864_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(KEYINPUT122), .A2(KEYINPUT62), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n868_), .ZN(new_n875_));
  AOI22_X1  g674(.A1(new_n872_), .A2(new_n874_), .B1(new_n307_), .B2(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n874_), .B2(new_n872_), .ZN(G1348gat));
  NAND3_X1  g676(.A1(new_n865_), .A2(new_n816_), .A3(new_n867_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n798_), .A2(new_n534_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n867_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n821_), .A2(new_n344_), .A3(new_n880_), .ZN(new_n881_));
  AOI22_X1  g680(.A1(new_n878_), .A2(new_n344_), .B1(new_n879_), .B2(new_n881_), .ZN(G1349gat));
  NOR3_X1   g681(.A1(new_n880_), .A2(new_n603_), .A3(new_n321_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n865_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT123), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n880_), .A2(new_n603_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n879_), .A2(new_n885_), .A3(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n310_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n885_), .B1(new_n879_), .B2(new_n886_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n884_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT124), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1350gat));
  NAND2_X1  g691(.A1(new_n865_), .A2(new_n867_), .ZN(new_n893_));
  OAI21_X1  g692(.A(G190gat), .B1(new_n893_), .B2(new_n650_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n612_), .A2(new_n322_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n893_), .B2(new_n895_), .ZN(G1351gat));
  NOR4_X1   g695(.A1(new_n798_), .A2(new_n532_), .A3(new_n474_), .A4(new_n866_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n235_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g698(.A(KEYINPUT125), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n900_), .A2(G204gat), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n901_), .B1(new_n897_), .B2(new_n816_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n900_), .A2(G204gat), .ZN(new_n903_));
  XOR2_X1   g702(.A(new_n903_), .B(KEYINPUT126), .Z(new_n904_));
  XNOR2_X1  g703(.A(new_n902_), .B(new_n904_), .ZN(G1353gat));
  AOI21_X1  g704(.A(new_n603_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n897_), .A2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(KEYINPUT127), .ZN(new_n908_));
  NOR2_X1   g707(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT127), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n897_), .A2(new_n910_), .A3(new_n906_), .ZN(new_n911_));
  AND3_X1   g710(.A1(new_n908_), .A2(new_n909_), .A3(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n909_), .B1(new_n908_), .B2(new_n911_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1354gat));
  INV_X1    g713(.A(G218gat), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n897_), .A2(new_n915_), .A3(new_n612_), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n897_), .A2(new_n586_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(new_n915_), .ZN(G1355gat));
endmodule


