//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n769_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n921_, new_n922_, new_n923_,
    new_n925_, new_n926_, new_n928_, new_n929_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_;
  XOR2_X1   g000(.A(G127gat), .B(G155gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G183gat), .B(G211gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XOR2_X1   g005(.A(KEYINPUT75), .B(KEYINPUT17), .Z(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT76), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G15gat), .B(G22gat), .ZN(new_n210_));
  INV_X1    g009(.A(G1gat), .ZN(new_n211_));
  INV_X1    g010(.A(G8gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT14), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G1gat), .B(G8gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G231gat), .A2(G233gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n216_), .B(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G57gat), .B(G64gat), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n219_), .A2(KEYINPUT11), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(KEYINPUT11), .ZN(new_n221_));
  XOR2_X1   g020(.A(G71gat), .B(G78gat), .Z(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n221_), .A2(new_n222_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n218_), .B(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n209_), .A2(new_n227_), .ZN(new_n228_));
  XOR2_X1   g027(.A(new_n228_), .B(KEYINPUT77), .Z(new_n229_));
  XNOR2_X1  g028(.A(new_n206_), .B(KEYINPUT78), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n227_), .B1(new_n231_), .B2(KEYINPUT17), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n232_), .B1(KEYINPUT17), .B2(new_n231_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n229_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT23), .ZN(new_n236_));
  INV_X1    g035(.A(G183gat), .ZN(new_n237_));
  INV_X1    g036(.A(G190gat), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n236_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n239_), .B(new_n240_), .C1(G183gat), .C2(G190gat), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G169gat), .A2(G176gat), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(G176gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT83), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT83), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(G176gat), .ZN(new_n248_));
  INV_X1    g047(.A(G169gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT22), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT22), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(G169gat), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n246_), .A2(new_n248_), .A3(new_n250_), .A4(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n244_), .B1(new_n253_), .B2(KEYINPUT84), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n246_), .A2(new_n248_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT22), .B(G169gat), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT84), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n254_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT85), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n254_), .A2(KEYINPUT85), .A3(new_n258_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n242_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(KEYINPUT82), .A2(G190gat), .ZN(new_n264_));
  XOR2_X1   g063(.A(new_n264_), .B(KEYINPUT26), .Z(new_n265_));
  INV_X1    g064(.A(KEYINPUT25), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(G183gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT81), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n237_), .A2(KEYINPUT25), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n267_), .A2(KEYINPUT81), .ZN(new_n270_));
  AND4_X1   g069(.A1(new_n265_), .A2(new_n268_), .A3(new_n269_), .A4(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n244_), .A2(new_n272_), .ZN(new_n273_));
  OR3_X1    g072(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n274_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n275_));
  NOR3_X1   g074(.A1(new_n271_), .A2(new_n273_), .A3(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n263_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G227gat), .A2(G233gat), .ZN(new_n278_));
  INV_X1    g077(.A(G15gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n277_), .B(new_n280_), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n281_), .B(KEYINPUT31), .Z(new_n282_));
  XNOR2_X1  g081(.A(G71gat), .B(G99gat), .ZN(new_n283_));
  INV_X1    g082(.A(G43gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT86), .B(KEYINPUT30), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XOR2_X1   g086(.A(G127gat), .B(G134gat), .Z(new_n288_));
  XNOR2_X1  g087(.A(G113gat), .B(G120gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n287_), .B(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n282_), .B(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT91), .ZN(new_n293_));
  AOI21_X1  g092(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT89), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT3), .ZN(new_n298_));
  NOR3_X1   g097(.A1(new_n298_), .A2(G141gat), .A3(G148gat), .ZN(new_n299_));
  INV_X1    g098(.A(G141gat), .ZN(new_n300_));
  INV_X1    g099(.A(G148gat), .ZN(new_n301_));
  AOI21_X1  g100(.A(KEYINPUT3), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n297_), .B1(new_n299_), .B2(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT90), .B1(new_n296_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G141gat), .A2(G148gat), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT2), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n295_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n294_), .A2(KEYINPUT89), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n297_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(G141gat), .A2(G148gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT3), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n298_), .B1(G141gat), .B2(G148gat), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n311_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT90), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n310_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n304_), .A2(new_n317_), .A3(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n318_), .B1(new_n320_), .B2(KEYINPUT1), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT87), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  OAI211_X1 g125(.A(KEYINPUT87), .B(new_n318_), .C1(new_n320_), .C2(KEYINPUT1), .ZN(new_n327_));
  OR3_X1    g126(.A1(new_n318_), .A2(KEYINPUT88), .A3(KEYINPUT1), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT88), .B1(new_n318_), .B2(KEYINPUT1), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n326_), .A2(new_n327_), .A3(new_n328_), .A4(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n305_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n331_), .A2(new_n312_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n322_), .A2(new_n323_), .A3(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT28), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT28), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n322_), .A2(new_n336_), .A3(new_n323_), .A4(new_n333_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G22gat), .B(G50gat), .ZN(new_n338_));
  AND3_X1   g137(.A1(new_n335_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n338_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n293_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n338_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n321_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n310_), .A2(new_n315_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n343_), .B1(new_n344_), .B2(KEYINPUT90), .ZN(new_n345_));
  AOI22_X1  g144(.A1(new_n345_), .A2(new_n317_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n336_), .B1(new_n346_), .B2(new_n323_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n337_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n342_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n335_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(KEYINPUT91), .A3(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n322_), .A2(new_n333_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT29), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G228gat), .A2(G233gat), .ZN(new_n354_));
  INV_X1    g153(.A(G204gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(G197gat), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT92), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  OR2_X1    g157(.A1(new_n355_), .A2(G197gat), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n355_), .A2(KEYINPUT92), .A3(G197gat), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n358_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT21), .ZN(new_n362_));
  INV_X1    g161(.A(G218gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(G211gat), .ZN(new_n364_));
  INV_X1    g163(.A(G211gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(G218gat), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n362_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n361_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT93), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n361_), .A2(new_n367_), .A3(KEYINPUT93), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n361_), .A2(KEYINPUT21), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n364_), .A2(new_n366_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n359_), .A2(new_n356_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n374_), .B1(new_n375_), .B2(KEYINPUT21), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n373_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n372_), .A2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n353_), .A2(new_n354_), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n354_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n323_), .B1(new_n322_), .B2(new_n333_), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n370_), .A2(new_n371_), .B1(new_n373_), .B2(new_n376_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n380_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G78gat), .B(G106gat), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n379_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n384_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n354_), .B1(new_n353_), .B2(new_n378_), .ZN(new_n387_));
  NOR3_X1   g186(.A1(new_n381_), .A2(new_n380_), .A3(new_n382_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n386_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n341_), .A2(new_n351_), .A3(new_n385_), .A4(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT94), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n387_), .A2(new_n388_), .A3(new_n386_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n384_), .B1(new_n379_), .B2(new_n383_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT94), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n394_), .A2(new_n395_), .A3(new_n351_), .A4(new_n341_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n391_), .A2(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n386_), .A2(KEYINPUT95), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n379_), .A2(new_n383_), .A3(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(new_n350_), .A3(new_n349_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n399_), .B1(new_n379_), .B2(new_n383_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n397_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n352_), .A2(new_n290_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n290_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n322_), .A2(new_n333_), .A3(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n406_), .A2(KEYINPUT98), .A3(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT98), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n346_), .A2(new_n410_), .A3(new_n407_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n409_), .A2(KEYINPUT4), .A3(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT4), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n406_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G225gat), .A2(G233gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT99), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G1gat), .B(G29gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(G85gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT0), .B(G57gat), .ZN(new_n421_));
  XOR2_X1   g220(.A(new_n420_), .B(new_n421_), .Z(new_n422_));
  AOI21_X1  g221(.A(new_n417_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n418_), .A2(new_n422_), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n422_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n417_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n427_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n426_), .B1(new_n428_), .B2(new_n423_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n425_), .A2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n275_), .B(KEYINPUT96), .ZN(new_n431_));
  AND2_X1   g230(.A1(new_n267_), .A2(new_n269_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT26), .B(G190gat), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n273_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n244_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n435_));
  AOI22_X1  g234(.A1(new_n431_), .A2(new_n434_), .B1(new_n241_), .B2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT20), .B1(new_n436_), .B2(new_n382_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n437_), .B1(new_n277_), .B2(new_n382_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G226gat), .A2(G233gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT19), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n438_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n262_), .ZN(new_n443_));
  AOI21_X1  g242(.A(KEYINPUT85), .B1(new_n254_), .B2(new_n258_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n241_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  OR3_X1    g244(.A1(new_n271_), .A2(new_n273_), .A3(new_n275_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n382_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n275_), .A2(KEYINPUT96), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n275_), .A2(KEYINPUT96), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n434_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n435_), .A2(new_n241_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT20), .B1(new_n378_), .B2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n440_), .B1(new_n447_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n442_), .A2(new_n454_), .ZN(new_n455_));
  XOR2_X1   g254(.A(G8gat), .B(G36gat), .Z(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G64gat), .B(G92gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n455_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT20), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n463_), .B1(new_n436_), .B2(new_n382_), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n441_), .B(new_n464_), .C1(new_n277_), .C2(new_n382_), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n465_), .B(new_n460_), .C1(new_n438_), .C2(new_n441_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n462_), .A2(KEYINPUT27), .A3(new_n466_), .ZN(new_n467_));
  NOR3_X1   g266(.A1(new_n447_), .A2(new_n453_), .A3(new_n440_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n445_), .A2(new_n446_), .A3(new_n382_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n463_), .B1(new_n378_), .B2(new_n452_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n441_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n461_), .B1(new_n468_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(new_n466_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT27), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n467_), .A2(new_n475_), .ZN(new_n476_));
  NOR4_X1   g275(.A1(new_n292_), .A2(new_n405_), .A3(new_n430_), .A4(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n403_), .B1(new_n391_), .B2(new_n396_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n423_), .B1(new_n415_), .B2(new_n417_), .ZN(new_n479_));
  AOI21_X1  g278(.A(KEYINPUT33), .B1(new_n479_), .B2(new_n422_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT33), .ZN(new_n481_));
  NOR4_X1   g280(.A1(new_n428_), .A2(new_n481_), .A3(new_n426_), .A4(new_n423_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n409_), .A2(new_n411_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(new_n417_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n426_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n417_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n466_), .B(new_n472_), .C1(new_n485_), .C2(new_n486_), .ZN(new_n487_));
  NOR3_X1   g286(.A1(new_n480_), .A2(new_n482_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n460_), .A2(KEYINPUT32), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n455_), .A2(new_n490_), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n465_), .B(new_n489_), .C1(new_n438_), .C2(new_n441_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n493_), .B1(new_n429_), .B2(new_n425_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n478_), .B1(new_n488_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT100), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n476_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n430_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n498_), .A2(new_n405_), .A3(new_n499_), .ZN(new_n500_));
  OAI211_X1 g299(.A(KEYINPUT100), .B(new_n478_), .C1(new_n488_), .C2(new_n494_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n497_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n477_), .B1(new_n502_), .B2(new_n292_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G29gat), .B(G36gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G43gat), .B(G50gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT15), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(new_n216_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n506_), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n216_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G229gat), .A2(G233gat), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n508_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n216_), .B(new_n509_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n511_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n512_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT80), .ZN(new_n517_));
  XOR2_X1   g316(.A(G113gat), .B(G141gat), .Z(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT79), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G169gat), .B(G197gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n517_), .B(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n503_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT13), .ZN(new_n526_));
  INV_X1    g325(.A(G230gat), .ZN(new_n527_));
  INV_X1    g326(.A(G233gat), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT8), .ZN(new_n530_));
  NOR2_X1   g329(.A1(G99gat), .A2(G106gat), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT7), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT6), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n535_), .B1(G99gat), .B2(G106gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G99gat), .A2(G106gat), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n537_), .A2(KEYINPUT6), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n533_), .B(new_n534_), .C1(new_n536_), .C2(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(G85gat), .B(G92gat), .Z(new_n540_));
  AOI21_X1  g339(.A(new_n530_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n530_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n533_), .A2(new_n534_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n537_), .A2(KEYINPUT6), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n535_), .A2(G99gat), .A3(G106gat), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n545_), .A2(new_n546_), .A3(KEYINPUT65), .ZN(new_n547_));
  AOI21_X1  g346(.A(KEYINPUT65), .B1(new_n545_), .B2(new_n546_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n544_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n542_), .B1(new_n549_), .B2(KEYINPUT66), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT65), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n551_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n545_), .A2(new_n546_), .A3(KEYINPUT65), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n543_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT66), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n541_), .B1(new_n550_), .B2(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(KEYINPUT10), .B(G99gat), .Z(new_n558_));
  INV_X1    g357(.A(G106gat), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n540_), .A2(KEYINPUT9), .ZN(new_n561_));
  XNOR2_X1  g360(.A(KEYINPUT64), .B(G85gat), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT9), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n562_), .A2(new_n563_), .A3(G92gat), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n560_), .A2(new_n561_), .A3(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n547_), .A2(new_n548_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT67), .B1(new_n557_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n541_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n542_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n570_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n549_), .A2(KEYINPUT66), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n569_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT67), .ZN(new_n574_));
  INV_X1    g373(.A(new_n567_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n568_), .A2(new_n576_), .A3(new_n225_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT68), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n568_), .A2(new_n576_), .A3(KEYINPUT68), .A4(new_n225_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n225_), .B1(new_n568_), .B2(new_n576_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n529_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n529_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n577_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NOR3_X1   g385(.A1(new_n557_), .A2(KEYINPUT67), .A3(new_n567_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n574_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n226_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT12), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n573_), .A2(new_n575_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n592_), .A2(KEYINPUT12), .A3(new_n226_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n586_), .A2(new_n591_), .A3(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(G120gat), .B(G148gat), .Z(new_n595_));
  XNOR2_X1  g394(.A(G176gat), .B(G204gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n583_), .A2(new_n594_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n600_), .B1(new_n583_), .B2(new_n594_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n526_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n603_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n605_), .A2(KEYINPUT13), .A3(new_n601_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n568_), .A2(new_n576_), .A3(new_n506_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT71), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n557_), .A2(new_n567_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n507_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n610_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n592_), .A2(KEYINPUT71), .A3(new_n507_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n609_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G232gat), .A2(G233gat), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT34), .Z(new_n617_));
  XNOR2_X1  g416(.A(KEYINPUT70), .B(KEYINPUT35), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n617_), .A2(new_n618_), .ZN(new_n620_));
  AOI211_X1 g419(.A(new_n619_), .B(new_n620_), .C1(new_n592_), .C2(new_n507_), .ZN(new_n621_));
  AOI22_X1  g420(.A1(new_n615_), .A2(new_n619_), .B1(new_n609_), .B2(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(G190gat), .B(G218gat), .Z(new_n623_));
  XNOR2_X1  g422(.A(G134gat), .B(G162gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT36), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT72), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n622_), .A2(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n625_), .B(new_n626_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n629_), .B1(new_n622_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT73), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n632_), .B1(new_n622_), .B2(new_n630_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n631_), .A2(KEYINPUT37), .A3(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT37), .ZN(new_n635_));
  OAI221_X1 g434(.A(new_n629_), .B1(new_n632_), .B2(new_n635_), .C1(new_n622_), .C2(new_n630_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  AND4_X1   g436(.A1(new_n235_), .A2(new_n525_), .A3(new_n608_), .A4(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n638_), .A2(new_n211_), .A3(new_n430_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT38), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n608_), .A2(new_n523_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n631_), .ZN(new_n642_));
  NOR4_X1   g441(.A1(new_n503_), .A2(new_n641_), .A3(new_n642_), .A4(new_n234_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n211_), .B1(new_n643_), .B2(new_n430_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT101), .Z(new_n645_));
  NAND2_X1  g444(.A1(new_n640_), .A2(new_n645_), .ZN(G1324gat));
  NAND3_X1  g445(.A1(new_n638_), .A2(new_n212_), .A3(new_n476_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n643_), .A2(new_n476_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT39), .ZN(new_n649_));
  AND4_X1   g448(.A1(KEYINPUT102), .A2(new_n648_), .A3(new_n649_), .A4(G8gat), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n212_), .B1(new_n651_), .B2(KEYINPUT39), .ZN(new_n652_));
  AOI22_X1  g451(.A1(new_n648_), .A2(new_n652_), .B1(KEYINPUT102), .B2(new_n649_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n647_), .B1(new_n650_), .B2(new_n653_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g454(.A(new_n292_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n279_), .B1(new_n643_), .B2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT41), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n638_), .A2(new_n279_), .A3(new_n656_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1326gat));
  INV_X1    g459(.A(G22gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n661_), .B1(new_n643_), .B2(new_n405_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT42), .Z(new_n663_));
  NOR2_X1   g462(.A1(new_n478_), .A2(G22gat), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT103), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n638_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n663_), .A2(new_n666_), .ZN(G1327gat));
  NAND2_X1  g466(.A1(new_n642_), .A2(new_n234_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n607_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n525_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(G29gat), .B1(new_n671_), .B2(new_n430_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n501_), .A2(new_n500_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n425_), .A2(new_n481_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n485_), .A2(new_n486_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n676_), .A2(new_n473_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n479_), .A2(KEYINPUT33), .A3(new_n422_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n675_), .A2(new_n677_), .A3(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n430_), .A2(new_n492_), .A3(new_n491_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT100), .B1(new_n681_), .B2(new_n478_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n292_), .B1(new_n674_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n477_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n637_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n673_), .B(KEYINPUT43), .C1(new_n685_), .C2(new_n686_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n641_), .A2(new_n235_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n637_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n478_), .A2(new_n476_), .A3(new_n430_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n405_), .B1(new_n680_), .B2(new_n679_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n691_), .B2(KEYINPUT100), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n656_), .B1(new_n692_), .B2(new_n497_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n689_), .B1(new_n693_), .B2(new_n477_), .ZN(new_n694_));
  AOI21_X1  g493(.A(KEYINPUT105), .B1(new_n694_), .B2(KEYINPUT104), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT43), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n696_), .B1(new_n685_), .B2(new_n673_), .ZN(new_n697_));
  OAI211_X1 g496(.A(new_n687_), .B(new_n688_), .C1(new_n695_), .C2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n673_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n694_), .A2(KEYINPUT105), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n701_), .A2(new_n702_), .A3(new_n696_), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n703_), .A2(KEYINPUT44), .A3(new_n687_), .A4(new_n688_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n700_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n430_), .A2(G29gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n672_), .B1(new_n706_), .B2(new_n707_), .ZN(G1328gat));
  NAND3_X1  g507(.A1(new_n700_), .A2(new_n476_), .A3(new_n704_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(G36gat), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n670_), .A2(G36gat), .A3(new_n498_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n711_), .B(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n710_), .A2(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n710_), .B(new_n713_), .C1(KEYINPUT107), .C2(KEYINPUT46), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1329gat));
  OAI21_X1  g517(.A(new_n284_), .B1(new_n670_), .B2(new_n292_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n656_), .A2(G43gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n705_), .B2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g521(.A(G50gat), .B1(new_n671_), .B2(new_n405_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n405_), .A2(G50gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n723_), .B1(new_n706_), .B2(new_n724_), .ZN(G1331gat));
  NOR2_X1   g524(.A1(new_n234_), .A2(new_n523_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n607_), .A2(new_n726_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n503_), .A2(new_n642_), .A3(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n728_), .A2(G57gat), .A3(new_n430_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n730_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n503_), .A2(new_n523_), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n608_), .A2(new_n234_), .A3(new_n689_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n735_), .A2(new_n499_), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n731_), .B(new_n732_), .C1(G57gat), .C2(new_n736_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT109), .Z(G1332gat));
  INV_X1    g537(.A(G64gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n728_), .B2(new_n476_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT48), .Z(new_n741_));
  INV_X1    g540(.A(new_n735_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n742_), .A2(new_n739_), .A3(new_n476_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1333gat));
  INV_X1    g543(.A(G71gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n728_), .B2(new_n656_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n746_), .B(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n742_), .A2(new_n745_), .A3(new_n656_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1334gat));
  INV_X1    g549(.A(G78gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n728_), .B2(new_n405_), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n752_), .B(KEYINPUT50), .Z(new_n753_));
  NAND3_X1  g552(.A1(new_n742_), .A2(new_n751_), .A3(new_n405_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1335gat));
  NOR2_X1   g554(.A1(new_n608_), .A2(new_n668_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n733_), .A2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT111), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n733_), .A2(KEYINPUT111), .A3(new_n756_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(G85gat), .B1(new_n761_), .B2(new_n430_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n607_), .A2(new_n234_), .A3(new_n524_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT112), .Z(new_n764_));
  OAI211_X1 g563(.A(new_n687_), .B(new_n764_), .C1(new_n695_), .C2(new_n697_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT113), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n430_), .A2(new_n562_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n762_), .B1(new_n766_), .B2(new_n767_), .ZN(G1336gat));
  INV_X1    g567(.A(G92gat), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n761_), .A2(new_n769_), .A3(new_n476_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n766_), .A2(new_n476_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(new_n769_), .ZN(G1337gat));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n656_), .A2(new_n558_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n760_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT111), .B1(new_n733_), .B2(new_n756_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n776_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT114), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n761_), .A2(KEYINPUT114), .A3(new_n776_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n775_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n773_), .A2(new_n774_), .ZN(new_n784_));
  OAI21_X1  g583(.A(G99gat), .B1(new_n765_), .B2(new_n292_), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n783_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n784_), .B1(new_n783_), .B2(new_n785_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n786_), .A2(new_n787_), .ZN(G1338gat));
  XNOR2_X1  g587(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n789_));
  OAI21_X1  g588(.A(G106gat), .B1(new_n765_), .B2(new_n478_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT52), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n792_), .B(G106gat), .C1(new_n765_), .C2(new_n478_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(new_n794_));
  AOI211_X1 g593(.A(G106gat), .B(new_n478_), .C1(new_n759_), .C2(new_n760_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n789_), .B1(new_n794_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n789_), .ZN(new_n798_));
  AOI211_X1 g597(.A(new_n795_), .B(new_n798_), .C1(new_n791_), .C2(new_n793_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n797_), .A2(new_n799_), .ZN(G1339gat));
  INV_X1    g599(.A(KEYINPUT123), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n508_), .A2(new_n510_), .A3(new_n514_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n513_), .A2(new_n511_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n521_), .A3(new_n803_), .ZN(new_n804_));
  XOR2_X1   g603(.A(new_n804_), .B(KEYINPUT119), .Z(new_n805_));
  NOR2_X1   g604(.A1(new_n516_), .A2(new_n521_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n807_), .A2(new_n601_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n593_), .B1(new_n582_), .B2(KEYINPUT12), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n529_), .B1(new_n581_), .B2(new_n809_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n586_), .A2(new_n591_), .A3(KEYINPUT55), .A4(new_n593_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n812_), .B1(new_n809_), .B2(new_n585_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n810_), .A2(new_n811_), .A3(new_n813_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n814_), .A2(KEYINPUT56), .A3(new_n599_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT56), .B1(new_n814_), .B2(new_n599_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n808_), .B(KEYINPUT58), .C1(new_n815_), .C2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n689_), .A2(new_n817_), .ZN(new_n818_));
  XOR2_X1   g617(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n814_), .A2(new_n599_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT56), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n814_), .A2(KEYINPUT56), .A3(new_n599_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n820_), .B1(new_n825_), .B2(new_n808_), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT121), .B1(new_n818_), .B2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n808_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n819_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT121), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n829_), .A2(new_n830_), .A3(new_n689_), .A4(new_n817_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n827_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT122), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT57), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n642_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n601_), .A2(new_n523_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n836_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n807_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n838_), .B1(new_n605_), .B2(new_n601_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n835_), .B1(new_n837_), .B2(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n833_), .A2(new_n834_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n840_), .B(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n235_), .B1(new_n832_), .B2(new_n842_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n637_), .A2(new_n606_), .A3(new_n604_), .A4(new_n726_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n845_), .B2(KEYINPUT54), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(KEYINPUT54), .ZN(new_n847_));
  XOR2_X1   g646(.A(new_n847_), .B(KEYINPUT118), .Z(new_n848_));
  XNOR2_X1  g647(.A(new_n846_), .B(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n801_), .B1(new_n843_), .B2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n841_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n840_), .B(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n827_), .A2(new_n831_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n234_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n855_), .A2(KEYINPUT123), .A3(new_n849_), .ZN(new_n856_));
  NOR4_X1   g655(.A1(new_n292_), .A2(new_n405_), .A3(new_n499_), .A4(new_n476_), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n851_), .A2(new_n856_), .A3(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(G113gat), .B1(new_n858_), .B2(new_n523_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n857_), .A2(new_n860_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n818_), .A2(new_n826_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n234_), .B1(new_n853_), .B2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n861_), .B1(new_n863_), .B2(new_n849_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n851_), .A2(new_n856_), .A3(new_n857_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(KEYINPUT59), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n524_), .A2(KEYINPUT124), .ZN(new_n867_));
  MUX2_X1   g666(.A(KEYINPUT124), .B(new_n867_), .S(G113gat), .Z(new_n868_));
  AOI21_X1  g667(.A(new_n859_), .B1(new_n866_), .B2(new_n868_), .ZN(G1340gat));
  INV_X1    g668(.A(G120gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n870_), .B1(new_n608_), .B2(KEYINPUT60), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n858_), .B(new_n871_), .C1(KEYINPUT60), .C2(new_n870_), .ZN(new_n872_));
  AND2_X1   g671(.A1(new_n866_), .A2(new_n607_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(new_n870_), .ZN(G1341gat));
  AOI21_X1  g673(.A(G127gat), .B1(new_n858_), .B2(new_n235_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n234_), .A2(KEYINPUT125), .ZN(new_n876_));
  MUX2_X1   g675(.A(KEYINPUT125), .B(new_n876_), .S(G127gat), .Z(new_n877_));
  AOI21_X1  g676(.A(new_n875_), .B1(new_n866_), .B2(new_n877_), .ZN(G1342gat));
  INV_X1    g677(.A(G134gat), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n637_), .A2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  AOI211_X1 g680(.A(new_n864_), .B(new_n881_), .C1(new_n865_), .C2(KEYINPUT59), .ZN(new_n882_));
  AOI21_X1  g681(.A(G134gat), .B1(new_n858_), .B2(new_n642_), .ZN(new_n883_));
  OAI21_X1  g682(.A(KEYINPUT126), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n866_), .A2(new_n880_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT126), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n879_), .B1(new_n865_), .B2(new_n631_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n885_), .A2(new_n886_), .A3(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n884_), .A2(new_n888_), .ZN(G1343gat));
  AND2_X1   g688(.A1(new_n851_), .A2(new_n856_), .ZN(new_n890_));
  NOR4_X1   g689(.A1(new_n656_), .A2(new_n499_), .A3(new_n478_), .A4(new_n476_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n893_), .A2(new_n300_), .A3(new_n523_), .ZN(new_n894_));
  OAI21_X1  g693(.A(G141gat), .B1(new_n892_), .B2(new_n524_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1344gat));
  NAND3_X1  g695(.A1(new_n893_), .A2(new_n301_), .A3(new_n607_), .ZN(new_n897_));
  OAI21_X1  g696(.A(G148gat), .B1(new_n892_), .B2(new_n608_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1345gat));
  XNOR2_X1  g698(.A(KEYINPUT61), .B(G155gat), .ZN(new_n900_));
  OR3_X1    g699(.A1(new_n892_), .A2(new_n234_), .A3(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n892_), .B2(new_n234_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1346gat));
  OAI21_X1  g702(.A(G162gat), .B1(new_n892_), .B2(new_n637_), .ZN(new_n904_));
  OR2_X1    g703(.A1(new_n631_), .A2(G162gat), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n892_), .B2(new_n905_), .ZN(G1347gat));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n498_), .A2(new_n430_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n656_), .A2(new_n908_), .ZN(new_n909_));
  AOI211_X1 g708(.A(new_n405_), .B(new_n909_), .C1(new_n863_), .C2(new_n849_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n523_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n907_), .B1(new_n912_), .B2(new_n249_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n256_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n911_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n913_), .A2(new_n914_), .A3(new_n915_), .ZN(G1348gat));
  AND2_X1   g715(.A1(new_n890_), .A2(new_n478_), .ZN(new_n917_));
  NOR3_X1   g716(.A1(new_n608_), .A2(new_n909_), .A3(new_n245_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n910_), .A2(new_n607_), .ZN(new_n919_));
  AOI22_X1  g718(.A1(new_n917_), .A2(new_n918_), .B1(new_n255_), .B2(new_n919_), .ZN(G1349gat));
  NOR2_X1   g719(.A1(new_n234_), .A2(new_n432_), .ZN(new_n921_));
  AND2_X1   g720(.A1(new_n910_), .A2(new_n921_), .ZN(new_n922_));
  NAND4_X1  g721(.A1(new_n917_), .A2(new_n656_), .A3(new_n235_), .A4(new_n908_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n922_), .B1(new_n923_), .B2(new_n237_), .ZN(G1350gat));
  NAND3_X1  g723(.A1(new_n910_), .A2(new_n433_), .A3(new_n642_), .ZN(new_n925_));
  AND2_X1   g724(.A1(new_n910_), .A2(new_n689_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n925_), .B1(new_n926_), .B2(new_n238_), .ZN(G1351gat));
  AND3_X1   g726(.A1(new_n908_), .A2(new_n405_), .A3(new_n292_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n890_), .A2(new_n523_), .A3(new_n928_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g729(.A1(new_n890_), .A2(new_n928_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n931_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(KEYINPUT127), .B(G204gat), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n932_), .A2(new_n607_), .A3(new_n933_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n933_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n935_), .B1(new_n931_), .B2(new_n608_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n934_), .A2(new_n936_), .ZN(G1353gat));
  NAND3_X1  g736(.A1(new_n890_), .A2(new_n235_), .A3(new_n928_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(KEYINPUT63), .B(G211gat), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n940_), .B1(new_n938_), .B2(new_n941_), .ZN(G1354gat));
  OAI21_X1  g741(.A(G218gat), .B1(new_n931_), .B2(new_n637_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n642_), .A2(new_n363_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n943_), .B1(new_n931_), .B2(new_n944_), .ZN(G1355gat));
endmodule


