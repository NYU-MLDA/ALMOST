//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 1 0 0 1 1 0 1 1 0 1 1 0 1 0 0 1 0 0 1 0 1 0 0 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n870_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n877_, new_n878_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_;
  XNOR2_X1  g000(.A(G85gat), .B(G92gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT6), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT66), .ZN(new_n206_));
  AOI211_X1 g005(.A(G99gat), .B(G106gat), .C1(KEYINPUT65), .C2(KEYINPUT7), .ZN(new_n207_));
  NOR2_X1   g006(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n203_), .B1(new_n206_), .B2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT8), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n202_), .A2(KEYINPUT8), .ZN(new_n212_));
  INV_X1    g011(.A(new_n205_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n212_), .B1(new_n209_), .B2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT10), .B(G99gat), .ZN(new_n217_));
  OAI22_X1  g016(.A1(new_n216_), .A2(new_n202_), .B1(new_n217_), .B2(G106gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G85gat), .ZN(new_n221_));
  INV_X1    g020(.A(G92gat), .ZN(new_n222_));
  NOR3_X1   g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  NOR3_X1   g022(.A1(new_n218_), .A2(new_n213_), .A3(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n215_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G43gat), .B(G50gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G29gat), .B(G36gat), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n229_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  XOR2_X1   g031(.A(new_n232_), .B(KEYINPUT15), .Z(new_n233_));
  NAND2_X1  g032(.A1(new_n226_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n215_), .A2(new_n225_), .A3(new_n230_), .A4(new_n231_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G232gat), .A2(G233gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT35), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n236_), .A2(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n239_), .A2(new_n240_), .ZN(new_n243_));
  NOR3_X1   g042(.A1(new_n235_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n235_), .A2(KEYINPUT71), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT72), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n242_), .A2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n236_), .A2(KEYINPUT72), .A3(new_n241_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT71), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n234_), .A2(new_n249_), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n245_), .A2(new_n247_), .A3(new_n248_), .A4(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n244_), .B1(new_n251_), .B2(new_n243_), .ZN(new_n252_));
  XOR2_X1   g051(.A(G190gat), .B(G218gat), .Z(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT73), .ZN(new_n254_));
  XOR2_X1   g053(.A(G134gat), .B(G162gat), .Z(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT36), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n252_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n256_), .B(new_n257_), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n259_), .B(KEYINPUT74), .C1(new_n252_), .C2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT37), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G15gat), .B(G22gat), .ZN(new_n263_));
  INV_X1    g062(.A(G1gat), .ZN(new_n264_));
  INV_X1    g063(.A(G8gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT14), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n263_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G1gat), .B(G8gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT75), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G57gat), .B(G64gat), .ZN(new_n271_));
  OR2_X1    g070(.A1(new_n271_), .A2(KEYINPUT11), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(KEYINPUT11), .ZN(new_n273_));
  XOR2_X1   g072(.A(G71gat), .B(G78gat), .Z(new_n274_));
  NAND3_X1  g073(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  OR2_X1    g074(.A1(new_n273_), .A2(new_n274_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n270_), .B(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G231gat), .A2(G233gat), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n280_), .B(KEYINPUT76), .Z(new_n281_));
  XNOR2_X1  g080(.A(new_n279_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G127gat), .B(G155gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT16), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G183gat), .B(G211gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n286_), .A2(KEYINPUT17), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n282_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(KEYINPUT17), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n282_), .A2(KEYINPUT77), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n262_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n226_), .A2(new_n278_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT12), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G230gat), .A2(G233gat), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n224_), .B1(new_n211_), .B2(new_n214_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(new_n277_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n226_), .A2(KEYINPUT12), .A3(new_n278_), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n297_), .A2(new_n298_), .A3(new_n300_), .A4(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n295_), .A2(new_n300_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n298_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G176gat), .B(G204gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT68), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G120gat), .B(G148gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n310_), .B(new_n311_), .Z(new_n312_));
  NAND2_X1  g111(.A1(new_n306_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n312_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n302_), .A2(new_n305_), .A3(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT69), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT13), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n313_), .A2(KEYINPUT69), .A3(new_n315_), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n318_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n319_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n294_), .A2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT78), .ZN(new_n326_));
  NOR3_X1   g125(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT24), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n328_), .B1(G169gat), .B2(G176gat), .ZN(new_n329_));
  INV_X1    g128(.A(G169gat), .ZN(new_n330_));
  INV_X1    g129(.A(G176gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n327_), .B1(new_n329_), .B2(new_n332_), .ZN(new_n333_));
  OR2_X1    g132(.A1(KEYINPUT79), .A2(KEYINPUT23), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G183gat), .A2(G190gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(KEYINPUT79), .A2(KEYINPUT23), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n334_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n335_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT23), .ZN(new_n339_));
  INV_X1    g138(.A(G183gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(KEYINPUT25), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT25), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(G183gat), .ZN(new_n343_));
  INV_X1    g142(.A(G190gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT26), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT26), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(G190gat), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n341_), .A2(new_n343_), .A3(new_n345_), .A4(new_n347_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n333_), .A2(new_n337_), .A3(new_n339_), .A4(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n330_), .A2(KEYINPUT22), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT22), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(G169gat), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n350_), .A2(new_n352_), .A3(new_n331_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n350_), .A2(new_n352_), .A3(KEYINPUT80), .A4(new_n331_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G169gat), .A2(G176gat), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n355_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n334_), .A2(new_n338_), .A3(new_n336_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n335_), .A2(KEYINPUT23), .ZN(new_n360_));
  AOI22_X1  g159(.A1(new_n359_), .A2(new_n360_), .B1(new_n340_), .B2(new_n344_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n349_), .B1(new_n358_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT81), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n349_), .B(KEYINPUT81), .C1(new_n358_), .C2(new_n361_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT30), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G15gat), .B(G43gat), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n368_), .B(KEYINPUT82), .Z(new_n369_));
  XOR2_X1   g168(.A(G71gat), .B(G99gat), .Z(new_n370_));
  NAND2_X1  g169(.A1(G227gat), .A2(G233gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n369_), .B(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n367_), .B(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT31), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G113gat), .B(G120gat), .ZN(new_n376_));
  INV_X1    g175(.A(G134gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(G127gat), .ZN(new_n378_));
  INV_X1    g177(.A(G127gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(G134gat), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n378_), .A2(new_n380_), .A3(KEYINPUT83), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(KEYINPUT83), .B1(new_n378_), .B2(new_n380_), .ZN(new_n383_));
  NOR3_X1   g182(.A1(new_n382_), .A2(new_n383_), .A3(KEYINPUT84), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT84), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n378_), .A2(new_n380_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT83), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n385_), .B1(new_n388_), .B2(new_n381_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n376_), .B1(new_n384_), .B2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT84), .B1(new_n382_), .B2(new_n383_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n388_), .A2(new_n385_), .A3(new_n381_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n376_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n391_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n390_), .A2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n375_), .B(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G8gat), .B(G36gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT18), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G64gat), .B(G92gat), .ZN(new_n400_));
  XOR2_X1   g199(.A(new_n399_), .B(new_n400_), .Z(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  OR2_X1    g201(.A1(G197gat), .A2(G204gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G197gat), .A2(G204gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT90), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT21), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  XOR2_X1   g207(.A(G211gat), .B(G218gat), .Z(new_n409_));
  NOR2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n406_), .A2(KEYINPUT21), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n407_), .B1(new_n405_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n405_), .A2(KEYINPUT91), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT91), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n403_), .A2(new_n415_), .A3(new_n404_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n409_), .A2(KEYINPUT21), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n413_), .A2(new_n419_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n337_), .B(new_n339_), .C1(G183gat), .C2(G190gat), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n421_), .A2(new_n353_), .A3(new_n357_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n359_), .A2(new_n360_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n423_), .A2(new_n348_), .A3(new_n333_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n420_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT20), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT93), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n429_), .B1(new_n366_), .B2(new_n420_), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n410_), .A2(new_n412_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n431_));
  AOI211_X1 g230(.A(KEYINPUT93), .B(new_n431_), .C1(new_n364_), .C2(new_n365_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n428_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G226gat), .A2(G233gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT19), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n364_), .A2(new_n365_), .A3(new_n431_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n427_), .B1(new_n420_), .B2(new_n425_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n435_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n437_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT97), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n402_), .B1(new_n436_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT99), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n439_), .B(new_n428_), .C1(new_n430_), .C2(new_n432_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n437_), .A2(new_n438_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n435_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n445_), .A2(new_n401_), .A3(new_n447_), .ZN(new_n448_));
  OAI211_X1 g247(.A(KEYINPUT99), .B(new_n402_), .C1(new_n436_), .C2(new_n441_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n444_), .A2(KEYINPUT27), .A3(new_n448_), .A4(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(G141gat), .A2(G148gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT3), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT3), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n453_), .B1(G141gat), .B2(G148gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G141gat), .A2(G148gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT2), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT2), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n458_), .A2(G141gat), .A3(G148gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n455_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G155gat), .A2(G162gat), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT86), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(KEYINPUT86), .A2(G155gat), .A3(G162gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  OR2_X1    g265(.A1(G155gat), .A2(G162gat), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n461_), .A2(KEYINPUT88), .A3(new_n466_), .A4(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT88), .ZN(new_n469_));
  AOI22_X1  g268(.A1(new_n454_), .A2(new_n452_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n466_), .A2(new_n467_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n469_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n468_), .A2(new_n472_), .ZN(new_n473_));
  AND3_X1   g272(.A1(KEYINPUT86), .A2(G155gat), .A3(G162gat), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT86), .B1(G155gat), .B2(G162gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT1), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT1), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n464_), .A2(new_n477_), .A3(new_n465_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n476_), .A2(new_n478_), .A3(new_n467_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT85), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n451_), .A2(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT85), .B1(G141gat), .B2(G148gat), .ZN(new_n482_));
  AOI22_X1  g281(.A1(new_n481_), .A2(new_n482_), .B1(G141gat), .B2(G148gat), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n479_), .A2(KEYINPUT87), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT87), .B1(new_n479_), .B2(new_n483_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n473_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  OR3_X1    g286(.A1(new_n487_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT28), .B1(new_n487_), .B2(KEYINPUT29), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G22gat), .B(G50gat), .Z(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n431_), .B1(new_n487_), .B2(KEYINPUT29), .ZN(new_n493_));
  NAND2_X1  g292(.A1(KEYINPUT89), .A2(G233gat), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(KEYINPUT89), .A2(G233gat), .ZN(new_n496_));
  OAI21_X1  g295(.A(G228gat), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  OR2_X1    g296(.A1(new_n493_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n493_), .A2(new_n497_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G78gat), .B(G106gat), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n498_), .A2(new_n499_), .A3(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT92), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n492_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n498_), .A2(new_n499_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(new_n500_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n504_), .A2(new_n502_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n502_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n508_), .A2(new_n492_), .A3(new_n503_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G225gat), .A2(G233gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n487_), .A2(new_n395_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT4), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n511_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n512_), .A2(KEYINPUT95), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT96), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n517_), .B1(new_n487_), .B2(new_n395_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n479_), .A2(new_n483_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT87), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  AOI22_X1  g320(.A1(new_n521_), .A2(new_n484_), .B1(new_n472_), .B2(new_n468_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n522_), .A2(KEYINPUT96), .A3(new_n394_), .A4(new_n390_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT95), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n487_), .A2(new_n524_), .A3(new_n395_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n516_), .A2(new_n518_), .A3(new_n523_), .A4(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n515_), .B1(new_n526_), .B2(new_n514_), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n523_), .A2(new_n518_), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n487_), .A2(new_n524_), .A3(new_n395_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n524_), .B1(new_n487_), .B2(new_n395_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n528_), .A2(new_n531_), .A3(new_n511_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G1gat), .B(G29gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT0), .ZN(new_n534_));
  INV_X1    g333(.A(G57gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(G85gat), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n527_), .A2(new_n532_), .A3(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n537_), .B1(new_n527_), .B2(new_n532_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(KEYINPUT100), .B(KEYINPUT27), .Z(new_n542_));
  AOI21_X1  g341(.A(new_n401_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT94), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n543_), .B1(new_n544_), .B2(new_n448_), .ZN(new_n545_));
  AOI211_X1 g344(.A(KEYINPUT94), .B(new_n401_), .C1(new_n445_), .C2(new_n447_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n542_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n450_), .A2(new_n510_), .A3(new_n541_), .A4(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n543_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n448_), .A2(new_n544_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n546_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n537_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n511_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n528_), .A2(new_n531_), .A3(KEYINPUT4), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n513_), .A2(new_n514_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n553_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n511_), .B1(new_n528_), .B2(new_n531_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n552_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n527_), .A2(KEYINPUT33), .A3(new_n532_), .A4(new_n537_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT33), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n538_), .A2(new_n560_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n551_), .A2(new_n558_), .A3(new_n559_), .A4(new_n561_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n401_), .A2(KEYINPUT32), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n563_), .B1(new_n436_), .B2(new_n441_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n445_), .A2(new_n447_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n565_), .A2(new_n563_), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n564_), .B(new_n566_), .C1(new_n539_), .C2(new_n540_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n510_), .B1(new_n562_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT98), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n548_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  AOI211_X1 g369(.A(KEYINPUT98), .B(new_n510_), .C1(new_n562_), .C2(new_n567_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n397_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n396_), .A2(new_n541_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n450_), .A2(new_n547_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n510_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n572_), .A2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n269_), .B(new_n232_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G229gat), .A2(G233gat), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n269_), .A2(new_n232_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n582_), .B1(new_n233_), .B2(new_n269_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n580_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n581_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(G113gat), .B(G141gat), .Z(new_n586_));
  XNOR2_X1  g385(.A(G169gat), .B(G197gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n585_), .A2(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n585_), .A2(new_n588_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n326_), .A2(new_n578_), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT101), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n594_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n541_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(new_n264_), .ZN(new_n599_));
  OR3_X1    g398(.A1(new_n597_), .A2(KEYINPUT38), .A3(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(KEYINPUT38), .B1(new_n597_), .B2(new_n599_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n573_), .A2(new_n576_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n558_), .A2(new_n561_), .A3(new_n559_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n550_), .A2(new_n549_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n546_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n567_), .B1(new_n604_), .B2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(new_n575_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(KEYINPUT98), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n568_), .A2(new_n569_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n610_), .A2(new_n611_), .A3(new_n548_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n603_), .B1(new_n612_), .B2(new_n397_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n259_), .B1(new_n252_), .B2(new_n260_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n324_), .A2(new_n591_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n616_), .A2(new_n617_), .A3(new_n293_), .ZN(new_n618_));
  OAI21_X1  g417(.A(G1gat), .B1(new_n618_), .B2(new_n541_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n602_), .A2(new_n619_), .ZN(G1324gat));
  INV_X1    g419(.A(new_n574_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n595_), .A2(new_n265_), .A3(new_n621_), .A4(new_n596_), .ZN(new_n622_));
  OAI21_X1  g421(.A(G8gat), .B1(new_n618_), .B2(new_n574_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT39), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT40), .Z(G1325gat));
  OR2_X1    g425(.A1(new_n397_), .A2(G15gat), .ZN(new_n627_));
  OR3_X1    g426(.A1(new_n597_), .A2(KEYINPUT102), .A3(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(KEYINPUT102), .B1(new_n597_), .B2(new_n627_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G15gat), .B1(new_n618_), .B2(new_n397_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT41), .Z(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(G1326gat));
  OAI21_X1  g432(.A(G22gat), .B1(new_n618_), .B2(new_n575_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT42), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n575_), .A2(G22gat), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT103), .Z(new_n637_));
  OAI21_X1  g436(.A(new_n635_), .B1(new_n597_), .B2(new_n637_), .ZN(G1327gat));
  NOR2_X1   g437(.A1(new_n293_), .A2(new_n614_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n617_), .A2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n640_), .A2(new_n613_), .ZN(new_n641_));
  AOI21_X1  g440(.A(G29gat), .B1(new_n641_), .B2(new_n598_), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n324_), .A2(new_n591_), .A3(new_n293_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT43), .ZN(new_n644_));
  INV_X1    g443(.A(new_n262_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n644_), .B1(new_n578_), .B2(new_n645_), .ZN(new_n646_));
  AOI211_X1 g445(.A(KEYINPUT43), .B(new_n262_), .C1(new_n572_), .C2(new_n577_), .ZN(new_n647_));
  OAI211_X1 g446(.A(KEYINPUT44), .B(new_n643_), .C1(new_n646_), .C2(new_n647_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n648_), .A2(G29gat), .A3(new_n598_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT44), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n646_), .A2(new_n647_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n643_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n650_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n642_), .B1(new_n649_), .B2(new_n653_), .ZN(G1328gat));
  INV_X1    g453(.A(KEYINPUT107), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT105), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n648_), .A2(new_n621_), .ZN(new_n657_));
  OAI21_X1  g456(.A(KEYINPUT43), .B1(new_n613_), .B2(new_n262_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n578_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(KEYINPUT44), .B1(new_n660_), .B2(new_n643_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G36gat), .B1(new_n657_), .B2(new_n661_), .ZN(new_n662_));
  XOR2_X1   g461(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n574_), .A2(G36gat), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n664_), .B1(new_n641_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n665_), .ZN(new_n667_));
  NOR4_X1   g466(.A1(new_n640_), .A2(new_n613_), .A3(new_n667_), .A4(new_n663_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n662_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT46), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n656_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  AOI211_X1 g472(.A(KEYINPUT105), .B(KEYINPUT46), .C1(new_n662_), .C2(new_n670_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n653_), .A2(new_n621_), .A3(new_n648_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n669_), .B1(new_n676_), .B2(G36gat), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n677_), .A2(KEYINPUT106), .A3(KEYINPUT46), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n662_), .A2(KEYINPUT46), .A3(new_n670_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT106), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n678_), .A2(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n655_), .B1(new_n675_), .B2(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n679_), .B(KEYINPUT106), .ZN(new_n684_));
  OAI21_X1  g483(.A(KEYINPUT105), .B1(new_n677_), .B2(KEYINPUT46), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n671_), .A2(new_n656_), .A3(new_n672_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n684_), .A2(new_n687_), .A3(KEYINPUT107), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n683_), .A2(new_n688_), .ZN(G1329gat));
  NAND3_X1  g488(.A1(new_n648_), .A2(G43gat), .A3(new_n396_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n641_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n691_), .A2(new_n397_), .ZN(new_n692_));
  OAI22_X1  g491(.A1(new_n690_), .A2(new_n661_), .B1(new_n692_), .B2(G43gat), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g493(.A1(new_n691_), .A2(G50gat), .A3(new_n575_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n648_), .A2(new_n510_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(new_n653_), .A3(KEYINPUT108), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(G50gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(KEYINPUT108), .B1(new_n696_), .B2(new_n653_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n695_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT109), .Z(G1331gat));
  NOR2_X1   g500(.A1(new_n323_), .A2(new_n592_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n616_), .A2(new_n293_), .A3(new_n702_), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n703_), .A2(new_n535_), .A3(new_n541_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT110), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n578_), .A2(new_n702_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n706_), .A2(new_n294_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n535_), .B1(new_n708_), .B2(new_n541_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n705_), .A2(new_n709_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT111), .Z(G1332gat));
  OAI21_X1  g510(.A(G64gat), .B1(new_n703_), .B2(new_n574_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT48), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n574_), .A2(G64gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n713_), .B1(new_n708_), .B2(new_n714_), .ZN(G1333gat));
  OAI21_X1  g514(.A(G71gat), .B1(new_n703_), .B2(new_n397_), .ZN(new_n716_));
  XOR2_X1   g515(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n717_));
  XNOR2_X1  g516(.A(new_n716_), .B(new_n717_), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n397_), .A2(G71gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n708_), .B2(new_n719_), .ZN(G1334gat));
  OAI21_X1  g519(.A(G78gat), .B1(new_n703_), .B2(new_n575_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT50), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n575_), .A2(G78gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(new_n708_), .B2(new_n723_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT113), .Z(G1335gat));
  INV_X1    g524(.A(new_n706_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(new_n639_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(G85gat), .B1(new_n728_), .B2(new_n598_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n702_), .A2(new_n292_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n651_), .A2(new_n730_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n541_), .A2(new_n221_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT114), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n729_), .B1(new_n731_), .B2(new_n733_), .ZN(G1336gat));
  NAND3_X1  g533(.A1(new_n728_), .A2(new_n222_), .A3(new_n621_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n651_), .A2(new_n574_), .A3(new_n730_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n735_), .B1(new_n736_), .B2(new_n222_), .ZN(G1337gat));
  NOR3_X1   g536(.A1(new_n727_), .A2(new_n217_), .A3(new_n397_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n731_), .A2(new_n396_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(G99gat), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g540(.A(G106gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n742_), .B1(new_n731_), .B2(new_n510_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT116), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n743_), .A2(KEYINPUT116), .A3(new_n744_), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n743_), .A2(new_n744_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n747_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n728_), .A2(new_n742_), .A3(new_n510_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT53), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT53), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n750_), .A2(new_n754_), .A3(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1339gat));
  NAND4_X1  g555(.A1(new_n396_), .A2(new_n574_), .A3(new_n598_), .A4(new_n575_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT57), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n583_), .B(KEYINPUT119), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(new_n584_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n588_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n589_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n318_), .A2(new_n320_), .A3(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n592_), .A2(new_n315_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n300_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n296_), .B2(new_n295_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n767_), .A2(KEYINPUT55), .A3(new_n298_), .A4(new_n301_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n302_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n297_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n304_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n768_), .A2(new_n770_), .A3(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT117), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n768_), .A2(new_n770_), .A3(KEYINPUT117), .A4(new_n772_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT118), .B1(new_n777_), .B2(new_n312_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n765_), .B1(new_n778_), .B2(KEYINPUT56), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT56), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n314_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n780_), .B1(new_n781_), .B2(KEYINPUT118), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n764_), .B1(new_n779_), .B2(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n758_), .B1(new_n783_), .B2(new_n615_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n777_), .A2(new_n312_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT118), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n785_), .A2(new_n786_), .A3(KEYINPUT56), .ZN(new_n787_));
  INV_X1    g586(.A(new_n765_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n782_), .A3(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n763_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n790_), .A2(KEYINPUT57), .A3(new_n614_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n762_), .A2(new_n315_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n792_), .B1(new_n781_), .B2(new_n780_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n793_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT58), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n793_), .B(KEYINPUT58), .C1(new_n780_), .C2(new_n781_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n645_), .A3(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n784_), .A2(new_n791_), .A3(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n292_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n262_), .A2(new_n591_), .A3(new_n323_), .A4(new_n293_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n801_), .B(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n757_), .B1(new_n800_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(G113gat), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n806_), .A3(new_n592_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n803_), .B1(new_n292_), .B2(new_n799_), .ZN(new_n808_));
  NOR3_X1   g607(.A1(new_n808_), .A2(KEYINPUT59), .A3(new_n757_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT120), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT59), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n810_), .B1(new_n805_), .B2(new_n811_), .ZN(new_n812_));
  OAI211_X1 g611(.A(KEYINPUT120), .B(KEYINPUT59), .C1(new_n808_), .C2(new_n757_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n809_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n814_), .A2(new_n592_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n807_), .B1(new_n815_), .B2(new_n806_), .ZN(G1340gat));
  AND2_X1   g615(.A1(new_n814_), .A2(new_n324_), .ZN(new_n817_));
  INV_X1    g616(.A(G120gat), .ZN(new_n818_));
  INV_X1    g617(.A(new_n805_), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n323_), .A2(KEYINPUT60), .A3(G120gat), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n820_), .B1(KEYINPUT60), .B2(G120gat), .ZN(new_n821_));
  OAI22_X1  g620(.A1(new_n817_), .A2(new_n818_), .B1(new_n819_), .B2(new_n821_), .ZN(G1341gat));
  NAND2_X1  g621(.A1(new_n293_), .A2(G127gat), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT121), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n814_), .A2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n379_), .B1(new_n819_), .B2(new_n292_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT122), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n825_), .A2(KEYINPUT122), .A3(new_n826_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(G1342gat));
  AOI21_X1  g630(.A(new_n377_), .B1(new_n814_), .B2(new_n645_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n805_), .A2(new_n377_), .A3(new_n615_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT123), .B1(new_n832_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT123), .ZN(new_n836_));
  AOI211_X1 g635(.A(new_n262_), .B(new_n809_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n836_), .B(new_n833_), .C1(new_n837_), .C2(new_n377_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n835_), .A2(new_n838_), .ZN(G1343gat));
  INV_X1    g638(.A(new_n808_), .ZN(new_n840_));
  NOR4_X1   g639(.A1(new_n621_), .A2(new_n396_), .A3(new_n541_), .A4(new_n575_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n592_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n324_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g646(.A(KEYINPUT124), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n843_), .A2(new_n848_), .A3(new_n293_), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT124), .B1(new_n842_), .B2(new_n292_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(KEYINPUT61), .B(G155gat), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n851_), .B(new_n852_), .ZN(G1346gat));
  NAND2_X1  g652(.A1(new_n843_), .A2(new_n615_), .ZN(new_n854_));
  INV_X1    g653(.A(G162gat), .ZN(new_n855_));
  AND3_X1   g654(.A1(new_n854_), .A2(KEYINPUT125), .A3(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(KEYINPUT125), .B1(new_n854_), .B2(new_n855_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n842_), .A2(new_n855_), .A3(new_n262_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n856_), .A2(new_n857_), .A3(new_n858_), .ZN(G1347gat));
  NOR3_X1   g658(.A1(new_n573_), .A2(new_n510_), .A3(new_n574_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n840_), .A2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n330_), .B1(new_n862_), .B2(new_n592_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT62), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n863_), .A2(new_n864_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n592_), .A2(new_n350_), .A3(new_n352_), .ZN(new_n867_));
  XOR2_X1   g666(.A(new_n867_), .B(KEYINPUT126), .Z(new_n868_));
  OAI22_X1  g667(.A1(new_n865_), .A2(new_n866_), .B1(new_n861_), .B2(new_n868_), .ZN(G1348gat));
  NOR2_X1   g668(.A1(new_n861_), .A2(new_n323_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(new_n331_), .ZN(G1349gat));
  NOR2_X1   g670(.A1(new_n861_), .A2(new_n292_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n340_), .A2(KEYINPUT127), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n872_), .A2(new_n341_), .A3(new_n343_), .A4(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(KEYINPUT127), .A2(G183gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n872_), .B2(new_n875_), .ZN(G1350gat));
  OAI21_X1  g675(.A(G190gat), .B1(new_n861_), .B2(new_n262_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n615_), .A2(new_n345_), .A3(new_n347_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n861_), .B2(new_n878_), .ZN(G1351gat));
  NAND3_X1  g678(.A1(new_n397_), .A2(new_n541_), .A3(new_n510_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n808_), .A2(new_n574_), .A3(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n592_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n324_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g684(.A(KEYINPUT63), .ZN(new_n886_));
  INV_X1    g685(.A(G211gat), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n881_), .B(new_n293_), .C1(new_n886_), .C2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n887_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1354gat));
  INV_X1    g689(.A(G218gat), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n881_), .A2(new_n891_), .A3(new_n615_), .ZN(new_n892_));
  AND2_X1   g691(.A1(new_n881_), .A2(new_n645_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n891_), .ZN(G1355gat));
endmodule


