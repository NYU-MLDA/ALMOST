//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1 0 0 0 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 0 1 1 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 1 1 1 0 1 1 1 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n903_, new_n904_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n934_, new_n935_,
    new_n936_, new_n938_, new_n939_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n946_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT23), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  OR2_X1    g003(.A1(G183gat), .A2(G190gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT80), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(G169gat), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n204_), .A2(new_n205_), .A3(KEYINPUT80), .A4(new_n206_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n209_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT26), .B(G190gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT79), .ZN(new_n215_));
  INV_X1    g014(.A(G183gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT25), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT25), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(KEYINPUT79), .A3(G183gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n214_), .A2(new_n217_), .A3(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(G169gat), .ZN(new_n223_));
  INV_X1    g022(.A(G176gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n222_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n204_), .A2(new_n206_), .ZN(new_n226_));
  NOR3_X1   g025(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n220_), .A2(new_n225_), .A3(new_n226_), .A4(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n213_), .A2(new_n229_), .A3(KEYINPUT81), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(KEYINPUT81), .B1(new_n213_), .B2(new_n229_), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT30), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n213_), .A2(new_n229_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT81), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT30), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n236_), .A2(new_n237_), .A3(new_n230_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT83), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n233_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n239_), .B1(new_n233_), .B2(new_n238_), .ZN(new_n242_));
  XOR2_X1   g041(.A(G15gat), .B(G71gat), .Z(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT82), .B(G43gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G227gat), .A2(G233gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(G99gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n245_), .B(new_n247_), .ZN(new_n248_));
  NOR3_X1   g047(.A1(new_n241_), .A2(new_n242_), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n242_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n248_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT85), .B1(new_n249_), .B2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n250_), .A2(new_n251_), .A3(new_n240_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT85), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n254_), .B(new_n255_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n256_));
  INV_X1    g055(.A(G113gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G127gat), .A2(G134gat), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(G127gat), .A2(G134gat), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT84), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(G127gat), .ZN(new_n262_));
  INV_X1    g061(.A(G134gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT84), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n264_), .A2(new_n265_), .A3(new_n258_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n257_), .B1(new_n261_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n261_), .A2(new_n266_), .A3(new_n257_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(G120gat), .A3(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(G120gat), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n261_), .A2(new_n266_), .A3(new_n257_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n271_), .B1(new_n272_), .B2(new_n267_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT31), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n253_), .A2(new_n256_), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n275_), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n277_), .B(KEYINPUT85), .C1(new_n249_), .C2(new_n252_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT29), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G155gat), .A2(G162gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT1), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT1), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n283_), .A2(G155gat), .A3(G162gat), .ZN(new_n284_));
  OR2_X1    g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n282_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(G141gat), .A2(G148gat), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n286_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT86), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n286_), .A2(KEYINPUT86), .A3(new_n288_), .A4(new_n289_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n287_), .B(KEYINPUT3), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n289_), .B(KEYINPUT2), .ZN(new_n296_));
  AOI22_X1  g095(.A1(new_n295_), .A2(new_n296_), .B1(G155gat), .B2(G162gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n285_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n280_), .B1(new_n294_), .B2(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G197gat), .B(G204gat), .Z(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT21), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G197gat), .B(G204gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT21), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G211gat), .B(G218gat), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n301_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n306_));
  OR3_X1    g105(.A1(new_n302_), .A2(new_n305_), .A3(new_n303_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G228gat), .A2(G233gat), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n310_), .A2(KEYINPUT88), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n310_), .A2(KEYINPUT88), .ZN(new_n312_));
  OAI22_X1  g111(.A1(new_n299_), .A2(new_n309_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G78gat), .B(G106gat), .ZN(new_n314_));
  XOR2_X1   g113(.A(new_n314_), .B(KEYINPUT89), .Z(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n310_), .A2(KEYINPUT88), .ZN(new_n317_));
  AOI22_X1  g116(.A1(new_n292_), .A2(new_n293_), .B1(new_n297_), .B2(new_n285_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n308_), .B(new_n317_), .C1(new_n318_), .C2(new_n280_), .ZN(new_n319_));
  AND3_X1   g118(.A1(new_n313_), .A2(new_n316_), .A3(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n316_), .B1(new_n313_), .B2(new_n319_), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT90), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n313_), .A2(new_n319_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n315_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT90), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n313_), .A2(new_n316_), .A3(new_n319_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n324_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n294_), .A2(new_n298_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n328_), .B1(new_n329_), .B2(KEYINPUT29), .ZN(new_n330_));
  XOR2_X1   g129(.A(G22gat), .B(G50gat), .Z(new_n331_));
  INV_X1    g130(.A(new_n328_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n318_), .A2(new_n280_), .A3(new_n332_), .ZN(new_n333_));
  AND3_X1   g132(.A1(new_n330_), .A2(new_n331_), .A3(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n331_), .B1(new_n330_), .B2(new_n333_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n322_), .A2(new_n327_), .A3(new_n337_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n336_), .B(KEYINPUT90), .C1(new_n321_), .C2(new_n320_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G8gat), .B(G36gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT18), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(G64gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(G92gat), .ZN(new_n344_));
  INV_X1    g143(.A(G64gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n342_), .B(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(G92gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n344_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G226gat), .A2(G233gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT19), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n236_), .A2(new_n230_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n308_), .B1(new_n207_), .B2(new_n211_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n221_), .B1(G169gat), .B2(G176gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n204_), .A2(new_n206_), .ZN(new_n356_));
  NOR3_X1   g155(.A1(new_n355_), .A2(new_n356_), .A3(new_n227_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT25), .B(G183gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n214_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  AOI22_X1  g159(.A1(new_n353_), .A2(new_n308_), .B1(new_n354_), .B2(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(KEYINPUT94), .B(KEYINPUT20), .Z(new_n362_));
  AOI21_X1  g161(.A(new_n352_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n236_), .A2(new_n309_), .A3(new_n230_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT91), .ZN(new_n365_));
  INV_X1    g164(.A(new_n207_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n210_), .B(new_n223_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n365_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n211_), .A2(KEYINPUT91), .A3(new_n207_), .ZN(new_n369_));
  AOI22_X1  g168(.A1(new_n368_), .A2(new_n369_), .B1(new_n357_), .B2(new_n359_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n364_), .B(KEYINPUT20), .C1(new_n309_), .C2(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n371_), .A2(new_n351_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n349_), .B1(new_n363_), .B2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n351_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT20), .ZN(new_n375_));
  AOI211_X1 g174(.A(new_n375_), .B(new_n351_), .C1(new_n370_), .C2(new_n309_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n353_), .A2(new_n308_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n349_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n374_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n373_), .A2(KEYINPUT27), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT27), .ZN(new_n382_));
  AOI221_X4 g181(.A(new_n349_), .B1(new_n376_), .B2(new_n377_), .C1(new_n371_), .C2(new_n351_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n379_), .B1(new_n374_), .B2(new_n378_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n382_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n381_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT92), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n274_), .A2(new_n329_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n387_), .B1(new_n388_), .B2(KEYINPUT4), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n270_), .A2(new_n294_), .A3(new_n273_), .A4(new_n298_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n388_), .A2(KEYINPUT4), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G225gat), .A2(G233gat), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT4), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n274_), .A2(new_n329_), .A3(KEYINPUT92), .A4(new_n394_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n389_), .A2(new_n391_), .A3(new_n393_), .A4(new_n395_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n388_), .A2(new_n390_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(new_n392_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G1gat), .B(G29gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(G85gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT0), .ZN(new_n401_));
  XOR2_X1   g200(.A(new_n401_), .B(G57gat), .Z(new_n402_));
  AND3_X1   g201(.A1(new_n396_), .A2(new_n398_), .A3(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n402_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NOR4_X1   g205(.A1(new_n279_), .A2(new_n340_), .A3(new_n386_), .A4(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n405_), .A2(new_n381_), .A3(new_n385_), .ZN(new_n409_));
  AOI22_X1  g208(.A1(new_n409_), .A2(new_n340_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n338_), .A2(new_n339_), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n379_), .A2(KEYINPUT32), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n363_), .B2(new_n372_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n374_), .A2(new_n378_), .ZN(new_n414_));
  OAI221_X1 g213(.A(new_n413_), .B1(new_n414_), .B2(new_n412_), .C1(new_n403_), .C2(new_n404_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n396_), .A2(new_n398_), .A3(KEYINPUT33), .A4(new_n402_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT93), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n383_), .A2(new_n384_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n396_), .A2(new_n398_), .A3(new_n402_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT33), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n402_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n389_), .A2(new_n391_), .A3(new_n392_), .A4(new_n395_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n397_), .A2(new_n393_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n419_), .A2(new_n422_), .A3(new_n426_), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n411_), .B(new_n415_), .C1(new_n418_), .C2(new_n427_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n410_), .A2(new_n428_), .A3(KEYINPUT95), .ZN(new_n429_));
  AOI21_X1  g228(.A(KEYINPUT95), .B1(new_n410_), .B2(new_n428_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n408_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  XOR2_X1   g230(.A(G71gat), .B(G78gat), .Z(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G57gat), .B(G64gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT11), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  OR2_X1    g235(.A1(new_n434_), .A2(KEYINPUT11), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n432_), .A2(KEYINPUT11), .A3(new_n434_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT66), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT64), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT10), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n442_), .A2(G99gat), .ZN(new_n443_));
  INV_X1    g242(.A(G99gat), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n444_), .A2(KEYINPUT10), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n441_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(KEYINPUT10), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n442_), .A2(G99gat), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(new_n448_), .A3(KEYINPUT64), .ZN(new_n449_));
  AOI21_X1  g248(.A(G106gat), .B1(new_n446_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT65), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n347_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT9), .ZN(new_n453_));
  NAND2_X1  g252(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n452_), .A2(new_n453_), .A3(G85gat), .A4(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G99gat), .A2(G106gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT6), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT6), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n458_), .A2(G99gat), .A3(G106gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G85gat), .B(G92gat), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n455_), .B(new_n460_), .C1(new_n453_), .C2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n440_), .B1(new_n450_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(G106gat), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n447_), .A2(new_n448_), .A3(KEYINPUT64), .ZN(new_n465_));
  AOI21_X1  g264(.A(KEYINPUT64), .B1(new_n447_), .B2(new_n448_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n464_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n461_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT9), .ZN(new_n469_));
  INV_X1    g268(.A(new_n454_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n453_), .A2(G85gat), .ZN(new_n473_));
  AOI22_X1  g272(.A1(new_n472_), .A2(new_n473_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n467_), .A2(KEYINPUT66), .A3(new_n469_), .A4(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n463_), .A2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT7), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(new_n444_), .A3(new_n464_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n460_), .A2(new_n477_), .A3(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT8), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n480_), .A2(new_n481_), .A3(new_n468_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n481_), .B1(new_n480_), .B2(new_n468_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n439_), .B1(new_n476_), .B2(new_n484_), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n457_), .A2(new_n459_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n479_), .A2(new_n477_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n468_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT8), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n480_), .A2(new_n481_), .A3(new_n468_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n439_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n491_), .A2(new_n492_), .A3(new_n463_), .A4(new_n475_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n485_), .A2(KEYINPUT12), .A3(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n491_), .A2(new_n463_), .A3(new_n475_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT12), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(new_n496_), .A3(new_n439_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n494_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(G230gat), .ZN(new_n499_));
  INV_X1    g298(.A(G233gat), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n498_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT67), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n485_), .A2(new_n504_), .A3(new_n493_), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n505_), .B(new_n501_), .C1(new_n504_), .C2(new_n485_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n503_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G120gat), .B(G148gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G176gat), .B(G204gat), .ZN(new_n511_));
  XOR2_X1   g310(.A(new_n510_), .B(new_n511_), .Z(new_n512_));
  NAND2_X1  g311(.A1(new_n507_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n512_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n503_), .A2(new_n506_), .A3(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT69), .ZN(new_n517_));
  OR2_X1    g316(.A1(new_n517_), .A2(KEYINPUT13), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(KEYINPUT13), .ZN(new_n520_));
  AND2_X1   g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n519_), .B1(new_n516_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G15gat), .B(G22gat), .ZN(new_n524_));
  INV_X1    g323(.A(G1gat), .ZN(new_n525_));
  INV_X1    g324(.A(G8gat), .ZN(new_n526_));
  OAI21_X1  g325(.A(KEYINPUT14), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G1gat), .B(G8gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(G29gat), .B(G36gat), .Z(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G43gat), .B(G50gat), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT72), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(G50gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(G43gat), .ZN(new_n538_));
  INV_X1    g337(.A(G43gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(G50gat), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n538_), .A2(new_n540_), .A3(new_n535_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n533_), .B1(new_n536_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n538_), .A2(new_n540_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT72), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n534_), .A2(new_n535_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(new_n545_), .A3(new_n532_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n542_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n531_), .A2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n530_), .A2(new_n546_), .A3(new_n542_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT78), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G229gat), .A2(G233gat), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n548_), .A2(KEYINPUT78), .A3(new_n549_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n552_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n542_), .A2(KEYINPUT15), .A3(new_n546_), .ZN(new_n557_));
  AOI21_X1  g356(.A(KEYINPUT15), .B1(new_n542_), .B2(new_n546_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(new_n530_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n560_), .A2(new_n553_), .A3(new_n548_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n556_), .A2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G113gat), .B(G141gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(new_n223_), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n564_), .B(G197gat), .Z(new_n565_));
  NAND2_X1  g364(.A1(new_n562_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n565_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n556_), .A2(new_n561_), .A3(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n523_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n431_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G190gat), .B(G218gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(G134gat), .ZN(new_n574_));
  INV_X1    g373(.A(G162gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT36), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n574_), .B(G162gat), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT36), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT73), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT73), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n578_), .A2(new_n580_), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G232gat), .A2(G233gat), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT70), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT34), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT35), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT71), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n559_), .A2(new_n495_), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n589_), .A2(KEYINPUT35), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n491_), .A2(new_n463_), .A3(new_n475_), .A4(new_n547_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n592_), .A2(new_n593_), .A3(new_n594_), .A4(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n593_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n592_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n585_), .A2(new_n596_), .A3(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT74), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n578_), .B1(new_n599_), .B2(new_n596_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT74), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n585_), .A2(new_n599_), .A3(new_n604_), .A4(new_n596_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n601_), .A2(new_n603_), .A3(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT37), .ZN(new_n607_));
  INV_X1    g406(.A(new_n581_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n599_), .A2(new_n608_), .A3(new_n596_), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n609_), .A2(KEYINPUT75), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n609_), .B1(new_n602_), .B2(KEYINPUT75), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT37), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n610_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n607_), .A2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G127gat), .B(G155gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT16), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(G183gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(G211gat), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(KEYINPUT17), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n619_), .B(KEYINPUT76), .Z(new_n620_));
  XNOR2_X1  g419(.A(new_n530_), .B(new_n439_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(G231gat), .A2(G233gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n620_), .A2(new_n623_), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n623_), .A2(KEYINPUT77), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n618_), .A2(KEYINPUT17), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n623_), .A2(KEYINPUT77), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n625_), .A2(new_n626_), .A3(new_n627_), .A4(new_n619_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n624_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n614_), .A2(new_n630_), .ZN(new_n631_));
  OR3_X1    g430(.A1(new_n572_), .A2(KEYINPUT96), .A3(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(KEYINPUT96), .B1(new_n572_), .B2(new_n631_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n634_), .A2(new_n525_), .A3(new_n406_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT38), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT97), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n410_), .A2(new_n428_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT95), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n410_), .A2(new_n428_), .A3(KEYINPUT95), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n407_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n610_), .A2(new_n611_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT99), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(KEYINPUT100), .B1(new_n644_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT100), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n431_), .A2(new_n649_), .A3(new_n646_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n522_), .A2(new_n630_), .A3(new_n569_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT98), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G1gat), .B1(new_n656_), .B2(new_n405_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n635_), .A2(new_n636_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT101), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n639_), .A2(new_n657_), .A3(new_n659_), .ZN(G1324gat));
  INV_X1    g459(.A(new_n386_), .ZN(new_n661_));
  AOI211_X1 g460(.A(new_n661_), .B(new_n654_), .C1(new_n648_), .C2(new_n650_), .ZN(new_n662_));
  OAI21_X1  g461(.A(KEYINPUT39), .B1(new_n662_), .B2(new_n526_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n654_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n651_), .A2(new_n386_), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT39), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n665_), .A2(new_n666_), .A3(G8gat), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n663_), .A2(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n661_), .A2(G8gat), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n632_), .A2(new_n633_), .A3(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n668_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT102), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT102), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n668_), .A2(new_n674_), .A3(new_n671_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n673_), .A2(KEYINPUT40), .A3(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT40), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n674_), .B1(new_n668_), .B2(new_n671_), .ZN(new_n678_));
  AOI211_X1 g477(.A(KEYINPUT102), .B(new_n670_), .C1(new_n663_), .C2(new_n667_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n677_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n676_), .A2(new_n680_), .ZN(G1325gat));
  INV_X1    g480(.A(G15gat), .ZN(new_n682_));
  INV_X1    g481(.A(new_n279_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n682_), .B1(new_n655_), .B2(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT41), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n634_), .A2(new_n682_), .A3(new_n683_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1326gat));
  INV_X1    g486(.A(G22gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n655_), .B2(new_n340_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT42), .Z(new_n690_));
  NAND3_X1  g489(.A1(new_n634_), .A2(new_n688_), .A3(new_n340_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1327gat));
  NAND2_X1  g491(.A1(new_n647_), .A2(new_n629_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n572_), .A2(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(G29gat), .B1(new_n694_), .B2(new_n406_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n571_), .A2(new_n629_), .ZN(new_n696_));
  OAI21_X1  g495(.A(KEYINPUT43), .B1(new_n644_), .B2(new_n614_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n607_), .A2(new_n613_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n431_), .A2(new_n698_), .A3(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n696_), .B1(new_n697_), .B2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(KEYINPUT44), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n702_), .A2(G29gat), .A3(new_n406_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n696_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n644_), .A2(KEYINPUT43), .A3(new_n614_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n698_), .B1(new_n431_), .B2(new_n699_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n704_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n695_), .B1(new_n703_), .B2(new_n709_), .ZN(G1328gat));
  INV_X1    g509(.A(G36gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n661_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n712_), .B2(new_n702_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n694_), .A2(new_n711_), .A3(new_n386_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT45), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n714_), .B(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(KEYINPUT103), .B1(new_n713_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT46), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n386_), .B1(new_n701_), .B2(KEYINPUT44), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n707_), .A2(new_n708_), .ZN(new_n720_));
  OAI21_X1  g519(.A(G36gat), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT103), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n714_), .B(KEYINPUT45), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n721_), .A2(new_n722_), .A3(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n717_), .A2(new_n718_), .A3(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n721_), .A2(KEYINPUT46), .A3(new_n723_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT104), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n717_), .A2(new_n724_), .A3(KEYINPUT104), .A4(new_n718_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1329gat));
  AND3_X1   g529(.A1(new_n709_), .A2(new_n702_), .A3(G43gat), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n694_), .A2(new_n683_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(KEYINPUT105), .B(G43gat), .ZN(new_n733_));
  AOI22_X1  g532(.A1(new_n731_), .A2(new_n683_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT47), .Z(G1330gat));
  NAND3_X1  g534(.A1(new_n709_), .A2(new_n702_), .A3(new_n340_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(G50gat), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT106), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n694_), .A2(new_n537_), .A3(new_n340_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1331gat));
  NOR2_X1   g539(.A1(new_n522_), .A2(new_n569_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n644_), .A2(new_n631_), .A3(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(G57gat), .B1(new_n743_), .B2(new_n406_), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n431_), .A2(new_n649_), .A3(new_n646_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n649_), .B1(new_n431_), .B2(new_n646_), .ZN(new_n746_));
  OAI211_X1 g545(.A(new_n630_), .B(new_n741_), .C1(new_n745_), .C2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n406_), .A2(G57gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n744_), .B1(new_n748_), .B2(new_n749_), .ZN(G1332gat));
  OAI21_X1  g549(.A(G64gat), .B1(new_n747_), .B2(new_n661_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT48), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n743_), .A2(new_n345_), .A3(new_n386_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(G1333gat));
  OAI21_X1  g553(.A(G71gat), .B1(new_n747_), .B2(new_n279_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT49), .ZN(new_n756_));
  INV_X1    g555(.A(G71gat), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n743_), .A2(new_n757_), .A3(new_n683_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1334gat));
  INV_X1    g558(.A(G78gat), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n743_), .A2(new_n760_), .A3(new_n340_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n651_), .A2(new_n630_), .A3(new_n340_), .A4(new_n741_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT108), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n762_), .A2(new_n763_), .A3(G78gat), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n763_), .B1(new_n762_), .B2(G78gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(KEYINPUT107), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(G78gat), .B1(new_n747_), .B2(new_n411_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT108), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT107), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n770_), .A3(new_n764_), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n767_), .A2(KEYINPUT50), .A3(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT50), .B1(new_n767_), .B2(new_n771_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n761_), .B1(new_n772_), .B2(new_n773_), .ZN(G1335gat));
  NOR3_X1   g573(.A1(new_n644_), .A2(new_n693_), .A3(new_n742_), .ZN(new_n775_));
  AOI21_X1  g574(.A(G85gat), .B1(new_n775_), .B2(new_n406_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n697_), .A2(new_n700_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n741_), .A2(new_n629_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT109), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n780_), .A2(KEYINPUT110), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n780_), .A2(KEYINPUT110), .ZN(new_n782_));
  OR2_X1    g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n406_), .A2(G85gat), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT111), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n776_), .B1(new_n783_), .B2(new_n785_), .ZN(G1336gat));
  OAI211_X1 g585(.A(new_n472_), .B(new_n386_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n775_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n347_), .B1(new_n788_), .B2(new_n661_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT112), .ZN(G1337gat));
  OAI21_X1  g590(.A(G99gat), .B1(new_n780_), .B2(new_n279_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n775_), .B(new_n683_), .C1(new_n466_), .C2(new_n465_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT113), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n792_), .A2(new_n796_), .A3(new_n793_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g598(.A1(new_n775_), .A2(new_n464_), .A3(new_n340_), .ZN(new_n800_));
  OAI21_X1  g599(.A(G106gat), .B1(new_n780_), .B2(new_n411_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n801_), .A2(KEYINPUT52), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n801_), .A2(KEYINPUT52), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n800_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g604(.A1(new_n522_), .A2(new_n614_), .A3(new_n630_), .A4(new_n570_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n806_), .A2(KEYINPUT114), .A3(KEYINPUT54), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT114), .B1(new_n806_), .B2(KEYINPUT54), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n806_), .A2(KEYINPUT54), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n807_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n515_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n498_), .A2(KEYINPUT115), .A3(KEYINPUT55), .A4(new_n501_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n813_), .B1(new_n501_), .B2(KEYINPUT115), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n814_), .B1(new_n498_), .B2(new_n502_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n813_), .B1(new_n494_), .B2(new_n497_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n512_), .B(new_n812_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT56), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT116), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n811_), .B1(new_n817_), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n498_), .A2(KEYINPUT55), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n501_), .B1(new_n494_), .B2(new_n497_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n822_), .B2(new_n814_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n819_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n823_), .A2(new_n512_), .A3(new_n812_), .A4(new_n824_), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n820_), .A2(new_n569_), .A3(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n552_), .A2(new_n553_), .A3(new_n555_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n560_), .A2(new_n554_), .A3(new_n548_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n827_), .A2(new_n565_), .A3(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n568_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n514_), .B1(new_n503_), .B2(new_n506_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n811_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT117), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n516_), .A2(new_n835_), .A3(new_n831_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n646_), .B1(new_n826_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  OR2_X1    g641(.A1(new_n838_), .A2(new_n839_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n823_), .A2(new_n818_), .A3(new_n512_), .A4(new_n812_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n844_), .A2(new_n515_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n830_), .B1(new_n817_), .B2(KEYINPUT56), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT58), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT119), .B1(new_n847_), .B2(new_n614_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n845_), .A2(KEYINPUT58), .A3(new_n846_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n817_), .A2(KEYINPUT56), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n850_), .A2(new_n515_), .A3(new_n831_), .A4(new_n844_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT58), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT119), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n699_), .A3(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n848_), .A2(new_n849_), .A3(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n838_), .A2(KEYINPUT118), .A3(new_n839_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n842_), .A2(new_n843_), .A3(new_n856_), .A4(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n810_), .B1(new_n858_), .B2(new_n629_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n386_), .A2(new_n405_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n683_), .A2(new_n860_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n859_), .A2(new_n340_), .A3(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(G113gat), .B1(new_n862_), .B2(new_n569_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n856_), .A2(new_n864_), .A3(new_n840_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n843_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n864_), .B1(new_n856_), .B2(new_n840_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n629_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n810_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n861_), .A2(KEYINPUT59), .A3(new_n340_), .ZN(new_n871_));
  AND2_X1   g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  OR3_X1    g671(.A1(new_n859_), .A2(new_n340_), .A3(new_n861_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT120), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n873_), .A2(new_n874_), .A3(KEYINPUT59), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT120), .B1(new_n862_), .B2(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n872_), .B1(new_n875_), .B2(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n570_), .A2(new_n257_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n863_), .B1(new_n878_), .B2(new_n879_), .ZN(G1340gat));
  OAI21_X1  g679(.A(new_n271_), .B1(new_n522_), .B2(KEYINPUT60), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n862_), .B(new_n881_), .C1(KEYINPUT60), .C2(new_n271_), .ZN(new_n882_));
  AOI211_X1 g681(.A(new_n522_), .B(new_n872_), .C1(new_n875_), .C2(new_n877_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(new_n271_), .ZN(G1341gat));
  AOI21_X1  g683(.A(G127gat), .B1(new_n862_), .B2(new_n630_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n262_), .B1(new_n630_), .B2(new_n886_), .ZN(new_n887_));
  AOI211_X1 g686(.A(new_n872_), .B(new_n887_), .C1(new_n875_), .C2(new_n877_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n262_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n885_), .B1(new_n888_), .B2(new_n889_), .ZN(G1342gat));
  AOI21_X1  g689(.A(G134gat), .B1(new_n862_), .B2(new_n647_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n614_), .A2(new_n263_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n893_), .B1(new_n878_), .B2(new_n894_), .ZN(G1343gat));
  NAND3_X1  g694(.A1(new_n860_), .A2(new_n340_), .A3(new_n279_), .ZN(new_n896_));
  XOR2_X1   g695(.A(new_n896_), .B(KEYINPUT124), .Z(new_n897_));
  NOR2_X1   g696(.A1(new_n859_), .A2(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n569_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n523_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g701(.A1(new_n898_), .A2(new_n630_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(KEYINPUT61), .B(G155gat), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1346gat));
  AOI21_X1  g704(.A(G162gat), .B1(new_n898_), .B2(new_n647_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n614_), .A2(new_n575_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n898_), .B2(new_n907_), .ZN(G1347gat));
  NOR2_X1   g707(.A1(new_n661_), .A2(new_n406_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(new_n683_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n910_), .A2(new_n340_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n912_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(KEYINPUT22), .B(G169gat), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n913_), .A2(new_n569_), .A3(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT62), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n856_), .A2(new_n840_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(KEYINPUT121), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n918_), .A2(new_n843_), .A3(new_n865_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n810_), .B1(new_n919_), .B2(new_n629_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT125), .ZN(new_n921_));
  NOR4_X1   g720(.A1(new_n920_), .A2(new_n921_), .A3(new_n570_), .A4(new_n912_), .ZN(new_n922_));
  AOI21_X1  g721(.A(KEYINPUT125), .B1(new_n913_), .B2(new_n569_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n916_), .B1(new_n924_), .B2(G169gat), .ZN(new_n925_));
  NOR4_X1   g724(.A1(new_n922_), .A2(new_n923_), .A3(KEYINPUT62), .A4(new_n223_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n915_), .B1(new_n925_), .B2(new_n926_), .ZN(G1348gat));
  AOI21_X1  g726(.A(G176gat), .B1(new_n913_), .B2(new_n523_), .ZN(new_n928_));
  OR3_X1    g727(.A1(new_n859_), .A2(KEYINPUT126), .A3(new_n340_), .ZN(new_n929_));
  OAI21_X1  g728(.A(KEYINPUT126), .B1(new_n859_), .B2(new_n340_), .ZN(new_n930_));
  AND4_X1   g729(.A1(new_n683_), .A2(new_n929_), .A3(new_n909_), .A4(new_n930_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n522_), .A2(new_n224_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n928_), .B1(new_n931_), .B2(new_n932_), .ZN(G1349gat));
  INV_X1    g732(.A(new_n913_), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n934_), .A2(new_n629_), .A3(new_n358_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n931_), .A2(new_n630_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n935_), .B1(new_n936_), .B2(new_n216_), .ZN(G1350gat));
  OAI21_X1  g736(.A(G190gat), .B1(new_n934_), .B2(new_n614_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n913_), .A2(new_n214_), .A3(new_n647_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1351gat));
  NOR3_X1   g739(.A1(new_n859_), .A2(new_n411_), .A3(new_n683_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(new_n909_), .ZN(new_n942_));
  INV_X1    g741(.A(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(new_n569_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g744(.A1(new_n943_), .A2(new_n523_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g746(.A1(new_n942_), .A2(new_n629_), .ZN(new_n948_));
  NOR3_X1   g747(.A1(new_n948_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n949_));
  XOR2_X1   g748(.A(KEYINPUT63), .B(G211gat), .Z(new_n950_));
  AOI21_X1  g749(.A(new_n949_), .B1(new_n948_), .B2(new_n950_), .ZN(G1354gat));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n952_), .B1(new_n942_), .B2(new_n646_), .ZN(new_n953_));
  INV_X1    g752(.A(G218gat), .ZN(new_n954_));
  NAND4_X1  g753(.A1(new_n941_), .A2(KEYINPUT127), .A3(new_n647_), .A4(new_n909_), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n953_), .A2(new_n954_), .A3(new_n955_), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n943_), .A2(G218gat), .A3(new_n699_), .ZN(new_n957_));
  AND2_X1   g756(.A1(new_n956_), .A2(new_n957_), .ZN(G1355gat));
endmodule


