//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 0 1 0 1 1 0 0 0 0 0 1 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n805_, new_n806_, new_n807_, new_n809_,
    new_n810_, new_n811_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n944_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n965_, new_n966_, new_n967_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n983_, new_n984_, new_n985_, new_n986_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n996_,
    new_n997_, new_n998_, new_n1000_, new_n1001_, new_n1002_, new_n1003_,
    new_n1005_, new_n1007_, new_n1008_, new_n1009_, new_n1011_, new_n1012_,
    new_n1013_;
  INV_X1    g000(.A(KEYINPUT66), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G57gat), .B(G64gat), .ZN(new_n203_));
  AOI21_X1  g002(.A(new_n202_), .B1(new_n203_), .B2(KEYINPUT11), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n203_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT11), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(G71gat), .B(G78gat), .Z(new_n209_));
  NAND3_X1  g008(.A1(new_n203_), .A2(new_n202_), .A3(KEYINPUT11), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n205_), .A2(new_n208_), .A3(new_n209_), .A4(new_n210_), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n209_), .B1(KEYINPUT11), .B2(new_n203_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n210_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n212_), .B1(new_n213_), .B2(new_n204_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G15gat), .B(G22gat), .ZN(new_n216_));
  INV_X1    g015(.A(G1gat), .ZN(new_n217_));
  INV_X1    g016(.A(G8gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT14), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G1gat), .B(G8gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n215_), .B(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G231gat), .A2(G233gat), .ZN(new_n224_));
  XOR2_X1   g023(.A(new_n224_), .B(KEYINPUT71), .Z(new_n225_));
  XNOR2_X1  g024(.A(new_n223_), .B(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(G127gat), .B(G155gat), .Z(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT16), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G183gat), .B(G211gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT17), .ZN(new_n231_));
  OR3_X1    g030(.A1(new_n230_), .A2(KEYINPUT72), .A3(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n231_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n226_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n225_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n223_), .B(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(new_n232_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT73), .ZN(new_n239_));
  AND3_X1   g038(.A1(new_n235_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n239_), .B1(new_n235_), .B2(new_n238_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G232gat), .A2(G233gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT34), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT35), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G29gat), .B(G36gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT69), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G43gat), .B(G50gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT15), .ZN(new_n253_));
  NOR2_X1   g052(.A1(G85gat), .A2(G92gat), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G85gat), .A2(G92gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT65), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  OAI211_X1 g060(.A(KEYINPUT65), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(G99gat), .A2(G106gat), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT7), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT6), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n267_), .B1(G99gat), .B2(G106gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G99gat), .A2(G106gat), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n269_), .A2(KEYINPUT6), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n266_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n258_), .B1(new_n263_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT8), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  OAI211_X1 g073(.A(KEYINPUT8), .B(new_n258_), .C1(new_n263_), .C2(new_n271_), .ZN(new_n275_));
  INV_X1    g074(.A(G92gat), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n276_), .A2(KEYINPUT9), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n277_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n256_), .ZN(new_n279_));
  NOR3_X1   g078(.A1(new_n279_), .A2(new_n254_), .A3(KEYINPUT9), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT64), .B1(new_n278_), .B2(new_n280_), .ZN(new_n281_));
  OAI22_X1  g080(.A1(new_n279_), .A2(new_n254_), .B1(KEYINPUT9), .B2(new_n276_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT64), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n282_), .B(new_n283_), .C1(new_n257_), .C2(KEYINPUT9), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n268_), .A2(new_n270_), .ZN(new_n285_));
  AND2_X1   g084(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n286_));
  NOR2_X1   g085(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n287_));
  NOR3_X1   g086(.A1(new_n286_), .A2(new_n287_), .A3(G106gat), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n285_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n281_), .A2(new_n284_), .A3(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n274_), .A2(new_n275_), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n253_), .A2(new_n291_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n252_), .A2(new_n275_), .A3(new_n290_), .A4(new_n274_), .ZN(new_n293_));
  AOI21_X1  g092(.A(KEYINPUT70), .B1(new_n245_), .B2(new_n246_), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n248_), .B1(new_n292_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G190gat), .B(G218gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G134gat), .B(G162gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n300_), .A2(KEYINPUT36), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n292_), .A2(new_n248_), .A3(new_n295_), .ZN(new_n302_));
  AND3_X1   g101(.A1(new_n297_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n300_), .B(KEYINPUT36), .Z(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n305_), .B1(new_n297_), .B2(new_n302_), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT37), .B1(new_n303_), .B2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n297_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT37), .ZN(new_n309_));
  INV_X1    g108(.A(new_n302_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n310_), .A2(new_n296_), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n308_), .B(new_n309_), .C1(new_n311_), .C2(new_n305_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n242_), .B1(new_n307_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n291_), .A2(new_n215_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT67), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(KEYINPUT12), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G230gat), .A2(G233gat), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n211_), .A2(new_n214_), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n318_), .A2(new_n275_), .A3(new_n290_), .A4(new_n274_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT67), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n320_), .B1(new_n291_), .B2(new_n215_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT12), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n316_), .A2(new_n317_), .A3(new_n319_), .A4(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n319_), .A2(new_n314_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n317_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n324_), .A2(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(G120gat), .B(G148gat), .Z(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G176gat), .B(G204gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n328_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n328_), .A2(new_n333_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT13), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n334_), .A2(KEYINPUT13), .A3(new_n335_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n313_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT74), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G155gat), .A2(G162gat), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT83), .B1(new_n342_), .B2(KEYINPUT1), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT83), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT1), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n344_), .A2(new_n345_), .A3(G155gat), .A4(G162gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n342_), .A2(KEYINPUT1), .ZN(new_n347_));
  OR2_X1    g146(.A1(G155gat), .A2(G162gat), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n343_), .A2(new_n346_), .A3(new_n347_), .A4(new_n348_), .ZN(new_n349_));
  XOR2_X1   g148(.A(G141gat), .B(G148gat), .Z(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT84), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n349_), .A2(KEYINPUT84), .A3(new_n350_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n356_));
  NAND3_X1  g155(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  OR3_X1    g157(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT85), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G141gat), .A2(G148gat), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT2), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n360_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  AND3_X1   g162(.A1(new_n361_), .A2(new_n360_), .A3(new_n362_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n358_), .B(new_n359_), .C1(new_n363_), .C2(new_n364_), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n348_), .A2(new_n342_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(KEYINPUT86), .A3(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(KEYINPUT86), .B1(new_n365_), .B2(new_n366_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n355_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT28), .B1(new_n370_), .B2(KEYINPUT29), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n364_), .A2(new_n363_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n359_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n366_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT86), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  AOI22_X1  g175(.A1(new_n376_), .A2(new_n367_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT28), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT29), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n377_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G22gat), .B(G50gat), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n371_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n381_), .B1(new_n371_), .B2(new_n380_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G228gat), .A2(G233gat), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n377_), .A2(new_n379_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G197gat), .B(G204gat), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT21), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(G218gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(G211gat), .ZN(new_n392_));
  INV_X1    g191(.A(G211gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(G218gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(G197gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(G204gat), .ZN(new_n398_));
  INV_X1    g197(.A(G204gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(G197gat), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n398_), .A2(new_n400_), .A3(KEYINPUT88), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT88), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(new_n397_), .A3(G204gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT21), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n390_), .B(new_n396_), .C1(new_n401_), .C2(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n388_), .A2(new_n389_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n395_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT87), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n386_), .B1(new_n387_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n370_), .A2(KEYINPUT29), .ZN(new_n411_));
  INV_X1    g210(.A(new_n386_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n409_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n411_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G78gat), .B(G106gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT89), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT90), .ZN(new_n419_));
  INV_X1    g218(.A(new_n417_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n410_), .A2(new_n414_), .A3(new_n420_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n385_), .A2(new_n418_), .A3(new_n419_), .A4(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n371_), .A2(new_n380_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n381_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(new_n419_), .A3(new_n382_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n421_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n420_), .B1(new_n410_), .B2(new_n414_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n426_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT90), .B1(new_n383_), .B2(new_n384_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n422_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G226gat), .A2(G233gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT19), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G183gat), .A2(G190gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT23), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT23), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n437_), .A2(G183gat), .A3(G190gat), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT78), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n436_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(G183gat), .A2(G190gat), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n437_), .A2(KEYINPUT78), .A3(G183gat), .A4(G190gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n440_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(G176gat), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT22), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n445_), .B1(new_n446_), .B2(KEYINPUT77), .ZN(new_n447_));
  INV_X1    g246(.A(G169gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  OAI211_X1 g248(.A(G169gat), .B(new_n445_), .C1(new_n446_), .C2(KEYINPUT77), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n444_), .A2(new_n451_), .ZN(new_n452_));
  NOR3_X1   g251(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT25), .B(G183gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(KEYINPUT26), .B(G190gat), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n453_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G169gat), .A2(G176gat), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n457_), .A2(KEYINPUT24), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n448_), .A2(new_n445_), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n458_), .A2(new_n459_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n456_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n452_), .A2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT20), .B1(new_n462_), .B2(new_n408_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n457_), .A2(KEYINPUT24), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT91), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT91), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n457_), .A2(new_n466_), .A3(KEYINPUT24), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n459_), .A3(new_n467_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n456_), .A2(new_n468_), .A3(new_n443_), .A4(new_n440_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT22), .B(G169gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n445_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n436_), .A2(new_n438_), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n471_), .B(new_n457_), .C1(new_n472_), .C2(new_n441_), .ZN(new_n473_));
  AOI22_X1  g272(.A1(new_n469_), .A2(new_n473_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n434_), .B1(new_n463_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n462_), .A2(new_n408_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n395_), .B1(new_n389_), .B2(new_n388_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n398_), .A2(new_n400_), .ZN(new_n478_));
  OAI211_X1 g277(.A(KEYINPUT21), .B(new_n403_), .C1(new_n478_), .C2(new_n402_), .ZN(new_n479_));
  AOI22_X1  g278(.A1(new_n477_), .A2(new_n479_), .B1(new_n395_), .B2(new_n406_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n480_), .A2(new_n473_), .A3(new_n469_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n434_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n476_), .A2(new_n481_), .A3(KEYINPUT20), .A4(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n475_), .A2(KEYINPUT92), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT20), .ZN(new_n485_));
  AOI22_X1  g284(.A1(new_n444_), .A2(new_n451_), .B1(new_n456_), .B2(new_n460_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n485_), .B1(new_n486_), .B2(new_n480_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n469_), .A2(new_n473_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n408_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT92), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n490_), .A2(new_n491_), .A3(new_n434_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G8gat), .B(G36gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G64gat), .B(G92gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n484_), .A2(new_n492_), .A3(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n498_), .B1(new_n484_), .B2(new_n492_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT94), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n499_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  AOI211_X1 g301(.A(KEYINPUT94), .B(new_n498_), .C1(new_n484_), .C2(new_n492_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(G127gat), .B(G134gat), .Z(new_n505_));
  XOR2_X1   g304(.A(G113gat), .B(G120gat), .Z(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G127gat), .B(G134gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G113gat), .B(G120gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n507_), .A2(KEYINPUT81), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT81), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n508_), .A2(new_n509_), .A3(new_n512_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n376_), .A2(new_n367_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n514_), .B1(new_n515_), .B2(new_n355_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT4), .ZN(new_n517_));
  AOI21_X1  g316(.A(KEYINPUT95), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT95), .ZN(new_n519_));
  NOR4_X1   g318(.A1(new_n377_), .A2(new_n519_), .A3(KEYINPUT4), .A4(new_n514_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n511_), .A2(new_n513_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n370_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n507_), .A2(new_n510_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n377_), .A2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(new_n525_), .A3(KEYINPUT4), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G225gat), .A2(G233gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT96), .B1(new_n521_), .B2(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n519_), .B1(new_n523_), .B2(KEYINPUT4), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n516_), .A2(KEYINPUT95), .A3(new_n517_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT96), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n532_), .A2(new_n533_), .A3(new_n527_), .A4(new_n526_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G1gat), .B(G29gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(G85gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT0), .B(G57gat), .ZN(new_n537_));
  XOR2_X1   g336(.A(new_n536_), .B(new_n537_), .Z(new_n538_));
  AOI21_X1  g337(.A(new_n516_), .B1(new_n377_), .B2(new_n524_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n527_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n538_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n529_), .A2(new_n534_), .A3(new_n541_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n526_), .B(new_n540_), .C1(new_n518_), .C2(new_n520_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n539_), .A2(new_n527_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n543_), .A2(KEYINPUT33), .A3(new_n544_), .A4(new_n538_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n543_), .A2(new_n544_), .A3(new_n538_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT33), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n504_), .A2(new_n542_), .A3(new_n545_), .A4(new_n548_), .ZN(new_n549_));
  AOI211_X1 g348(.A(KEYINPUT92), .B(new_n482_), .C1(new_n487_), .C2(new_n489_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n491_), .B1(new_n490_), .B2(new_n434_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n550_), .B1(new_n551_), .B2(new_n483_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n497_), .A2(KEYINPUT32), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(KEYINPUT97), .B1(new_n552_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n484_), .A2(new_n492_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT97), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n556_), .A2(new_n557_), .A3(new_n553_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n555_), .A2(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT20), .B1(new_n488_), .B2(new_n408_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n486_), .A2(new_n480_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n434_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT98), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT98), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n564_), .B(new_n434_), .C1(new_n560_), .C2(new_n561_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n487_), .A2(new_n489_), .A3(new_n482_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n563_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(new_n554_), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n543_), .A2(new_n544_), .A3(new_n538_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n538_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n559_), .B(new_n568_), .C1(new_n569_), .C2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n549_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT27), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n573_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(KEYINPUT99), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT99), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n576_), .B(new_n573_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n575_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n567_), .A2(new_n498_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n556_), .A2(new_n497_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n579_), .A2(KEYINPUT27), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n543_), .A2(new_n544_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n538_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n581_), .A2(new_n584_), .A3(new_n546_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n432_), .A2(new_n585_), .ZN(new_n586_));
  AOI22_X1  g385(.A1(new_n432_), .A2(new_n572_), .B1(new_n578_), .B2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G71gat), .B(G99gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(KEYINPUT79), .B(G43gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n462_), .B(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT82), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n522_), .B(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT31), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n595_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(new_n597_), .A3(KEYINPUT80), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G227gat), .A2(G233gat), .ZN(new_n599_));
  INV_X1    g398(.A(G15gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT30), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n598_), .A2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n598_), .A2(new_n602_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n592_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n598_), .A2(new_n602_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n598_), .A2(new_n602_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n606_), .A2(new_n591_), .A3(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n605_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(KEYINPUT100), .B1(new_n587_), .B2(new_n610_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n578_), .A2(new_n581_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n569_), .A2(new_n570_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n609_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n612_), .A2(new_n432_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT100), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n430_), .B(new_n426_), .C1(new_n427_), .C2(new_n428_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n613_), .A2(new_n422_), .A3(new_n618_), .A4(new_n581_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n619_), .B1(new_n575_), .B2(new_n577_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n618_), .A2(new_n422_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n621_), .B1(new_n549_), .B2(new_n571_), .ZN(new_n622_));
  OAI211_X1 g421(.A(new_n617_), .B(new_n609_), .C1(new_n620_), .C2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n611_), .A2(new_n616_), .A3(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G229gat), .A2(G233gat), .ZN(new_n625_));
  INV_X1    g424(.A(new_n222_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n252_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n252_), .A2(new_n626_), .ZN(new_n629_));
  OAI21_X1  g428(.A(KEYINPUT75), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n252_), .A2(new_n626_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT75), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n631_), .A2(new_n632_), .A3(new_n627_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n625_), .B1(new_n630_), .B2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n627_), .A2(new_n625_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n253_), .B2(new_n222_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  XOR2_X1   g436(.A(G113gat), .B(G141gat), .Z(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT76), .ZN(new_n639_));
  XNOR2_X1  g438(.A(G169gat), .B(G197gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n637_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n641_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n643_), .B1(new_n634_), .B2(new_n636_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n341_), .A2(new_n624_), .A3(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n645_), .ZN(new_n649_));
  AND4_X1   g448(.A1(new_n432_), .A2(new_n615_), .A3(new_n578_), .A4(new_n581_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n572_), .A2(new_n432_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n578_), .A2(new_n586_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n610_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n650_), .B1(new_n653_), .B2(new_n617_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n649_), .B1(new_n654_), .B2(new_n611_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n655_), .A2(KEYINPUT101), .A3(new_n341_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n648_), .A2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(new_n217_), .A3(new_n614_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT38), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(KEYINPUT102), .B1(new_n303_), .B2(new_n306_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT102), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n308_), .B(new_n662_), .C1(new_n311_), .C2(new_n305_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n624_), .A2(KEYINPUT103), .A3(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT103), .B1(new_n624_), .B2(new_n665_), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n338_), .A2(new_n339_), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n669_), .A2(new_n649_), .A3(new_n242_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n668_), .A2(new_n614_), .A3(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(G1gat), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n658_), .A2(new_n659_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n660_), .A2(new_n672_), .A3(new_n673_), .ZN(G1324gat));
  NOR2_X1   g473(.A1(new_n612_), .A2(G8gat), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n648_), .A2(new_n656_), .A3(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n676_), .B(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n578_), .A2(new_n581_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n679_), .B(new_n670_), .C1(new_n666_), .C2(new_n667_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n680_), .A2(KEYINPUT39), .A3(G8gat), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(G8gat), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT39), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n678_), .A2(new_n681_), .A3(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT40), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n678_), .A2(KEYINPUT40), .A3(new_n684_), .A4(new_n681_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1325gat));
  NAND3_X1  g488(.A1(new_n657_), .A2(new_n600_), .A3(new_n610_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n668_), .A2(new_n610_), .A3(new_n670_), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n691_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(KEYINPUT41), .B1(new_n691_), .B2(G15gat), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n690_), .B1(new_n692_), .B2(new_n693_), .ZN(G1326gat));
  INV_X1    g493(.A(G22gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n657_), .A2(new_n695_), .A3(new_n621_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n668_), .A2(new_n621_), .A3(new_n670_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(G22gat), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n698_), .A2(KEYINPUT42), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n698_), .A2(KEYINPUT42), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n696_), .B1(new_n699_), .B2(new_n700_), .ZN(G1327gat));
  INV_X1    g500(.A(new_n242_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n665_), .A2(new_n702_), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n703_), .A2(KEYINPUT106), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(KEYINPUT106), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n669_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n706_), .A2(new_n624_), .A3(new_n645_), .A4(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(KEYINPUT107), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n655_), .A2(new_n710_), .A3(new_n707_), .A4(new_n706_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n709_), .A2(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(G29gat), .B1(new_n712_), .B2(new_n614_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n669_), .A2(new_n649_), .A3(new_n702_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n307_), .A2(new_n312_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n623_), .A2(new_n616_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n651_), .A2(new_n652_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n617_), .B1(new_n720_), .B2(new_n609_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n718_), .B1(new_n719_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT43), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT43), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n624_), .A2(new_n724_), .A3(new_n718_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n716_), .B1(new_n723_), .B2(new_n725_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n714_), .B1(new_n726_), .B2(KEYINPUT44), .ZN(new_n727_));
  AOI211_X1 g526(.A(KEYINPUT43), .B(new_n717_), .C1(new_n654_), .C2(new_n611_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n724_), .B1(new_n624_), .B2(new_n718_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n715_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(KEYINPUT105), .A3(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n727_), .A2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n723_), .A2(new_n725_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(KEYINPUT44), .A3(new_n715_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n614_), .A2(G29gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n713_), .B1(new_n737_), .B2(new_n738_), .ZN(G1328gat));
  INV_X1    g538(.A(KEYINPUT46), .ZN(new_n740_));
  INV_X1    g539(.A(G36gat), .ZN(new_n741_));
  AOI211_X1 g540(.A(new_n731_), .B(new_n716_), .C1(new_n723_), .C2(new_n725_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n742_), .A2(new_n612_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n741_), .B1(new_n733_), .B2(new_n743_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n612_), .A2(G36gat), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n709_), .A2(new_n711_), .A3(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT45), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n746_), .B(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n740_), .B1(new_n744_), .B2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n746_), .B(KEYINPUT45), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n735_), .A2(new_n679_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n727_), .B2(new_n732_), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n750_), .B(KEYINPUT46), .C1(new_n752_), .C2(new_n741_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n749_), .A2(new_n753_), .ZN(G1329gat));
  NAND2_X1  g553(.A1(new_n610_), .A2(G43gat), .ZN(new_n755_));
  AOI211_X1 g554(.A(new_n755_), .B(new_n742_), .C1(new_n727_), .C2(new_n732_), .ZN(new_n756_));
  AOI21_X1  g555(.A(G43gat), .B1(new_n712_), .B2(new_n610_), .ZN(new_n757_));
  OAI21_X1  g556(.A(KEYINPUT47), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n757_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT47), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n759_), .B(new_n760_), .C1(new_n736_), .C2(new_n755_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n758_), .A2(new_n761_), .ZN(G1330gat));
  AOI21_X1  g561(.A(G50gat), .B1(new_n712_), .B2(new_n621_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n621_), .A2(G50gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n737_), .B2(new_n764_), .ZN(G1331gat));
  NAND2_X1  g564(.A1(new_n669_), .A2(new_n649_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n766_), .A2(new_n242_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n668_), .A2(new_n614_), .A3(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(G57gat), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n766_), .B1(new_n654_), .B2(new_n611_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n770_), .A2(new_n313_), .ZN(new_n771_));
  INV_X1    g570(.A(G57gat), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n772_), .A3(new_n614_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n769_), .A2(new_n773_), .ZN(G1332gat));
  INV_X1    g573(.A(G64gat), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n771_), .A2(new_n775_), .A3(new_n679_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n668_), .A2(new_n679_), .A3(new_n767_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(G64gat), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n778_), .A2(KEYINPUT48), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n778_), .A2(KEYINPUT48), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n776_), .B1(new_n779_), .B2(new_n780_), .ZN(G1333gat));
  INV_X1    g580(.A(G71gat), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n771_), .A2(new_n782_), .A3(new_n610_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n668_), .A2(new_n610_), .A3(new_n767_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(G71gat), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n785_), .A2(KEYINPUT49), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n785_), .A2(KEYINPUT49), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n783_), .B1(new_n786_), .B2(new_n787_), .ZN(G1334gat));
  NOR2_X1   g587(.A1(new_n432_), .A2(G78gat), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT108), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n771_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n668_), .A2(new_n621_), .A3(new_n767_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(G78gat), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n793_), .A2(KEYINPUT50), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n793_), .A2(KEYINPUT50), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n791_), .B1(new_n794_), .B2(new_n795_), .ZN(G1335gat));
  AND2_X1   g595(.A1(new_n770_), .A2(new_n706_), .ZN(new_n797_));
  AOI21_X1  g596(.A(G85gat), .B1(new_n797_), .B2(new_n614_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT109), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n766_), .A2(new_n702_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n723_), .B2(new_n725_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n802_), .A2(G85gat), .A3(new_n614_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n799_), .A2(new_n803_), .ZN(G1336gat));
  AOI21_X1  g603(.A(G92gat), .B1(new_n797_), .B2(new_n679_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(KEYINPUT110), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n612_), .A2(new_n276_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n802_), .B2(new_n807_), .ZN(G1337gat));
  NAND2_X1  g607(.A1(new_n802_), .A2(new_n610_), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n609_), .A2(new_n287_), .A3(new_n286_), .ZN(new_n810_));
  AOI22_X1  g609(.A1(new_n809_), .A2(G99gat), .B1(new_n797_), .B2(new_n810_), .ZN(new_n811_));
  XOR2_X1   g610(.A(new_n811_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g611(.A(G106gat), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n621_), .B(new_n800_), .C1(new_n728_), .C2(new_n729_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n813_), .B1(new_n815_), .B2(KEYINPUT112), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT112), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n814_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT52), .B1(new_n816_), .B2(new_n818_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n734_), .A2(KEYINPUT112), .A3(new_n621_), .A4(new_n800_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n818_), .A2(KEYINPUT52), .A3(new_n820_), .A4(G106gat), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n770_), .A2(new_n813_), .A3(new_n706_), .A4(new_n621_), .ZN(new_n822_));
  XOR2_X1   g621(.A(new_n822_), .B(KEYINPUT111), .Z(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(KEYINPUT53), .B1(new_n819_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n826_));
  INV_X1    g625(.A(new_n818_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n820_), .A2(G106gat), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n826_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n829_), .A2(new_n830_), .A3(new_n821_), .A4(new_n823_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n825_), .A2(new_n831_), .ZN(G1339gat));
  NOR4_X1   g631(.A1(new_n679_), .A2(new_n609_), .A3(new_n621_), .A4(new_n613_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n645_), .A2(new_n334_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n319_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n835_));
  AOI211_X1 g634(.A(new_n320_), .B(KEYINPUT12), .C1(new_n291_), .C2(new_n215_), .ZN(new_n836_));
  NOR3_X1   g635(.A1(new_n835_), .A2(new_n326_), .A3(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT55), .B1(new_n837_), .B2(KEYINPUT114), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT114), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n324_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT115), .B1(new_n835_), .B2(new_n836_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n316_), .A2(new_n843_), .A3(new_n319_), .A4(new_n323_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n842_), .A2(new_n844_), .A3(new_n326_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n838_), .A2(new_n841_), .A3(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n333_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT56), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n846_), .A2(KEYINPUT56), .A3(new_n333_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n834_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n630_), .A2(new_n633_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n625_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n253_), .A2(new_n222_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n628_), .A2(new_n625_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n641_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  AOI22_X1  g655(.A1(new_n637_), .A2(new_n641_), .B1(new_n853_), .B2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n336_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  OAI211_X1 g658(.A(KEYINPUT57), .B(new_n665_), .C1(new_n851_), .C2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT116), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n645_), .A2(new_n334_), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n846_), .A2(KEYINPUT56), .A3(new_n333_), .ZN(new_n864_));
  AOI21_X1  g663(.A(KEYINPUT56), .B1(new_n846_), .B2(new_n333_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n863_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n664_), .B1(new_n866_), .B2(new_n858_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(KEYINPUT116), .A3(KEYINPUT57), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n862_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n866_), .A2(new_n858_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n665_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n857_), .A2(new_n334_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n874_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT58), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n717_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n874_), .B(KEYINPUT58), .C1(new_n864_), .C2(new_n865_), .ZN(new_n878_));
  AOI22_X1  g677(.A1(new_n871_), .A2(new_n872_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n702_), .B1(new_n869_), .B2(new_n879_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n718_), .A2(new_n669_), .A3(new_n242_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n881_), .A2(KEYINPUT113), .A3(new_n882_), .A4(new_n649_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT113), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n707_), .A2(new_n649_), .A3(new_n313_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(KEYINPUT54), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(KEYINPUT54), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n883_), .A2(new_n886_), .A3(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n833_), .B1(new_n880_), .B2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT118), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n875_), .A2(new_n876_), .ZN(new_n894_));
  AND3_X1   g693(.A1(new_n894_), .A2(new_n718_), .A3(new_n878_), .ZN(new_n895_));
  AOI21_X1  g694(.A(KEYINPUT57), .B1(new_n870_), .B2(new_n665_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n893_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n894_), .A2(new_n718_), .A3(new_n878_), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n898_), .B(KEYINPUT118), .C1(KEYINPUT57), .C2(new_n867_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n897_), .A2(new_n869_), .A3(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n889_), .B1(new_n900_), .B2(new_n242_), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n833_), .A2(KEYINPUT117), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n833_), .A2(KEYINPUT117), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n902_), .A2(new_n892_), .A3(new_n903_), .ZN(new_n904_));
  OAI22_X1  g703(.A1(new_n891_), .A2(new_n892_), .B1(new_n901_), .B2(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(G113gat), .B1(new_n905_), .B2(new_n649_), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n649_), .A2(G113gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n890_), .B2(new_n907_), .ZN(G1340gat));
  XNOR2_X1  g707(.A(KEYINPUT119), .B(G120gat), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n909_), .B1(new_n905_), .B2(new_n707_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT60), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n909_), .B1(new_n669_), .B2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(KEYINPUT120), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT120), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n914_), .B1(new_n909_), .B2(new_n911_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n913_), .B1(new_n912_), .B2(new_n915_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n910_), .B1(new_n890_), .B2(new_n916_), .ZN(G1341gat));
  OAI21_X1  g716(.A(G127gat), .B1(new_n905_), .B2(new_n242_), .ZN(new_n918_));
  OR2_X1    g717(.A1(new_n242_), .A2(G127gat), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n890_), .B2(new_n919_), .ZN(G1342gat));
  INV_X1    g719(.A(G134gat), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n900_), .A2(new_n242_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(new_n888_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n904_), .ZN(new_n924_));
  AOI22_X1  g723(.A1(new_n923_), .A2(new_n924_), .B1(KEYINPUT59), .B2(new_n890_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n921_), .B1(new_n925_), .B2(new_n718_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n891_), .A2(new_n921_), .A3(new_n664_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(KEYINPUT121), .B1(new_n926_), .B2(new_n928_), .ZN(new_n929_));
  OAI21_X1  g728(.A(G134gat), .B1(new_n905_), .B2(new_n717_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT121), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n930_), .A2(new_n931_), .A3(new_n927_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n929_), .A2(new_n932_), .ZN(G1343gat));
  NOR2_X1   g732(.A1(new_n610_), .A2(new_n432_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  NOR3_X1   g734(.A1(new_n935_), .A2(new_n679_), .A3(new_n613_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n936_), .B1(new_n880_), .B2(new_n889_), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT122), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n937_), .A2(new_n938_), .ZN(new_n939_));
  OAI211_X1 g738(.A(KEYINPUT122), .B(new_n936_), .C1(new_n880_), .C2(new_n889_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(new_n645_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g742(.A1(new_n941_), .A2(new_n669_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g744(.A(KEYINPUT61), .B(G155gat), .ZN(new_n946_));
  INV_X1    g745(.A(new_n946_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT123), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n948_), .B1(new_n941_), .B2(new_n702_), .ZN(new_n949_));
  AOI211_X1 g748(.A(KEYINPUT123), .B(new_n242_), .C1(new_n939_), .C2(new_n940_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n947_), .B1(new_n949_), .B2(new_n950_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n873_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n718_), .B1(new_n952_), .B2(KEYINPUT58), .ZN(new_n953_));
  INV_X1    g752(.A(new_n878_), .ZN(new_n954_));
  OAI22_X1  g753(.A1(new_n953_), .A2(new_n954_), .B1(new_n867_), .B2(KEYINPUT57), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n955_), .B1(new_n862_), .B2(new_n868_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n888_), .B1(new_n956_), .B2(new_n702_), .ZN(new_n957_));
  AOI21_X1  g756(.A(KEYINPUT122), .B1(new_n957_), .B2(new_n936_), .ZN(new_n958_));
  INV_X1    g757(.A(new_n940_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n702_), .B1(new_n958_), .B2(new_n959_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n960_), .A2(KEYINPUT123), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n941_), .A2(new_n948_), .A3(new_n702_), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n961_), .A2(new_n962_), .A3(new_n946_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n951_), .A2(new_n963_), .ZN(G1346gat));
  INV_X1    g763(.A(new_n941_), .ZN(new_n965_));
  OR3_X1    g764(.A1(new_n965_), .A2(G162gat), .A3(new_n665_), .ZN(new_n966_));
  OAI21_X1  g765(.A(G162gat), .B1(new_n965_), .B2(new_n717_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n966_), .A2(new_n967_), .ZN(G1347gat));
  AND2_X1   g767(.A1(new_n679_), .A2(new_n615_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n969_), .A2(new_n432_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(new_n901_), .A2(new_n970_), .ZN(new_n971_));
  NAND3_X1  g770(.A1(new_n971_), .A2(new_n470_), .A3(new_n645_), .ZN(new_n972_));
  AOI21_X1  g771(.A(KEYINPUT124), .B1(new_n969_), .B2(new_n645_), .ZN(new_n973_));
  AND3_X1   g772(.A1(new_n969_), .A2(KEYINPUT124), .A3(new_n645_), .ZN(new_n974_));
  OAI211_X1 g773(.A(new_n923_), .B(new_n432_), .C1(new_n973_), .C2(new_n974_), .ZN(new_n975_));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n976_));
  NOR2_X1   g775(.A1(new_n976_), .A2(KEYINPUT62), .ZN(new_n977_));
  AOI21_X1  g776(.A(new_n448_), .B1(new_n976_), .B2(KEYINPUT62), .ZN(new_n978_));
  NAND3_X1  g777(.A1(new_n975_), .A2(new_n977_), .A3(new_n978_), .ZN(new_n979_));
  INV_X1    g778(.A(new_n979_), .ZN(new_n980_));
  AOI21_X1  g779(.A(new_n977_), .B1(new_n975_), .B2(new_n978_), .ZN(new_n981_));
  OAI21_X1  g780(.A(new_n972_), .B1(new_n980_), .B2(new_n981_), .ZN(G1348gat));
  AOI21_X1  g781(.A(G176gat), .B1(new_n971_), .B2(new_n669_), .ZN(new_n983_));
  NOR2_X1   g782(.A1(new_n880_), .A2(new_n889_), .ZN(new_n984_));
  NOR2_X1   g783(.A1(new_n984_), .A2(new_n621_), .ZN(new_n985_));
  AND3_X1   g784(.A1(new_n969_), .A2(G176gat), .A3(new_n669_), .ZN(new_n986_));
  AOI21_X1  g785(.A(new_n983_), .B1(new_n985_), .B2(new_n986_), .ZN(G1349gat));
  INV_X1    g786(.A(new_n454_), .ZN(new_n988_));
  NAND3_X1  g787(.A1(new_n971_), .A2(new_n988_), .A3(new_n702_), .ZN(new_n989_));
  INV_X1    g788(.A(KEYINPUT126), .ZN(new_n990_));
  AND2_X1   g789(.A1(new_n989_), .A2(new_n990_), .ZN(new_n991_));
  NOR2_X1   g790(.A1(new_n989_), .A2(new_n990_), .ZN(new_n992_));
  AND2_X1   g791(.A1(new_n969_), .A2(new_n702_), .ZN(new_n993_));
  AOI21_X1  g792(.A(G183gat), .B1(new_n985_), .B2(new_n993_), .ZN(new_n994_));
  NOR3_X1   g793(.A1(new_n991_), .A2(new_n992_), .A3(new_n994_), .ZN(G1350gat));
  NAND3_X1  g794(.A1(new_n971_), .A2(new_n455_), .A3(new_n664_), .ZN(new_n996_));
  NOR3_X1   g795(.A1(new_n901_), .A2(new_n717_), .A3(new_n970_), .ZN(new_n997_));
  INV_X1    g796(.A(G190gat), .ZN(new_n998_));
  OAI21_X1  g797(.A(new_n996_), .B1(new_n997_), .B2(new_n998_), .ZN(G1351gat));
  NOR3_X1   g798(.A1(new_n935_), .A2(new_n612_), .A3(new_n614_), .ZN(new_n1000_));
  NAND2_X1  g799(.A1(new_n957_), .A2(new_n1000_), .ZN(new_n1001_));
  INV_X1    g800(.A(new_n1001_), .ZN(new_n1002_));
  NAND2_X1  g801(.A1(new_n1002_), .A2(new_n645_), .ZN(new_n1003_));
  XNOR2_X1  g802(.A(new_n1003_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g803(.A1(new_n1002_), .A2(new_n669_), .ZN(new_n1005_));
  XNOR2_X1  g804(.A(new_n1005_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g805(.A(KEYINPUT63), .ZN(new_n1007_));
  OAI211_X1 g806(.A(new_n1002_), .B(new_n702_), .C1(new_n1007_), .C2(new_n393_), .ZN(new_n1008_));
  NAND2_X1  g807(.A1(new_n1007_), .A2(new_n393_), .ZN(new_n1009_));
  XNOR2_X1  g808(.A(new_n1008_), .B(new_n1009_), .ZN(G1354gat));
  OAI21_X1  g809(.A(G218gat), .B1(new_n1001_), .B2(new_n717_), .ZN(new_n1011_));
  NAND2_X1  g810(.A1(new_n664_), .A2(new_n391_), .ZN(new_n1012_));
  OAI21_X1  g811(.A(new_n1011_), .B1(new_n1001_), .B2(new_n1012_), .ZN(new_n1013_));
  XNOR2_X1  g812(.A(new_n1013_), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


