//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1 0 1 0 1 0 0 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 0 1 0 0 0 0 0 1 0 1 1 1 1 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n800_, new_n801_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n812_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n844_,
    new_n845_, new_n846_, new_n848_, new_n849_, new_n851_, new_n852_,
    new_n853_, new_n855_, new_n856_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT4), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G127gat), .B(G134gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G113gat), .B(G120gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT84), .ZN(new_n208_));
  AND2_X1   g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(G141gat), .ZN(new_n212_));
  INV_X1    g011(.A(G148gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT88), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n214_), .B(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  XOR2_X1   g017(.A(new_n218_), .B(KEYINPUT2), .Z(new_n219_));
  OAI21_X1  g018(.A(new_n211_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT1), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n211_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n209_), .A2(KEYINPUT1), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n222_), .A2(new_n218_), .A3(new_n214_), .A4(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n220_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n208_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n207_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n204_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n208_), .A2(new_n226_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n230_), .A2(KEYINPUT4), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n203_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n227_), .A2(new_n202_), .A3(new_n228_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G1gat), .B(G29gat), .Z(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(G85gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT0), .B(G57gat), .ZN(new_n236_));
  XOR2_X1   g035(.A(new_n235_), .B(new_n236_), .Z(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n232_), .A2(new_n233_), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT33), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT98), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT98), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n239_), .A2(new_n243_), .A3(new_n240_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G197gat), .B(G204gat), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT21), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G211gat), .B(G218gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n246_), .A2(new_n247_), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n251_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT91), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT26), .B(G190gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT25), .B(G183gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  OR2_X1    g058(.A1(G169gat), .A2(G176gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G169gat), .A2(G176gat), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(KEYINPUT24), .A3(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n259_), .A2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT80), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n260_), .A2(KEYINPUT24), .ZN(new_n265_));
  INV_X1    g064(.A(G183gat), .ZN(new_n266_));
  INV_X1    g065(.A(G190gat), .ZN(new_n267_));
  OR3_X1    g066(.A1(new_n266_), .A2(new_n267_), .A3(KEYINPUT23), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT23), .B1(new_n266_), .B2(new_n267_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n265_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT81), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n264_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n261_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT22), .B(G169gat), .ZN(new_n274_));
  INV_X1    g073(.A(G176gat), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n273_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT82), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n268_), .A2(new_n277_), .A3(new_n269_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n278_), .B1(new_n277_), .B2(new_n268_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(G183gat), .A2(G190gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n276_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n272_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n256_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT97), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n256_), .A2(KEYINPUT97), .A3(new_n282_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n258_), .B(KEYINPUT95), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n287_), .A2(new_n257_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n262_), .ZN(new_n289_));
  NOR4_X1   g088(.A1(new_n288_), .A2(new_n279_), .A3(new_n289_), .A4(new_n265_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n276_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n280_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n290_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n254_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n285_), .A2(new_n286_), .A3(KEYINPUT20), .A4(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G226gat), .A2(G233gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT19), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT96), .B1(new_n294_), .B2(new_n295_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT96), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n303_), .B(new_n254_), .C1(new_n290_), .C2(new_n293_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n256_), .A2(new_n282_), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n305_), .A2(KEYINPUT20), .A3(new_n299_), .A4(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n301_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G8gat), .B(G36gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(G92gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT18), .B(G64gat), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n310_), .B(new_n311_), .Z(new_n312_));
  NAND2_X1  g111(.A1(new_n308_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n312_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n301_), .A2(new_n307_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n239_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT33), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n245_), .A2(new_n313_), .A3(new_n315_), .A4(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n202_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n227_), .A2(new_n203_), .A3(new_n228_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(new_n237_), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT99), .B1(new_n318_), .B2(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n238_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n324_), .A2(KEYINPUT100), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(KEYINPUT100), .ZN(new_n326_));
  NOR3_X1   g125(.A1(new_n325_), .A2(new_n326_), .A3(new_n316_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT32), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n308_), .B1(new_n329_), .B2(new_n314_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n297_), .A2(new_n299_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n305_), .A2(KEYINPUT20), .A3(new_n300_), .A4(new_n306_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n333_), .A2(KEYINPUT32), .A3(new_n312_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n328_), .A2(new_n330_), .A3(new_n334_), .ZN(new_n335_));
  AND3_X1   g134(.A1(new_n313_), .A2(new_n315_), .A3(new_n317_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT99), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n336_), .A2(new_n337_), .A3(new_n321_), .A4(new_n245_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n323_), .A2(new_n335_), .A3(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n225_), .A2(KEYINPUT29), .ZN(new_n340_));
  INV_X1    g139(.A(G50gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  XOR2_X1   g141(.A(KEYINPUT89), .B(G22gat), .Z(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n342_), .B(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G228gat), .A2(G233gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n225_), .A2(KEYINPUT29), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n348_), .B1(new_n349_), .B2(new_n254_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT92), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n351_), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n349_), .A2(new_n348_), .ZN(new_n354_));
  AOI22_X1  g153(.A1(new_n352_), .A2(new_n353_), .B1(new_n256_), .B2(new_n354_), .ZN(new_n355_));
  XOR2_X1   g154(.A(G78gat), .B(G106gat), .Z(new_n356_));
  AND2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n355_), .A2(new_n356_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n347_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT93), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n358_), .A2(KEYINPUT94), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT94), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n363_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n355_), .A2(new_n356_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n362_), .A2(new_n346_), .A3(new_n364_), .A4(new_n365_), .ZN(new_n366_));
  OAI211_X1 g165(.A(KEYINPUT93), .B(new_n347_), .C1(new_n357_), .C2(new_n358_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n361_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n339_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT27), .ZN(new_n371_));
  INV_X1    g170(.A(new_n315_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n314_), .B1(new_n301_), .B2(new_n307_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n371_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n333_), .A2(new_n314_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n313_), .A2(new_n375_), .A3(KEYINPUT27), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n368_), .A2(new_n374_), .A3(new_n376_), .A4(new_n327_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT101), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n370_), .A2(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n282_), .B(KEYINPUT30), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT83), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G15gat), .B(G43gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(G99gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G227gat), .A2(G233gat), .ZN(new_n385_));
  XOR2_X1   g184(.A(new_n385_), .B(G71gat), .Z(new_n386_));
  XNOR2_X1  g185(.A(new_n384_), .B(new_n386_), .ZN(new_n387_));
  OR2_X1    g186(.A1(new_n382_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n208_), .B(KEYINPUT31), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT30), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n282_), .B(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT83), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n382_), .A2(new_n392_), .A3(new_n387_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n388_), .A2(new_n389_), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT85), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n394_), .A2(new_n395_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT86), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n388_), .A2(new_n393_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n389_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n398_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  AOI211_X1 g200(.A(KEYINPUT86), .B(new_n389_), .C1(new_n388_), .C2(new_n393_), .ZN(new_n402_));
  OAI22_X1  g201(.A1(new_n396_), .A2(new_n397_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT87), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT87), .ZN(new_n405_));
  OAI221_X1 g204(.A(new_n405_), .B1(new_n401_), .B2(new_n402_), .C1(new_n396_), .C2(new_n397_), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n379_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n404_), .A2(new_n406_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n374_), .A2(new_n376_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n410_), .A2(new_n328_), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n409_), .A2(new_n369_), .A3(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n408_), .A2(new_n413_), .ZN(new_n414_));
  AND3_X1   g213(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n415_));
  AOI21_X1  g214(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT65), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G99gat), .A2(G106gat), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT6), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT65), .ZN(new_n421_));
  NAND3_X1  g220(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n420_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n417_), .A2(new_n423_), .ZN(new_n424_));
  XOR2_X1   g223(.A(KEYINPUT10), .B(G99gat), .Z(new_n425_));
  INV_X1    g224(.A(G106gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  XOR2_X1   g226(.A(G85gat), .B(G92gat), .Z(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT9), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT9), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(G85gat), .A3(G92gat), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n424_), .A2(new_n427_), .A3(new_n429_), .A4(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT8), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n428_), .A2(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(G99gat), .A2(G106gat), .ZN(new_n435_));
  AND2_X1   g234(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n436_));
  NOR2_X1   g235(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n435_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  OAI22_X1  g237(.A1(KEYINPUT66), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n434_), .B1(new_n440_), .B2(new_n424_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n415_), .A2(new_n416_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n442_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n433_), .B1(new_n443_), .B2(new_n428_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n432_), .B1(new_n441_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT67), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  OAI211_X1 g246(.A(KEYINPUT67), .B(new_n432_), .C1(new_n441_), .C2(new_n444_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G57gat), .B(G64gat), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n450_), .A2(KEYINPUT11), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(KEYINPUT11), .ZN(new_n452_));
  XOR2_X1   g251(.A(G71gat), .B(G78gat), .Z(new_n453_));
  NAND3_X1  g252(.A1(new_n451_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n452_), .A2(new_n453_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n449_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT68), .ZN(new_n458_));
  INV_X1    g257(.A(new_n456_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n447_), .A2(new_n448_), .A3(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n457_), .A2(new_n458_), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G230gat), .A2(G233gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT64), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n447_), .A2(new_n448_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n465_), .A2(KEYINPUT68), .A3(new_n459_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n461_), .A2(new_n464_), .A3(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT69), .B(KEYINPUT12), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n460_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n445_), .A2(KEYINPUT12), .A3(new_n459_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n469_), .A2(new_n457_), .A3(new_n463_), .A4(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n467_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G120gat), .B(G148gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(G204gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT5), .B(G176gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n474_), .B(new_n475_), .Z(new_n476_));
  NAND2_X1  g275(.A1(new_n472_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n476_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n467_), .A2(new_n471_), .A3(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT13), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n477_), .A2(KEYINPUT13), .A3(new_n479_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G229gat), .A2(G233gat), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(G1gat), .ZN(new_n487_));
  INV_X1    g286(.A(G8gat), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT14), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT74), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G15gat), .B(G22gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G1gat), .B(G8gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT75), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n492_), .A2(new_n494_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G29gat), .B(G36gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(new_n341_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT70), .B(G43gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n498_), .B(G50gat), .ZN(new_n502_));
  INV_X1    g301(.A(new_n500_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n501_), .A2(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n497_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n505_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n507_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n486_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT15), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n505_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n501_), .A2(new_n504_), .A3(KEYINPUT15), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n511_), .A2(new_n495_), .A3(new_n496_), .A4(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n497_), .A2(new_n505_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(new_n514_), .A3(new_n485_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n509_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT79), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G113gat), .B(G141gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G169gat), .B(G197gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n517_), .A2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n516_), .A2(KEYINPUT79), .A3(new_n520_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G127gat), .B(G155gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(G211gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT16), .B(G183gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  XOR2_X1   g328(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n531_), .B(KEYINPUT77), .Z(new_n532_));
  NAND2_X1  g331(.A1(G231gat), .A2(G233gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n456_), .B(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(new_n497_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n532_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT78), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n529_), .B(KEYINPUT17), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n535_), .A2(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NOR3_X1   g340(.A1(new_n484_), .A2(new_n525_), .A3(new_n541_), .ZN(new_n542_));
  OR2_X1    g341(.A1(KEYINPUT73), .A2(KEYINPUT37), .ZN(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT71), .B1(new_n465_), .B2(new_n507_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT71), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n449_), .A2(new_n547_), .A3(new_n505_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n511_), .A2(new_n512_), .A3(new_n445_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n546_), .A2(new_n548_), .A3(new_n549_), .A4(KEYINPUT72), .ZN(new_n550_));
  INV_X1    g349(.A(G232gat), .ZN(new_n551_));
  INV_X1    g350(.A(G233gat), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n550_), .A2(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n550_), .A2(new_n554_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n545_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n550_), .A2(new_n554_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n550_), .A2(new_n554_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n558_), .A2(new_n544_), .A3(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G190gat), .B(G218gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G134gat), .B(G162gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n561_), .B(new_n562_), .Z(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT36), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n546_), .A2(new_n548_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(new_n549_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT35), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n557_), .A2(new_n560_), .A3(new_n565_), .A4(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n564_), .A2(KEYINPUT36), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n570_), .A2(new_n571_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n543_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n557_), .A2(new_n560_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n571_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n575_), .A2(new_n576_), .A3(new_n565_), .A4(new_n569_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n570_), .A2(new_n571_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(KEYINPUT73), .B(KEYINPUT37), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n577_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n574_), .A2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n414_), .A2(new_n542_), .A3(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n582_), .B(KEYINPUT102), .Z(new_n583_));
  NAND3_X1  g382(.A1(new_n583_), .A2(new_n487_), .A3(new_n328_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT38), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n542_), .B(KEYINPUT103), .Z(new_n586_));
  NAND2_X1  g385(.A1(new_n577_), .A2(new_n578_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n414_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT104), .ZN(new_n589_));
  OAI21_X1  g388(.A(G1gat), .B1(new_n589_), .B2(new_n327_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n585_), .A2(new_n590_), .ZN(G1324gat));
  INV_X1    g390(.A(new_n410_), .ZN(new_n592_));
  OAI21_X1  g391(.A(G8gat), .B1(new_n588_), .B2(new_n592_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n593_), .A2(KEYINPUT105), .ZN(new_n594_));
  OAI21_X1  g393(.A(KEYINPUT39), .B1(new_n593_), .B2(KEYINPUT105), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n583_), .A2(new_n488_), .A3(new_n410_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n594_), .A2(new_n595_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n596_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT40), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n596_), .A2(KEYINPUT40), .A3(new_n597_), .A4(new_n598_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(G1325gat));
  OAI21_X1  g402(.A(G15gat), .B1(new_n589_), .B2(new_n407_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT41), .Z(new_n605_));
  INV_X1    g404(.A(G15gat), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n583_), .A2(new_n606_), .A3(new_n409_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(G1326gat));
  OAI21_X1  g407(.A(G22gat), .B1(new_n589_), .B2(new_n369_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT42), .ZN(new_n610_));
  INV_X1    g409(.A(G22gat), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n583_), .A2(new_n611_), .A3(new_n368_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(G1327gat));
  INV_X1    g412(.A(new_n587_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n484_), .A2(new_n525_), .A3(new_n540_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n414_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(G29gat), .B1(new_n617_), .B2(new_n328_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT43), .ZN(new_n619_));
  INV_X1    g418(.A(new_n581_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n414_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n412_), .B1(new_n379_), .B2(new_n407_), .ZN(new_n622_));
  OAI21_X1  g421(.A(KEYINPUT43), .B1(new_n622_), .B2(new_n581_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(new_n615_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT44), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n627_), .A2(G29gat), .A3(new_n328_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n619_), .B1(new_n414_), .B2(new_n620_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n622_), .A2(KEYINPUT43), .A3(new_n581_), .ZN(new_n630_));
  OAI211_X1 g429(.A(KEYINPUT44), .B(new_n615_), .C1(new_n629_), .C2(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n618_), .B1(new_n628_), .B2(new_n631_), .ZN(G1328gat));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n410_), .ZN(new_n633_));
  AOI21_X1  g432(.A(KEYINPUT44), .B1(new_n624_), .B2(new_n615_), .ZN(new_n634_));
  OAI21_X1  g433(.A(G36gat), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n616_), .A2(G36gat), .A3(new_n592_), .ZN(new_n636_));
  XOR2_X1   g435(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n636_), .B(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n635_), .A2(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(KEYINPUT46), .B1(new_n640_), .B2(KEYINPUT107), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT107), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT46), .ZN(new_n643_));
  AOI211_X1 g442(.A(new_n642_), .B(new_n643_), .C1(new_n635_), .C2(new_n639_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n641_), .A2(new_n644_), .ZN(G1329gat));
  INV_X1    g444(.A(G43gat), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n646_), .B1(new_n616_), .B2(new_n407_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n627_), .A2(G43gat), .A3(new_n409_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n631_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n647_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g450(.A(G50gat), .B1(new_n617_), .B2(new_n368_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n649_), .A2(new_n341_), .A3(new_n369_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n652_), .B1(new_n653_), .B2(new_n627_), .ZN(G1331gat));
  INV_X1    g453(.A(new_n484_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n655_), .A2(new_n524_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n414_), .A2(new_n540_), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(new_n587_), .ZN(new_n659_));
  INV_X1    g458(.A(G57gat), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n659_), .A2(new_n660_), .A3(new_n327_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n658_), .A2(new_n581_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT108), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(new_n328_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n661_), .B1(new_n664_), .B2(new_n660_), .ZN(G1332gat));
  OAI21_X1  g464(.A(G64gat), .B1(new_n659_), .B2(new_n592_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT48), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n592_), .A2(G64gat), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n667_), .B1(new_n662_), .B2(new_n668_), .ZN(G1333gat));
  OAI21_X1  g468(.A(G71gat), .B1(new_n659_), .B2(new_n407_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT49), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n407_), .A2(G71gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(new_n662_), .B2(new_n672_), .ZN(G1334gat));
  OAI21_X1  g472(.A(G78gat), .B1(new_n659_), .B2(new_n369_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(KEYINPUT109), .B(KEYINPUT110), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(new_n677_));
  OAI211_X1 g476(.A(G78gat), .B(new_n675_), .C1(new_n659_), .C2(new_n369_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n677_), .A2(KEYINPUT50), .A3(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(KEYINPUT50), .B1(new_n677_), .B2(new_n678_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n369_), .A2(G78gat), .ZN(new_n681_));
  OAI22_X1  g480(.A1(new_n679_), .A2(new_n680_), .B1(new_n662_), .B2(new_n681_), .ZN(G1335gat));
  NAND4_X1  g481(.A1(new_n414_), .A2(new_n541_), .A3(new_n614_), .A4(new_n656_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT111), .ZN(new_n684_));
  AOI21_X1  g483(.A(G85gat), .B1(new_n684_), .B2(new_n328_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n656_), .A2(new_n541_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(new_n621_), .B2(new_n623_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n328_), .A2(G85gat), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT112), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n685_), .B1(new_n687_), .B2(new_n689_), .ZN(G1336gat));
  NAND3_X1  g489(.A1(new_n687_), .A2(G92gat), .A3(new_n410_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n684_), .A2(new_n410_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n691_), .B1(new_n692_), .B2(G92gat), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT113), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  OAI211_X1 g494(.A(KEYINPUT113), .B(new_n691_), .C1(new_n692_), .C2(G92gat), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1337gat));
  AND2_X1   g496(.A1(new_n409_), .A2(new_n425_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n687_), .A2(new_n409_), .ZN(new_n699_));
  AOI22_X1  g498(.A1(new_n684_), .A2(new_n698_), .B1(new_n699_), .B2(G99gat), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g500(.A1(new_n684_), .A2(new_n426_), .A3(new_n368_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n426_), .B1(new_n687_), .B2(new_n368_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT52), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n703_), .A2(new_n704_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n702_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT53), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT53), .ZN(new_n709_));
  OAI211_X1 g508(.A(new_n702_), .B(new_n709_), .C1(new_n705_), .C2(new_n706_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(G1339gat));
  INV_X1    g510(.A(KEYINPUT55), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n469_), .A2(new_n457_), .A3(new_n470_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(new_n464_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n471_), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n471_), .A2(KEYINPUT55), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n715_), .A2(new_n716_), .A3(new_n476_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT56), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n478_), .B1(new_n714_), .B2(new_n471_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(KEYINPUT56), .A3(new_n716_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n485_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n506_), .A2(new_n508_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n723_), .B1(new_n485_), .B2(new_n724_), .ZN(new_n725_));
  MUX2_X1   g524(.A(new_n516_), .B(new_n725_), .S(new_n520_), .Z(new_n726_));
  NAND4_X1  g525(.A1(new_n722_), .A2(KEYINPUT58), .A3(new_n479_), .A4(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n722_), .A2(new_n479_), .A3(new_n726_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT58), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n574_), .A2(new_n580_), .A3(new_n727_), .A4(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n479_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n523_), .B2(new_n522_), .ZN(new_n733_));
  AND4_X1   g532(.A1(KEYINPUT56), .A2(new_n715_), .A3(new_n716_), .A4(new_n476_), .ZN(new_n734_));
  AOI21_X1  g533(.A(KEYINPUT56), .B1(new_n720_), .B2(new_n716_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n733_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT115), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n722_), .A2(KEYINPUT115), .A3(new_n733_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n478_), .B1(new_n467_), .B2(new_n471_), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n726_), .B(KEYINPUT116), .C1(new_n732_), .C2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(KEYINPUT116), .B1(new_n480_), .B2(new_n726_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n738_), .A2(new_n739_), .A3(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT57), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n745_), .A2(new_n746_), .A3(new_n587_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n745_), .B2(new_n587_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n731_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT117), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  OAI211_X1 g550(.A(KEYINPUT117), .B(new_n731_), .C1(new_n747_), .C2(new_n748_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(new_n541_), .A3(new_n752_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n484_), .A2(new_n541_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n581_), .A2(new_n525_), .A3(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(KEYINPUT114), .B1(new_n755_), .B2(KEYINPUT54), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(KEYINPUT54), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n524_), .B1(new_n574_), .B2(new_n580_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT114), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT54), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n758_), .A2(new_n759_), .A3(new_n760_), .A4(new_n754_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n756_), .A2(new_n757_), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n753_), .A2(new_n762_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n410_), .A2(new_n327_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n407_), .A2(new_n368_), .A3(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n763_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(G113gat), .B1(new_n768_), .B2(new_n524_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n749_), .A2(new_n541_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT118), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n749_), .A2(KEYINPUT118), .A3(new_n541_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n762_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  NOR4_X1   g573(.A1(new_n407_), .A2(KEYINPUT59), .A3(new_n765_), .A4(new_n368_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT119), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n774_), .A2(KEYINPUT119), .A3(new_n775_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n767_), .A2(KEYINPUT59), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n524_), .A2(G113gat), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n769_), .B1(new_n782_), .B2(new_n783_), .ZN(G1340gat));
  NAND3_X1  g583(.A1(new_n780_), .A2(new_n484_), .A3(new_n781_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT60), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n655_), .A2(G120gat), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n767_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(G120gat), .B1(new_n785_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n786_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(G1341gat));
  NAND4_X1  g590(.A1(new_n778_), .A2(new_n781_), .A3(new_n540_), .A4(new_n779_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(G127gat), .ZN(new_n793_));
  OR3_X1    g592(.A1(new_n767_), .A2(G127gat), .A3(new_n541_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT120), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n793_), .A2(KEYINPUT120), .A3(new_n794_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(G1342gat));
  AOI21_X1  g598(.A(G134gat), .B1(new_n768_), .B2(new_n614_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n620_), .A2(G134gat), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n782_), .B2(new_n801_), .ZN(G1343gat));
  NOR2_X1   g601(.A1(new_n409_), .A2(new_n369_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n753_), .B2(new_n762_), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT121), .B1(new_n805_), .B2(new_n764_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n805_), .A2(KEYINPUT121), .A3(new_n764_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n524_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n484_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(G148gat), .ZN(G1345gat));
  AND4_X1   g612(.A1(KEYINPUT121), .A2(new_n763_), .A3(new_n764_), .A4(new_n803_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n540_), .B1(new_n814_), .B2(new_n806_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(KEYINPUT123), .B(G155gat), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n818_));
  INV_X1    g617(.A(new_n816_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n540_), .B(new_n819_), .C1(new_n814_), .C2(new_n806_), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n817_), .A2(new_n818_), .A3(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n818_), .B1(new_n817_), .B2(new_n820_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n821_), .A2(new_n822_), .ZN(G1346gat));
  NAND2_X1  g622(.A1(new_n809_), .A2(new_n614_), .ZN(new_n824_));
  INV_X1    g623(.A(G162gat), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n824_), .A2(KEYINPUT124), .A3(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT124), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n587_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n827_), .B1(new_n828_), .B2(G162gat), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n581_), .A2(new_n825_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(KEYINPUT125), .ZN(new_n831_));
  AOI22_X1  g630(.A1(new_n826_), .A2(new_n829_), .B1(new_n809_), .B2(new_n831_), .ZN(G1347gat));
  NOR2_X1   g631(.A1(new_n592_), .A2(new_n328_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n409_), .A2(new_n833_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(KEYINPUT126), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n835_), .A2(new_n368_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n774_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n524_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(G169gat), .ZN(new_n840_));
  INV_X1    g639(.A(new_n274_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n839_), .B2(new_n841_), .ZN(new_n842_));
  MUX2_X1   g641(.A(new_n840_), .B(new_n842_), .S(KEYINPUT62), .Z(G1348gat));
  AOI21_X1  g642(.A(G176gat), .B1(new_n838_), .B2(new_n484_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n763_), .A2(new_n836_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n655_), .A2(new_n275_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n844_), .B1(new_n845_), .B2(new_n846_), .ZN(G1349gat));
  AOI21_X1  g646(.A(G183gat), .B1(new_n845_), .B2(new_n540_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n837_), .A2(new_n541_), .A3(new_n287_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n848_), .A2(new_n849_), .ZN(G1350gat));
  OAI21_X1  g649(.A(G190gat), .B1(new_n837_), .B2(new_n581_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(KEYINPUT127), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n838_), .A2(new_n257_), .A3(new_n614_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(G1351gat));
  AND2_X1   g653(.A1(new_n805_), .A2(new_n833_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n524_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n484_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g658(.A1(new_n855_), .A2(new_n540_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n861_));
  AND2_X1   g660(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n862_));
  NOR3_X1   g661(.A1(new_n860_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n863_), .B1(new_n860_), .B2(new_n861_), .ZN(G1354gat));
  AOI21_X1  g663(.A(G218gat), .B1(new_n855_), .B2(new_n614_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n620_), .A2(G218gat), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n865_), .B1(new_n855_), .B2(new_n866_), .ZN(G1355gat));
endmodule


