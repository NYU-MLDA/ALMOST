//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 0 0 0 1 0 1 1 1 1 1 0 1 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 0 1 1 1 1 0 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n917_, new_n918_, new_n919_,
    new_n921_, new_n922_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n932_, new_n933_;
  XOR2_X1   g000(.A(G15gat), .B(G22gat), .Z(new_n202_));
  NAND2_X1  g001(.A1(G1gat), .A2(G8gat), .ZN(new_n203_));
  AOI21_X1  g002(.A(new_n202_), .B1(KEYINPUT14), .B2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT76), .ZN(new_n205_));
  OR2_X1    g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n203_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G1gat), .A2(G8gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n204_), .A2(new_n205_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n206_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n209_), .B1(new_n206_), .B2(new_n210_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G231gat), .A2(G233gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT66), .B(G71gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(G78gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G57gat), .B(G64gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT11), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n219_), .A2(KEYINPUT11), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n218_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G78gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n217_), .B(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(new_n220_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n223_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n216_), .B(new_n228_), .ZN(new_n229_));
  XOR2_X1   g028(.A(G127gat), .B(G155gat), .Z(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT16), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G183gat), .B(G211gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT17), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT77), .ZN(new_n236_));
  NOR3_X1   g035(.A1(new_n233_), .A2(new_n236_), .A3(new_n234_), .ZN(new_n237_));
  OR3_X1    g036(.A1(new_n229_), .A2(new_n235_), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n229_), .A2(new_n237_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G85gat), .B(G92gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(KEYINPUT8), .B1(new_n243_), .B2(KEYINPUT64), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G99gat), .A2(G106gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT6), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(G99gat), .A2(G106gat), .ZN(new_n248_));
  XOR2_X1   g047(.A(new_n248_), .B(KEYINPUT7), .Z(new_n249_));
  OAI21_X1  g048(.A(new_n243_), .B1(new_n247_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n244_), .A2(new_n250_), .ZN(new_n251_));
  OAI221_X1 g050(.A(new_n243_), .B1(KEYINPUT64), .B2(KEYINPUT8), .C1(new_n247_), .C2(new_n249_), .ZN(new_n252_));
  XOR2_X1   g051(.A(KEYINPUT10), .B(G99gat), .Z(new_n253_));
  INV_X1    g052(.A(G106gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(G85gat), .B(G92gat), .Z(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT9), .ZN(new_n257_));
  INV_X1    g056(.A(G85gat), .ZN(new_n258_));
  INV_X1    g057(.A(G92gat), .ZN(new_n259_));
  OR3_X1    g058(.A1(new_n258_), .A2(new_n259_), .A3(KEYINPUT9), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n255_), .A2(new_n257_), .A3(new_n246_), .A4(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n251_), .A2(new_n252_), .A3(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(G29gat), .B(G36gat), .Z(new_n263_));
  XOR2_X1   g062(.A(G43gat), .B(G50gat), .Z(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n262_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT73), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G232gat), .A2(G233gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(KEYINPUT72), .B(KEYINPUT35), .Z(new_n273_));
  NOR2_X1   g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n261_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n261_), .A2(new_n276_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n251_), .A2(new_n277_), .A3(new_n252_), .A4(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n265_), .B(KEYINPUT15), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n279_), .A2(new_n280_), .B1(new_n273_), .B2(new_n272_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n268_), .A2(new_n275_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n275_), .B1(new_n268_), .B2(new_n281_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G190gat), .B(G218gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G134gat), .B(G162gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n288_), .A2(KEYINPUT36), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n285_), .A2(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(new_n288_), .B(KEYINPUT36), .Z(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT75), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n292_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n290_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(KEYINPUT74), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(KEYINPUT37), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT37), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n290_), .B(new_n293_), .C1(KEYINPUT74), .C2(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n240_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G230gat), .A2(G233gat), .ZN(new_n300_));
  INV_X1    g099(.A(new_n262_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT12), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n228_), .A2(new_n302_), .ZN(new_n303_));
  AOI22_X1  g102(.A1(new_n301_), .A2(new_n228_), .B1(new_n303_), .B2(new_n279_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n262_), .A2(new_n227_), .ZN(new_n305_));
  AOI21_X1  g104(.A(KEYINPUT68), .B1(new_n305_), .B2(new_n302_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT68), .ZN(new_n307_));
  AOI211_X1 g106(.A(new_n307_), .B(KEYINPUT12), .C1(new_n262_), .C2(new_n227_), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n300_), .B(new_n304_), .C1(new_n306_), .C2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n301_), .A2(new_n228_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(new_n305_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n311_), .A2(G230gat), .A3(G233gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  XOR2_X1   g112(.A(G120gat), .B(G148gat), .Z(new_n314_));
  XNOR2_X1  g113(.A(G176gat), .B(G204gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n316_), .B(new_n317_), .Z(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n313_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n309_), .A2(new_n312_), .A3(new_n318_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT13), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n320_), .B(new_n321_), .C1(KEYINPUT70), .C2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n299_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT78), .ZN(new_n329_));
  XOR2_X1   g128(.A(G127gat), .B(G134gat), .Z(new_n330_));
  XOR2_X1   g129(.A(G113gat), .B(G120gat), .Z(new_n331_));
  XOR2_X1   g130(.A(new_n330_), .B(new_n331_), .Z(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G71gat), .B(G99gat), .ZN(new_n334_));
  INV_X1    g133(.A(G43gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G227gat), .A2(G233gat), .ZN(new_n337_));
  INV_X1    g136(.A(G15gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n336_), .B(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G183gat), .A2(G190gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT23), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT23), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n343_), .A2(G183gat), .A3(G190gat), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT83), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n342_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n341_), .A2(KEYINPUT23), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT83), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n346_), .B(new_n348_), .C1(G183gat), .C2(G190gat), .ZN(new_n349_));
  OAI21_X1  g148(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT22), .ZN(new_n351_));
  INV_X1    g150(.A(G169gat), .ZN(new_n352_));
  INV_X1    g151(.A(G176gat), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n349_), .A2(new_n350_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT82), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G169gat), .A2(G176gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT26), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT81), .B1(new_n361_), .B2(G190gat), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT81), .ZN(new_n363_));
  INV_X1    g162(.A(G190gat), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n363_), .A2(new_n364_), .A3(KEYINPUT26), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n362_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n361_), .A2(G190gat), .ZN(new_n367_));
  INV_X1    g166(.A(G183gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT25), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT25), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(G183gat), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n367_), .A2(new_n369_), .A3(new_n371_), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n356_), .B(new_n360_), .C1(new_n366_), .C2(new_n372_), .ZN(new_n373_));
  NOR3_X1   g172(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n374_), .B1(new_n344_), .B2(new_n342_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT25), .B(G183gat), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n377_), .A2(new_n367_), .A3(new_n362_), .A4(new_n365_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n356_), .B1(new_n378_), .B2(new_n360_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n355_), .B1(new_n376_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT84), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT84), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n355_), .B(new_n382_), .C1(new_n376_), .C2(new_n379_), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n381_), .A2(KEYINPUT30), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(KEYINPUT30), .B1(new_n381_), .B2(new_n383_), .ZN(new_n385_));
  OAI21_X1  g184(.A(KEYINPUT85), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT30), .ZN(new_n387_));
  INV_X1    g186(.A(new_n383_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n360_), .B1(new_n366_), .B2(new_n372_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT82), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n390_), .A2(new_n373_), .A3(new_n375_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n382_), .B1(new_n391_), .B2(new_n355_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n387_), .B1(new_n388_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT85), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n381_), .A2(KEYINPUT30), .A3(new_n383_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n393_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n340_), .B1(new_n386_), .B2(new_n396_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n396_), .A2(new_n340_), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT31), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n340_), .ZN(new_n400_));
  NOR3_X1   g199(.A1(new_n384_), .A2(new_n385_), .A3(KEYINPUT85), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n394_), .B1(new_n393_), .B2(new_n395_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n400_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT31), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n396_), .A2(new_n340_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n403_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT86), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n399_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n407_), .B1(new_n399_), .B2(new_n406_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n333_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NOR3_X1   g209(.A1(new_n397_), .A2(new_n398_), .A3(KEYINPUT31), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n404_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT86), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n399_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(new_n332_), .A3(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G155gat), .B(G162gat), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT3), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n417_), .B1(G141gat), .B2(G148gat), .ZN(new_n418_));
  INV_X1    g217(.A(G141gat), .ZN(new_n419_));
  INV_X1    g218(.A(G148gat), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(new_n420_), .A3(KEYINPUT3), .ZN(new_n421_));
  AND3_X1   g220(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT88), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n418_), .A2(new_n421_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G141gat), .A2(G148gat), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT2), .ZN(new_n427_));
  AOI22_X1  g226(.A1(new_n425_), .A2(KEYINPUT88), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n416_), .B1(new_n424_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT89), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n419_), .A2(new_n420_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n432_), .A2(new_n426_), .A3(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n434_), .B1(KEYINPUT1), .B2(new_n416_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n435_), .B1(new_n429_), .B2(KEYINPUT89), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT90), .B1(new_n431_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT89), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n424_), .A2(new_n428_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n438_), .B1(new_n439_), .B2(new_n416_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT90), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n440_), .A2(new_n441_), .A3(new_n430_), .A4(new_n435_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n437_), .A2(new_n442_), .A3(new_n332_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n431_), .A2(new_n436_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n333_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G225gat), .A2(G233gat), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n443_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT4), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n437_), .A2(new_n442_), .A3(new_n448_), .A4(new_n332_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT98), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n443_), .A2(new_n445_), .A3(KEYINPUT4), .ZN(new_n452_));
  INV_X1    g251(.A(new_n446_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n447_), .B1(new_n451_), .B2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G1gat), .B(G29gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(G85gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT0), .B(G57gat), .ZN(new_n458_));
  XOR2_X1   g257(.A(new_n457_), .B(new_n458_), .Z(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n455_), .A2(new_n460_), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n447_), .B(new_n459_), .C1(new_n451_), .C2(new_n454_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n410_), .A2(new_n415_), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT29), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n444_), .A2(new_n466_), .ZN(new_n467_));
  OR2_X1    g266(.A1(G197gat), .A2(G204gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G197gat), .A2(G204gat), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n468_), .A2(KEYINPUT21), .A3(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G211gat), .B(G218gat), .ZN(new_n471_));
  OR2_X1    g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT21), .ZN(new_n473_));
  INV_X1    g272(.A(new_n469_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(G197gat), .A2(G204gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n473_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n476_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n472_), .A2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT92), .ZN(new_n479_));
  OAI211_X1 g278(.A(G228gat), .B(G233gat), .C1(new_n467_), .C2(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n478_), .B1(G228gat), .B2(G233gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n437_), .A2(new_n442_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n481_), .B1(new_n482_), .B2(new_n466_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n480_), .A2(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(G78gat), .B(G106gat), .Z(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n485_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n480_), .A2(new_n483_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G22gat), .B(G50gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n490_), .B(KEYINPUT91), .Z(new_n491_));
  INV_X1    g290(.A(KEYINPUT28), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n482_), .A2(new_n492_), .A3(new_n466_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n492_), .B1(new_n482_), .B2(new_n466_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n491_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n495_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n491_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n497_), .A2(new_n493_), .A3(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n496_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n489_), .A2(new_n500_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n486_), .A2(new_n496_), .A3(new_n499_), .A4(new_n488_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G8gat), .B(G36gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT18), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G64gat), .B(G92gat), .ZN(new_n506_));
  XOR2_X1   g305(.A(new_n505_), .B(new_n506_), .Z(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n381_), .A2(new_n478_), .A3(new_n383_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT20), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n374_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n364_), .A2(KEYINPUT26), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n367_), .A2(new_n369_), .A3(new_n371_), .A4(new_n512_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n511_), .A2(new_n346_), .A3(new_n348_), .A4(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n343_), .B1(G183gat), .B2(G190gat), .ZN(new_n515_));
  OAI22_X1  g314(.A1(new_n515_), .A2(new_n347_), .B1(G183gat), .B2(G190gat), .ZN(new_n516_));
  INV_X1    g315(.A(new_n350_), .ZN(new_n517_));
  NOR3_X1   g316(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n518_));
  OAI21_X1  g317(.A(KEYINPUT94), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT94), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n354_), .A2(new_n520_), .A3(new_n350_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n516_), .A2(new_n519_), .A3(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n514_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n472_), .A2(new_n477_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n510_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n509_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G226gat), .A2(G233gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n526_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n529_), .ZN(new_n531_));
  XOR2_X1   g330(.A(KEYINPUT100), .B(KEYINPUT20), .Z(new_n532_));
  INV_X1    g331(.A(new_n523_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n532_), .B1(new_n479_), .B2(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n524_), .B1(new_n388_), .B2(new_n392_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n531_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n508_), .B1(new_n530_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n526_), .A2(new_n529_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n478_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT95), .B1(new_n523_), .B2(new_n524_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT95), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n478_), .A2(new_n541_), .A3(new_n514_), .A4(new_n522_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n529_), .A2(new_n510_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT96), .B1(new_n539_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT96), .ZN(new_n547_));
  INV_X1    g346(.A(new_n544_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n548_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n535_), .A2(new_n547_), .A3(new_n549_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n538_), .A2(new_n546_), .A3(new_n550_), .A4(new_n507_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n537_), .A2(KEYINPUT27), .A3(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT101), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n539_), .A2(new_n545_), .ZN(new_n554_));
  AOI22_X1  g353(.A1(new_n554_), .A2(new_n547_), .B1(new_n526_), .B2(new_n529_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n555_), .A2(KEYINPUT97), .A3(new_n507_), .A4(new_n546_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT97), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n551_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n538_), .A2(new_n546_), .A3(new_n550_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(new_n508_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n556_), .A2(new_n558_), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT103), .ZN(new_n562_));
  XOR2_X1   g361(.A(KEYINPUT102), .B(KEYINPUT27), .Z(new_n563_));
  AND3_X1   g362(.A1(new_n561_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n562_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n503_), .B(new_n553_), .C1(new_n564_), .C2(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n465_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT87), .ZN(new_n568_));
  NOR3_X1   g367(.A1(new_n408_), .A2(new_n409_), .A3(new_n333_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n332_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n568_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n410_), .A2(new_n415_), .A3(KEYINPUT87), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n530_), .A2(new_n536_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n507_), .A2(KEYINPUT32), .ZN(new_n575_));
  MUX2_X1   g374(.A(new_n574_), .B(new_n559_), .S(new_n575_), .Z(new_n576_));
  NAND2_X1  g375(.A1(new_n463_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT33), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n462_), .A2(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n449_), .B(KEYINPUT98), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n580_), .A2(new_n453_), .A3(new_n452_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n581_), .A2(KEYINPUT33), .A3(new_n447_), .A4(new_n459_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n443_), .A2(new_n445_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n460_), .B1(new_n583_), .B2(new_n446_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n584_), .A2(KEYINPUT99), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n580_), .A2(new_n446_), .A3(new_n452_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(KEYINPUT99), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n579_), .B(new_n582_), .C1(new_n585_), .C2(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n577_), .B1(new_n589_), .B2(new_n561_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(new_n503_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n503_), .A2(new_n463_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n592_), .B(new_n553_), .C1(new_n564_), .C2(new_n565_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n567_), .B1(new_n573_), .B2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n266_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n213_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n597_), .A2(new_n265_), .A3(new_n211_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT79), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n596_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  OAI211_X1 g399(.A(KEYINPUT79), .B(new_n266_), .C1(new_n212_), .C2(new_n213_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT80), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G229gat), .A2(G233gat), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n600_), .A2(new_n601_), .A3(new_n602_), .A4(new_n604_), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n600_), .A2(new_n601_), .A3(new_n604_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n280_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(new_n598_), .ZN(new_n608_));
  OAI21_X1  g407(.A(KEYINPUT80), .B1(new_n608_), .B2(new_n604_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n605_), .B1(new_n606_), .B2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G113gat), .B(G141gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G169gat), .B(G197gat), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n611_), .B(new_n612_), .Z(new_n613_));
  OR2_X1    g412(.A1(new_n610_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n610_), .A2(new_n613_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n595_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n329_), .A2(new_n618_), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n619_), .A2(G1gat), .A3(new_n464_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT38), .Z(new_n621_));
  XNOR2_X1  g420(.A(new_n294_), .B(KEYINPUT104), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n595_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n327_), .A2(new_n616_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n624_), .A2(new_n240_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G1gat), .B1(new_n626_), .B2(new_n464_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(KEYINPUT105), .Z(new_n628_));
  NAND2_X1  g427(.A1(new_n621_), .A2(new_n628_), .ZN(G1324gat));
  OR2_X1    g428(.A1(new_n564_), .A2(new_n565_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(new_n553_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  OR3_X1    g431(.A1(new_n619_), .A2(G8gat), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT39), .ZN(new_n634_));
  INV_X1    g433(.A(new_n625_), .ZN(new_n635_));
  NOR4_X1   g434(.A1(new_n595_), .A2(new_n635_), .A3(new_n632_), .A4(new_n622_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT106), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n637_), .A2(G8gat), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n636_), .A2(KEYINPUT106), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n634_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  AND4_X1   g439(.A1(new_n634_), .A2(new_n639_), .A3(G8gat), .A4(new_n637_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n633_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT40), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  OAI211_X1 g443(.A(KEYINPUT40), .B(new_n633_), .C1(new_n640_), .C2(new_n641_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(G1325gat));
  NOR3_X1   g445(.A1(new_n619_), .A2(G15gat), .A3(new_n573_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT107), .Z(new_n648_));
  INV_X1    g447(.A(new_n626_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n573_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n338_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT41), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n652_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n648_), .A2(new_n653_), .A3(new_n654_), .ZN(G1326gat));
  INV_X1    g454(.A(G22gat), .ZN(new_n656_));
  INV_X1    g455(.A(new_n503_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n329_), .A2(new_n656_), .A3(new_n657_), .A4(new_n618_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT42), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n649_), .A2(new_n657_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n660_), .B2(G22gat), .ZN(new_n661_));
  AOI211_X1 g460(.A(KEYINPUT42), .B(new_n656_), .C1(new_n649_), .C2(new_n657_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n658_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT108), .ZN(G1327gat));
  INV_X1    g463(.A(new_n327_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n240_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n665_), .A2(new_n666_), .A3(new_n294_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n618_), .A2(new_n667_), .ZN(new_n668_));
  OR3_X1    g467(.A1(new_n668_), .A2(G29gat), .A3(new_n464_), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n296_), .A2(KEYINPUT109), .A3(new_n298_), .ZN(new_n670_));
  AOI21_X1  g469(.A(KEYINPUT109), .B1(new_n296_), .B2(new_n298_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(KEYINPUT43), .B1(new_n595_), .B2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n296_), .A2(new_n298_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n674_), .A2(KEYINPUT43), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(KEYINPUT110), .B1(new_n595_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT110), .ZN(new_n678_));
  AOI22_X1  g477(.A1(new_n571_), .A2(new_n572_), .B1(new_n591_), .B2(new_n593_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n678_), .B(new_n675_), .C1(new_n679_), .C2(new_n567_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n673_), .A2(new_n677_), .A3(new_n680_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n624_), .A2(new_n666_), .ZN(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT44), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n681_), .A2(KEYINPUT44), .A3(new_n682_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n684_), .A2(new_n463_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT111), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n686_), .A2(new_n687_), .A3(G29gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n686_), .B2(G29gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n669_), .B1(new_n688_), .B2(new_n689_), .ZN(G1328gat));
  INV_X1    g489(.A(G36gat), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n618_), .A2(new_n691_), .A3(new_n631_), .A4(new_n667_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT45), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n681_), .A2(KEYINPUT44), .A3(new_n682_), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n694_), .A2(new_n683_), .A3(new_n632_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n693_), .B1(new_n695_), .B2(new_n691_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT46), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  OAI211_X1 g497(.A(KEYINPUT46), .B(new_n693_), .C1(new_n695_), .C2(new_n691_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1329gat));
  NOR2_X1   g499(.A1(new_n569_), .A2(new_n570_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(G43gat), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n694_), .A2(new_n683_), .A3(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT47), .ZN(new_n705_));
  INV_X1    g504(.A(new_n668_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(new_n650_), .ZN(new_n707_));
  AOI21_X1  g506(.A(KEYINPUT112), .B1(new_n707_), .B2(new_n335_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT112), .ZN(new_n709_));
  AOI211_X1 g508(.A(new_n709_), .B(G43gat), .C1(new_n706_), .C2(new_n650_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n704_), .B(new_n705_), .C1(new_n708_), .C2(new_n710_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n708_), .A2(new_n710_), .ZN(new_n712_));
  OAI21_X1  g511(.A(KEYINPUT47), .B1(new_n712_), .B2(new_n703_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1330gat));
  AOI21_X1  g513(.A(G50gat), .B1(new_n706_), .B2(new_n657_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n694_), .A2(new_n683_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n657_), .A2(G50gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n715_), .B1(new_n716_), .B2(new_n717_), .ZN(G1331gat));
  INV_X1    g517(.A(new_n623_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n665_), .A2(new_n617_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n719_), .A2(new_n240_), .A3(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(G57gat), .B1(new_n722_), .B2(new_n464_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n299_), .A2(new_n665_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT113), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n725_), .A2(new_n595_), .A3(new_n616_), .ZN(new_n726_));
  INV_X1    g525(.A(G57gat), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n726_), .A2(new_n727_), .A3(new_n463_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n723_), .A2(new_n728_), .ZN(G1332gat));
  INV_X1    g528(.A(G64gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n730_), .B1(new_n721_), .B2(new_n631_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT48), .Z(new_n732_));
  NAND2_X1  g531(.A1(new_n631_), .A2(new_n730_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT114), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n726_), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n732_), .A2(new_n735_), .ZN(G1333gat));
  INV_X1    g535(.A(G71gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n721_), .B2(new_n650_), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT49), .Z(new_n739_));
  NAND3_X1  g538(.A1(new_n726_), .A2(new_n737_), .A3(new_n650_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1334gat));
  AOI21_X1  g540(.A(new_n224_), .B1(new_n721_), .B2(new_n657_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT50), .Z(new_n743_));
  NAND3_X1  g542(.A1(new_n726_), .A2(new_n224_), .A3(new_n657_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1335gat));
  INV_X1    g544(.A(new_n292_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n268_), .A2(new_n281_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(new_n274_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n746_), .B1(new_n748_), .B2(new_n282_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n289_), .B2(new_n285_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n665_), .A2(new_n750_), .A3(new_n240_), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n595_), .A2(new_n616_), .A3(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n752_), .A2(new_n258_), .A3(new_n463_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n720_), .A2(new_n666_), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n681_), .A2(new_n463_), .A3(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n753_), .B1(new_n755_), .B2(new_n258_), .ZN(G1336gat));
  NAND3_X1  g555(.A1(new_n752_), .A2(new_n259_), .A3(new_n631_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n681_), .A2(new_n631_), .A3(new_n754_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n758_), .B2(new_n259_), .ZN(G1337gat));
  NAND3_X1  g558(.A1(new_n681_), .A2(new_n650_), .A3(new_n754_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(G99gat), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n701_), .A2(new_n253_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT115), .ZN(new_n763_));
  AOI22_X1  g562(.A1(new_n752_), .A2(new_n762_), .B1(new_n763_), .B2(KEYINPUT51), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n761_), .A2(new_n764_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n763_), .A2(KEYINPUT51), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n765_), .B(new_n766_), .Z(G1338gat));
  NAND3_X1  g566(.A1(new_n752_), .A2(new_n254_), .A3(new_n657_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n681_), .A2(new_n657_), .A3(new_n754_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n769_), .A2(new_n770_), .A3(G106gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n769_), .B2(G106gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT53), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n775_), .B(new_n768_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1339gat));
  INV_X1    g576(.A(new_n321_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n778_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n309_), .A2(KEYINPUT117), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT55), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n309_), .A2(KEYINPUT117), .A3(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT118), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n303_), .A2(new_n279_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n310_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n305_), .A2(new_n302_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n307_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n305_), .A2(KEYINPUT68), .A3(new_n302_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n786_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n784_), .B1(new_n790_), .B2(new_n300_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n304_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n792_), .A2(KEYINPUT118), .A3(G230gat), .A4(G233gat), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n781_), .A2(new_n783_), .A3(new_n791_), .A4(new_n793_), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n794_), .A2(KEYINPUT56), .A3(new_n319_), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT56), .B1(new_n794_), .B2(new_n319_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n779_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT119), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n603_), .B1(new_n608_), .B2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n799_), .B1(new_n798_), .B2(new_n608_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n613_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n600_), .A2(new_n601_), .A3(new_n603_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n800_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n322_), .A2(new_n615_), .A3(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n750_), .B1(new_n797_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT120), .ZN(new_n806_));
  OAI21_X1  g605(.A(KEYINPUT57), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808_));
  INV_X1    g607(.A(new_n804_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n794_), .A2(new_n319_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT56), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n794_), .A2(KEYINPUT56), .A3(new_n319_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n809_), .B1(new_n814_), .B2(new_n779_), .ZN(new_n815_));
  OAI211_X1 g614(.A(KEYINPUT120), .B(new_n808_), .C1(new_n815_), .C2(new_n750_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n615_), .A2(new_n321_), .A3(new_n803_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT121), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT121), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n615_), .A2(new_n819_), .A3(new_n321_), .A4(new_n803_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n821_), .B1(new_n796_), .B2(new_n795_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT58), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n674_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n814_), .A2(KEYINPUT58), .A3(new_n821_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n824_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n807_), .A2(new_n816_), .A3(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n240_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n674_), .A2(new_n666_), .A3(new_n617_), .A4(new_n327_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT116), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n831_), .A2(KEYINPUT54), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n299_), .A2(new_n617_), .A3(new_n327_), .A4(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n829_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT122), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n836_), .B1(new_n828_), .B2(new_n240_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT122), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n839_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(G113gat), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n701_), .A2(new_n463_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n845_), .A2(new_n566_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n843_), .A2(new_n844_), .A3(new_n616_), .A4(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n846_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n840_), .A2(KEYINPUT59), .A3(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n841_), .B1(new_n829_), .B2(new_n837_), .ZN(new_n850_));
  AOI211_X1 g649(.A(KEYINPUT122), .B(new_n836_), .C1(new_n828_), .C2(new_n240_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n846_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  AOI211_X1 g651(.A(new_n617_), .B(new_n849_), .C1(new_n852_), .C2(KEYINPUT59), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n847_), .B1(new_n853_), .B2(new_n844_), .ZN(G1340gat));
  INV_X1    g653(.A(G120gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n327_), .B2(KEYINPUT60), .ZN(new_n856_));
  OR2_X1    g655(.A1(new_n855_), .A2(KEYINPUT60), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n843_), .A2(new_n846_), .A3(new_n856_), .A4(new_n857_), .ZN(new_n858_));
  AOI211_X1 g657(.A(new_n327_), .B(new_n849_), .C1(new_n852_), .C2(KEYINPUT59), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n859_), .B2(new_n855_), .ZN(G1341gat));
  OAI211_X1 g659(.A(new_n666_), .B(new_n846_), .C1(new_n850_), .C2(new_n851_), .ZN(new_n861_));
  INV_X1    g660(.A(G127gat), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT123), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT123), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n861_), .A2(new_n865_), .A3(new_n862_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n849_), .B1(new_n852_), .B2(KEYINPUT59), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n240_), .A2(new_n862_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(KEYINPUT124), .ZN(new_n869_));
  AOI22_X1  g668(.A1(new_n864_), .A2(new_n866_), .B1(new_n867_), .B2(new_n869_), .ZN(G1342gat));
  INV_X1    g669(.A(G134gat), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n843_), .A2(new_n871_), .A3(new_n622_), .A4(new_n846_), .ZN(new_n872_));
  AOI211_X1 g671(.A(new_n674_), .B(new_n849_), .C1(new_n852_), .C2(KEYINPUT59), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(new_n871_), .ZN(G1343gat));
  NOR2_X1   g673(.A1(new_n650_), .A2(new_n503_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n875_), .A2(new_n463_), .A3(new_n632_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n843_), .A2(new_n616_), .A3(new_n877_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g678(.A1(new_n843_), .A2(new_n665_), .A3(new_n877_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g680(.A1(new_n843_), .A2(new_n666_), .A3(new_n877_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT61), .B(G155gat), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1346gat));
  AOI21_X1  g683(.A(new_n876_), .B1(new_n839_), .B2(new_n842_), .ZN(new_n885_));
  AOI21_X1  g684(.A(G162gat), .B1(new_n885_), .B2(new_n622_), .ZN(new_n886_));
  INV_X1    g685(.A(G162gat), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n672_), .A2(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n886_), .B1(new_n885_), .B2(new_n888_), .ZN(G1347gat));
  NOR2_X1   g688(.A1(new_n632_), .A2(new_n463_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n890_), .A2(new_n503_), .A3(new_n650_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n840_), .A2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(KEYINPUT125), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT125), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n894_), .B1(new_n840_), .B2(new_n891_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n893_), .A2(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n351_), .A2(new_n352_), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n896_), .B(new_n616_), .C1(new_n897_), .C2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT62), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n892_), .A2(new_n616_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(G169gat), .ZN(new_n902_));
  AOI211_X1 g701(.A(KEYINPUT62), .B(new_n352_), .C1(new_n892_), .C2(new_n616_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n899_), .B1(new_n902_), .B2(new_n903_), .ZN(G1348gat));
  AOI21_X1  g703(.A(G176gat), .B1(new_n896_), .B2(new_n665_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n657_), .B1(new_n839_), .B2(new_n842_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n890_), .A2(new_n650_), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n907_), .A2(new_n353_), .A3(new_n327_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n905_), .B1(new_n906_), .B2(new_n908_), .ZN(G1349gat));
  NOR2_X1   g708(.A1(new_n907_), .A2(new_n240_), .ZN(new_n910_));
  AOI21_X1  g709(.A(G183gat), .B1(new_n906_), .B2(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n240_), .A2(new_n377_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n911_), .B1(new_n896_), .B2(new_n912_), .ZN(G1350gat));
  NAND4_X1  g712(.A1(new_n896_), .A2(new_n367_), .A3(new_n512_), .A4(new_n622_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n674_), .B1(new_n893_), .B2(new_n895_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n915_), .B2(new_n364_), .ZN(G1351gat));
  NAND2_X1  g715(.A1(new_n875_), .A2(new_n890_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n843_), .A2(new_n616_), .A3(new_n918_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g719(.A1(new_n843_), .A2(new_n665_), .A3(new_n918_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n921_), .B1(KEYINPUT126), .B2(G204gat), .ZN(new_n922_));
  XOR2_X1   g721(.A(KEYINPUT126), .B(G204gat), .Z(new_n923_));
  OAI21_X1  g722(.A(new_n922_), .B1(new_n921_), .B2(new_n923_), .ZN(G1353gat));
  AOI21_X1  g723(.A(new_n240_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n843_), .A2(new_n918_), .A3(new_n925_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n927_));
  XOR2_X1   g726(.A(new_n927_), .B(KEYINPUT127), .Z(new_n928_));
  XNOR2_X1  g727(.A(new_n926_), .B(new_n928_), .ZN(G1354gat));
  NAND2_X1  g728(.A1(new_n843_), .A2(new_n918_), .ZN(new_n930_));
  OAI21_X1  g729(.A(G218gat), .B1(new_n930_), .B2(new_n674_), .ZN(new_n931_));
  INV_X1    g730(.A(G218gat), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n622_), .A2(new_n932_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n931_), .B1(new_n930_), .B2(new_n933_), .ZN(G1355gat));
endmodule


