//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 0 0 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n961_, new_n962_, new_n963_, new_n964_, new_n965_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n987_, new_n988_,
    new_n990_, new_n991_, new_n992_, new_n994_, new_n995_, new_n997_,
    new_n998_, new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_,
    new_n1004_, new_n1006_, new_n1007_, new_n1008_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1015_, new_n1016_;
  XNOR2_X1  g000(.A(KEYINPUT99), .B(KEYINPUT27), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G226gat), .A2(G233gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT19), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT83), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207_));
  INV_X1    g006(.A(G176gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT81), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT81), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G176gat), .ZN(new_n211_));
  INV_X1    g010(.A(G169gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT22), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT22), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(G169gat), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n209_), .A2(new_n211_), .A3(new_n213_), .A4(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n207_), .B1(new_n216_), .B2(KEYINPUT82), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT82), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT81), .B(G176gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT22), .B(G169gat), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n218_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n206_), .B1(new_n217_), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT23), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n225_), .A2(G183gat), .A3(G190gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT84), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n224_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(G183gat), .ZN(new_n229_));
  INV_X1    g028(.A(G190gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n225_), .A2(KEYINPUT84), .A3(G183gat), .A4(G190gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n228_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n216_), .A2(KEYINPUT82), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n219_), .A2(new_n220_), .A3(new_n218_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n234_), .A2(KEYINPUT83), .A3(new_n207_), .A4(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n222_), .A2(new_n233_), .A3(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT21), .ZN(new_n238_));
  INV_X1    g037(.A(G218gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(G211gat), .ZN(new_n240_));
  INV_X1    g039(.A(G211gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(G218gat), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n238_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT90), .ZN(new_n244_));
  INV_X1    g043(.A(G204gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(KEYINPUT90), .A2(G204gat), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n246_), .A2(G197gat), .A3(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT91), .B1(new_n245_), .B2(G197gat), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT91), .ZN(new_n250_));
  INV_X1    g049(.A(G197gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(new_n251_), .A3(G204gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n249_), .A2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n243_), .B1(new_n248_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT92), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  OAI211_X1 g055(.A(KEYINPUT92), .B(new_n243_), .C1(new_n248_), .C2(new_n253_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n246_), .A2(G197gat), .A3(new_n247_), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n258_), .A2(new_n238_), .A3(new_n252_), .A4(new_n249_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n240_), .A2(new_n242_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n246_), .A2(new_n251_), .A3(new_n247_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n238_), .B1(G197gat), .B2(G204gat), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n260_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  AOI22_X1  g062(.A1(new_n256_), .A2(new_n257_), .B1(new_n259_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n229_), .A2(KEYINPUT25), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT25), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(G183gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n230_), .A2(KEYINPUT26), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT26), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(G190gat), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n265_), .A2(new_n267_), .A3(new_n268_), .A4(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n212_), .A2(new_n208_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n272_), .A2(KEYINPUT24), .A3(new_n207_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n224_), .A2(new_n226_), .ZN(new_n276_));
  OR3_X1    g075(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n237_), .A2(new_n264_), .A3(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT95), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n228_), .A2(new_n232_), .A3(new_n277_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n274_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n228_), .A2(KEYINPUT95), .A3(new_n232_), .A4(new_n277_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT96), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n220_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n220_), .A2(new_n284_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n285_), .A2(new_n286_), .A3(new_n219_), .ZN(new_n287_));
  AOI22_X1  g086(.A1(new_n276_), .A2(new_n231_), .B1(G169gat), .B2(G176gat), .ZN(new_n288_));
  AOI22_X1  g087(.A1(new_n282_), .A2(new_n283_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT20), .B1(new_n289_), .B2(new_n264_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n205_), .B1(new_n279_), .B2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G8gat), .B(G36gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT18), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G64gat), .B(G92gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n237_), .A2(new_n278_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n263_), .A2(new_n259_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n257_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n258_), .A2(new_n252_), .A3(new_n249_), .ZN(new_n300_));
  AOI21_X1  g099(.A(KEYINPUT92), .B1(new_n300_), .B2(new_n243_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n298_), .B1(new_n299_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n205_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT20), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n305_), .B1(new_n289_), .B2(new_n264_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n303_), .A2(new_n304_), .A3(new_n306_), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n291_), .A2(new_n296_), .A3(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n296_), .B1(new_n291_), .B2(new_n307_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n203_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n264_), .B1(new_n237_), .B2(new_n278_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n281_), .A2(new_n280_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n312_), .A2(new_n275_), .A3(new_n283_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n287_), .A2(new_n288_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT20), .B1(new_n315_), .B2(new_n302_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n205_), .B1(new_n311_), .B2(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n305_), .B1(new_n315_), .B2(new_n302_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n237_), .A2(new_n264_), .A3(new_n278_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n318_), .A2(new_n319_), .A3(new_n304_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n317_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(new_n295_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n291_), .A2(new_n307_), .A3(new_n296_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n322_), .A2(KEYINPUT27), .A3(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n310_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT29), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT3), .ZN(new_n327_));
  INV_X1    g126(.A(G141gat), .ZN(new_n328_));
  INV_X1    g127(.A(G148gat), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .A4(KEYINPUT89), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT89), .ZN(new_n331_));
  OAI22_X1  g130(.A1(new_n331_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G141gat), .A2(G148gat), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT2), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n330_), .A2(new_n332_), .A3(new_n335_), .A4(new_n336_), .ZN(new_n337_));
  XOR2_X1   g136(.A(G155gat), .B(G162gat), .Z(new_n338_));
  INV_X1    g137(.A(G155gat), .ZN(new_n339_));
  INV_X1    g138(.A(G162gat), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT1), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT1), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(G155gat), .A3(G162gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n339_), .A2(new_n340_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n341_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  XOR2_X1   g144(.A(G141gat), .B(G148gat), .Z(new_n346_));
  AOI22_X1  g145(.A1(new_n337_), .A2(new_n338_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n302_), .B1(new_n326_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G78gat), .B(G106gat), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT93), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n302_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G228gat), .A2(G233gat), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n350_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n350_), .ZN(new_n356_));
  AOI211_X1 g155(.A(new_n353_), .B(new_n356_), .C1(new_n302_), .C2(new_n351_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n349_), .B1(new_n355_), .B2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G22gat), .B(G50gat), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n337_), .A2(new_n338_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n345_), .A2(new_n346_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n361_), .A2(new_n326_), .A3(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n363_), .A2(KEYINPUT28), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT28), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n365_), .B1(new_n347_), .B2(new_n326_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n360_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n363_), .A2(KEYINPUT28), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n347_), .A2(new_n365_), .A3(new_n326_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(new_n369_), .A3(new_n359_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n367_), .A2(KEYINPUT94), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n256_), .A2(new_n257_), .ZN(new_n373_));
  AOI21_X1  g172(.A(KEYINPUT93), .B1(new_n373_), .B2(new_n298_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n356_), .B1(new_n374_), .B2(new_n353_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n352_), .A2(new_n354_), .A3(new_n350_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(new_n348_), .A3(new_n376_), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n358_), .A2(new_n372_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT94), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n368_), .A2(new_n369_), .A3(new_n359_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n359_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n379_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(new_n371_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n383_), .B1(new_n358_), .B2(new_n377_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n378_), .A2(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n325_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G227gat), .A2(G233gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(G15gat), .ZN(new_n388_));
  INV_X1    g187(.A(G43gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G71gat), .B(G99gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n237_), .A2(KEYINPUT30), .A3(new_n278_), .ZN(new_n394_));
  AOI21_X1  g193(.A(KEYINPUT30), .B1(new_n237_), .B2(new_n278_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n393_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT30), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n297_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n237_), .A2(KEYINPUT30), .A3(new_n278_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n398_), .A2(new_n399_), .A3(new_n392_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT85), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n396_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G113gat), .B(G120gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(G134gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(G127gat), .ZN(new_n406_));
  INV_X1    g205(.A(G127gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(G134gat), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n406_), .A2(new_n408_), .A3(KEYINPUT86), .ZN(new_n409_));
  AOI21_X1  g208(.A(KEYINPUT86), .B1(new_n406_), .B2(new_n408_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n404_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT86), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n407_), .A2(G134gat), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n405_), .A2(G127gat), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n412_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n406_), .A2(new_n408_), .A3(KEYINPUT86), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n415_), .A2(new_n416_), .A3(new_n403_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n411_), .A2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT31), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n402_), .A2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n401_), .B1(new_n396_), .B2(new_n400_), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT87), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n400_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n392_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT85), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT87), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n426_), .A2(new_n427_), .A3(new_n420_), .A4(new_n402_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n396_), .A2(new_n400_), .A3(new_n419_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n423_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G1gat), .B(G29gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(G85gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT0), .B(G57gat), .ZN(new_n433_));
  XOR2_X1   g232(.A(new_n432_), .B(new_n433_), .Z(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n361_), .A2(new_n362_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT4), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n418_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G225gat), .A2(G233gat), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n438_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n418_), .A2(new_n436_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT97), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n411_), .A2(new_n361_), .A3(new_n417_), .A4(new_n362_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n347_), .A2(KEYINPUT97), .A3(new_n417_), .A4(new_n411_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n441_), .B1(new_n447_), .B2(KEYINPUT4), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n440_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n435_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n447_), .A2(new_n439_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n437_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n451_), .B(new_n434_), .C1(new_n452_), .C2(new_n441_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n450_), .A2(KEYINPUT98), .A3(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT98), .ZN(new_n455_));
  OAI211_X1 g254(.A(new_n455_), .B(new_n435_), .C1(new_n448_), .C2(new_n449_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n386_), .A2(new_n430_), .A3(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT88), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n430_), .A2(new_n459_), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n423_), .A2(new_n428_), .A3(KEYINPUT88), .A4(new_n429_), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n323_), .A2(KEYINPUT27), .ZN(new_n463_));
  NOR3_X1   g262(.A1(new_n311_), .A2(new_n316_), .A3(new_n205_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n304_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n295_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n323_), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n463_), .A2(new_n322_), .B1(new_n467_), .B2(new_n203_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT100), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n468_), .A2(new_n469_), .A3(new_n457_), .A4(new_n385_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n385_), .A2(new_n457_), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT100), .B1(new_n471_), .B2(new_n325_), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n296_), .A2(KEYINPUT32), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n317_), .A2(new_n320_), .A3(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n473_), .B1(new_n291_), .B2(new_n307_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT33), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n453_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n447_), .A2(KEYINPUT4), .ZN(new_n479_));
  INV_X1    g278(.A(new_n441_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n481_), .A2(KEYINPUT33), .A3(new_n451_), .A4(new_n434_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n434_), .B1(new_n447_), .B2(new_n440_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n438_), .A2(new_n439_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n483_), .B1(new_n452_), .B2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n478_), .A2(new_n482_), .A3(new_n485_), .ZN(new_n486_));
  OAI22_X1  g285(.A1(new_n457_), .A2(new_n476_), .B1(new_n486_), .B2(new_n467_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n385_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n470_), .A2(new_n472_), .A3(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n458_), .B1(new_n462_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT79), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT75), .B(G8gat), .ZN(new_n493_));
  INV_X1    g292(.A(G1gat), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT14), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT76), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G15gat), .B(G22gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G1gat), .B(G8gat), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n497_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n499_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G29gat), .B(G36gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT72), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G43gat), .B(G50gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n492_), .B1(new_n502_), .B2(new_n506_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n504_), .A2(new_n505_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n504_), .A2(new_n505_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  OAI211_X1 g309(.A(KEYINPUT79), .B(new_n510_), .C1(new_n500_), .C2(new_n501_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n507_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G229gat), .A2(G233gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT80), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n510_), .A2(KEYINPUT15), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT15), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n506_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n515_), .B1(new_n519_), .B2(new_n502_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n512_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G113gat), .B(G141gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G169gat), .B(G197gat), .ZN(new_n523_));
  XOR2_X1   g322(.A(new_n522_), .B(new_n523_), .Z(new_n524_));
  NAND2_X1  g323(.A1(new_n502_), .A2(new_n506_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n512_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n521_), .B(new_n524_), .C1(new_n527_), .C2(new_n513_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n524_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n521_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n513_), .B1(new_n512_), .B2(new_n525_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n529_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  AND2_X1   g331(.A1(new_n528_), .A2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n491_), .A2(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT78), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G127gat), .B(G155gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G183gat), .B(G211gat), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n538_), .B(new_n539_), .Z(new_n540_));
  XOR2_X1   g339(.A(new_n540_), .B(KEYINPUT17), .Z(new_n541_));
  NAND2_X1  g340(.A1(G231gat), .A2(G233gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n502_), .B(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G71gat), .B(G78gat), .ZN(new_n544_));
  INV_X1    g343(.A(G64gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(G57gat), .ZN(new_n546_));
  INV_X1    g345(.A(G57gat), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(G64gat), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n546_), .A2(new_n548_), .A3(KEYINPUT67), .ZN(new_n549_));
  AOI21_X1  g348(.A(KEYINPUT67), .B1(new_n546_), .B2(new_n548_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT11), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n544_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT11), .B1(new_n549_), .B2(new_n550_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT68), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT67), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n547_), .A2(G64gat), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n545_), .A2(G57gat), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n556_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n546_), .A2(new_n548_), .A3(KEYINPUT67), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT68), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n561_), .A2(new_n562_), .A3(KEYINPUT11), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n553_), .A2(new_n555_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n553_), .B1(new_n555_), .B2(new_n563_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n543_), .A2(new_n567_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n543_), .A2(new_n567_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n541_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n554_), .A2(KEYINPUT68), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n562_), .B1(new_n561_), .B2(KEYINPUT11), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n561_), .A2(KEYINPUT11), .ZN(new_n573_));
  OAI22_X1  g372(.A1(new_n571_), .A2(new_n572_), .B1(new_n573_), .B2(new_n544_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n574_), .A2(KEYINPUT70), .A3(new_n564_), .ZN(new_n575_));
  AOI21_X1  g374(.A(KEYINPUT70), .B1(new_n574_), .B2(new_n564_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n543_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n543_), .A2(new_n577_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n578_), .A2(KEYINPUT17), .A3(new_n540_), .A4(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n570_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT66), .ZN(new_n582_));
  OAI22_X1  g381(.A1(new_n582_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT7), .ZN(new_n584_));
  INV_X1    g383(.A(G99gat), .ZN(new_n585_));
  INV_X1    g384(.A(G106gat), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n584_), .A2(new_n585_), .A3(new_n586_), .A4(KEYINPUT66), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G99gat), .A2(G106gat), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n588_), .A2(KEYINPUT6), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n588_), .A2(KEYINPUT6), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n583_), .B(new_n587_), .C1(new_n589_), .C2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(G85gat), .ZN(new_n592_));
  INV_X1    g391(.A(G92gat), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G85gat), .A2(G92gat), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(KEYINPUT8), .B1(new_n591_), .B2(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n588_), .B(KEYINPUT6), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT9), .ZN(new_n599_));
  INV_X1    g398(.A(new_n595_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT65), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n599_), .B(new_n594_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n602_));
  OR2_X1    g401(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n586_), .A2(KEYINPUT64), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT64), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(G106gat), .ZN(new_n606_));
  NAND2_X1  g405(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n603_), .A2(new_n604_), .A3(new_n606_), .A4(new_n607_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n594_), .A2(KEYINPUT65), .A3(KEYINPUT9), .A4(new_n595_), .ZN(new_n609_));
  AND4_X1   g408(.A1(new_n598_), .A2(new_n602_), .A3(new_n608_), .A4(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n597_), .A2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n591_), .A2(KEYINPUT8), .A3(new_n596_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(G232gat), .A2(G233gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT34), .ZN(new_n615_));
  OAI22_X1  g414(.A1(new_n613_), .A2(new_n506_), .B1(KEYINPUT35), .B2(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n616_), .B1(new_n519_), .B2(new_n613_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(KEYINPUT35), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G190gat), .B(G218gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G134gat), .B(G162gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT36), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT74), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n619_), .A2(new_n624_), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n617_), .A2(new_n618_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n622_), .A2(KEYINPUT36), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n617_), .A2(new_n618_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n626_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n625_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT73), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n625_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n630_), .A2(new_n632_), .A3(KEYINPUT37), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT37), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n625_), .B(new_n629_), .C1(new_n631_), .C2(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n581_), .B1(new_n633_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n613_), .A2(KEYINPUT12), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n639_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n613_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n574_), .A2(new_n564_), .A3(new_n612_), .A4(new_n611_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT12), .ZN(new_n643_));
  AOI22_X1  g442(.A1(new_n640_), .A2(KEYINPUT71), .B1(new_n641_), .B2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(G230gat), .A2(G233gat), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT70), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n646_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n574_), .A2(KEYINPUT70), .A3(new_n564_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n638_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT71), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n644_), .A2(new_n645_), .A3(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n645_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT69), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(G120gat), .B(G148gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT5), .ZN(new_n657_));
  XNOR2_X1  g456(.A(G176gat), .B(G204gat), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n657_), .B(new_n658_), .Z(new_n659_));
  NAND2_X1  g458(.A1(new_n655_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n659_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n652_), .A2(new_n654_), .A3(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT13), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n660_), .A2(KEYINPUT13), .A3(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n637_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n534_), .A2(new_n668_), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n669_), .A2(G1gat), .A3(new_n457_), .ZN(new_n670_));
  XOR2_X1   g469(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n671_));
  OR2_X1    g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n458_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n470_), .A2(new_n472_), .A3(new_n489_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n460_), .A2(new_n461_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n673_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(new_n630_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n667_), .A2(new_n533_), .A3(new_n581_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G1gat), .B1(new_n680_), .B2(new_n457_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n670_), .A2(new_n671_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n672_), .A2(new_n681_), .A3(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT102), .ZN(G1324gat));
  NAND3_X1  g483(.A1(new_n678_), .A2(new_n325_), .A3(new_n679_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT39), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n685_), .A2(new_n686_), .A3(G8gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n685_), .B2(G8gat), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n325_), .A2(new_n493_), .ZN(new_n689_));
  OAI22_X1  g488(.A1(new_n687_), .A2(new_n688_), .B1(new_n669_), .B2(new_n689_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g490(.A1(new_n678_), .A2(new_n675_), .A3(new_n679_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n692_), .A2(new_n693_), .A3(G15gat), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT41), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n693_), .B1(new_n692_), .B2(G15gat), .ZN(new_n697_));
  OR3_X1    g496(.A1(new_n695_), .A2(new_n696_), .A3(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n696_), .B1(new_n695_), .B2(new_n697_), .ZN(new_n699_));
  OR3_X1    g498(.A1(new_n669_), .A2(G15gat), .A3(new_n462_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n698_), .A2(new_n699_), .A3(new_n700_), .ZN(G1326gat));
  OAI21_X1  g500(.A(G22gat), .B1(new_n680_), .B2(new_n488_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT42), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n488_), .A2(G22gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n703_), .B1(new_n669_), .B2(new_n704_), .ZN(G1327gat));
  INV_X1    g504(.A(new_n630_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n581_), .A2(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n667_), .A2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n534_), .A2(new_n708_), .ZN(new_n709_));
  OR3_X1    g508(.A1(new_n709_), .A2(G29gat), .A3(new_n457_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n581_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n667_), .A2(new_n533_), .A3(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(KEYINPUT104), .A2(KEYINPUT43), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(KEYINPUT104), .A2(KEYINPUT43), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n633_), .A2(new_n635_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n716_), .B1(new_n676_), .B2(new_n718_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n491_), .A2(new_n717_), .A3(new_n714_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n712_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT105), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n723_));
  INV_X1    g522(.A(new_n712_), .ZN(new_n724_));
  OAI22_X1  g523(.A1(new_n491_), .A2(new_n717_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n385_), .A2(new_n457_), .A3(new_n310_), .A4(new_n324_), .ZN(new_n726_));
  AOI22_X1  g525(.A1(KEYINPUT100), .A2(new_n726_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n675_), .B1(new_n470_), .B2(new_n727_), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n718_), .B(new_n713_), .C1(new_n728_), .C2(new_n458_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n724_), .B1(new_n725_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n722_), .A2(new_n723_), .A3(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n457_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n730_), .A2(KEYINPUT44), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n733_), .A2(new_n734_), .A3(new_n735_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n736_), .A2(KEYINPUT106), .A3(G29gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT106), .B1(new_n736_), .B2(G29gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n710_), .B1(new_n737_), .B2(new_n738_), .ZN(G1328gat));
  INV_X1    g538(.A(KEYINPUT107), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT46), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n743_));
  INV_X1    g542(.A(G36gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n468_), .B1(new_n730_), .B2(KEYINPUT44), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n733_), .B2(new_n745_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n709_), .A2(G36gat), .A3(new_n468_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT45), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n742_), .B(new_n743_), .C1(new_n746_), .C2(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n723_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n750_));
  AOI211_X1 g549(.A(KEYINPUT105), .B(new_n724_), .C1(new_n725_), .C2(new_n729_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n745_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(G36gat), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT45), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n747_), .B(new_n754_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n753_), .A2(new_n740_), .A3(new_n741_), .A4(new_n755_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n749_), .A2(new_n756_), .ZN(G1329gat));
  OAI21_X1  g556(.A(new_n389_), .B1(new_n709_), .B2(new_n462_), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT108), .Z(new_n759_));
  NAND2_X1  g558(.A1(new_n733_), .A2(new_n735_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n430_), .A2(G43gat), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n759_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT47), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT47), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n759_), .B(new_n764_), .C1(new_n760_), .C2(new_n761_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(G1330gat));
  OAI211_X1 g565(.A(new_n385_), .B(new_n735_), .C1(new_n750_), .C2(new_n751_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(G50gat), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n488_), .A2(G50gat), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT109), .Z(new_n770_));
  NAND3_X1  g569(.A1(new_n534_), .A2(new_n708_), .A3(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n768_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n768_), .A2(KEYINPUT110), .A3(new_n771_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1331gat));
  NAND2_X1  g575(.A1(new_n528_), .A2(new_n532_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n491_), .A2(new_n777_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n778_), .A2(KEYINPUT112), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n778_), .A2(KEYINPUT112), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n667_), .A2(new_n636_), .A3(KEYINPUT111), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT111), .B1(new_n667_), .B2(new_n636_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(KEYINPUT113), .B1(new_n781_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n781_), .A2(new_n784_), .A3(KEYINPUT113), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n457_), .A2(G57gat), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n786_), .A2(new_n787_), .A3(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n667_), .A2(new_n533_), .A3(new_n711_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n677_), .A2(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n547_), .B1(new_n792_), .B2(new_n734_), .ZN(new_n793_));
  OAI21_X1  g592(.A(KEYINPUT114), .B1(new_n790_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n787_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n795_), .A2(new_n785_), .A3(new_n788_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT114), .ZN(new_n797_));
  INV_X1    g596(.A(new_n793_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n796_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n794_), .A2(new_n799_), .ZN(G1332gat));
  NOR2_X1   g599(.A1(new_n468_), .A2(G64gat), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n786_), .A2(new_n787_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT48), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n792_), .A2(new_n325_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(G64gat), .ZN(new_n806_));
  AOI211_X1 g605(.A(KEYINPUT48), .B(new_n545_), .C1(new_n792_), .C2(new_n325_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT115), .B1(new_n803_), .B2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n795_), .A2(new_n785_), .A3(new_n801_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n811_));
  INV_X1    g610(.A(new_n808_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n810_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n809_), .A2(new_n813_), .ZN(G1333gat));
  NOR2_X1   g613(.A1(new_n786_), .A2(new_n787_), .ZN(new_n815_));
  INV_X1    g614(.A(G71gat), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n816_), .A3(new_n675_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n816_), .B1(new_n792_), .B2(new_n675_), .ZN(new_n818_));
  XOR2_X1   g617(.A(new_n818_), .B(KEYINPUT49), .Z(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(G1334gat));
  INV_X1    g619(.A(G78gat), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n815_), .A2(new_n821_), .A3(new_n385_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n821_), .B1(new_n792_), .B2(new_n385_), .ZN(new_n823_));
  XOR2_X1   g622(.A(new_n823_), .B(KEYINPUT50), .Z(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(G1335gat));
  INV_X1    g624(.A(new_n667_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n781_), .A2(new_n826_), .A3(new_n707_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n827_), .A2(new_n592_), .A3(new_n734_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n667_), .A2(new_n533_), .A3(new_n581_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n829_), .B1(new_n725_), .B2(new_n729_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(G85gat), .B1(new_n831_), .B2(new_n457_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n828_), .A2(new_n832_), .ZN(G1336gat));
  NAND3_X1  g632(.A1(new_n827_), .A2(new_n593_), .A3(new_n325_), .ZN(new_n834_));
  OAI21_X1  g633(.A(G92gat), .B1(new_n831_), .B2(new_n468_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(G1337gat));
  NAND2_X1  g635(.A1(KEYINPUT117), .A2(KEYINPUT51), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n826_), .A2(new_n707_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n430_), .A2(new_n603_), .A3(new_n607_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n837_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n585_), .B1(new_n830_), .B2(new_n675_), .ZN(new_n842_));
  OR2_X1    g641(.A1(new_n842_), .A2(KEYINPUT116), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(KEYINPUT116), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n841_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(KEYINPUT117), .A2(KEYINPUT51), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n845_), .B(new_n846_), .ZN(G1338gat));
  AND2_X1   g646(.A1(new_n604_), .A2(new_n606_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n827_), .A2(new_n385_), .A3(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT52), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n830_), .A2(new_n385_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(G106gat), .ZN(new_n852_));
  AOI211_X1 g651(.A(KEYINPUT52), .B(new_n586_), .C1(new_n830_), .C2(new_n385_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n849_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(KEYINPUT53), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n849_), .B(new_n856_), .C1(new_n852_), .C2(new_n853_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(G1339gat));
  NAND4_X1  g657(.A1(new_n636_), .A2(new_n666_), .A3(new_n665_), .A4(new_n533_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(KEYINPUT118), .A2(KEYINPUT54), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n859_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n514_), .B1(new_n519_), .B2(new_n502_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n524_), .B1(new_n512_), .B2(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n866_), .B1(new_n527_), .B2(new_n515_), .ZN(new_n867_));
  AND3_X1   g666(.A1(new_n663_), .A2(new_n528_), .A3(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n643_), .A2(new_n641_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n645_), .ZN(new_n871_));
  AOI211_X1 g670(.A(KEYINPUT71), .B(new_n638_), .C1(new_n647_), .C2(new_n648_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n870_), .A2(new_n871_), .A3(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n871_), .B1(new_n870_), .B2(new_n872_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n873_), .B1(KEYINPUT55), .B2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT55), .ZN(new_n876_));
  NOR4_X1   g675(.A1(new_n870_), .A2(new_n872_), .A3(new_n876_), .A4(new_n871_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n659_), .B1(new_n875_), .B2(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n662_), .A2(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n533_), .B1(new_n878_), .B2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n879_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n645_), .B1(new_n644_), .B2(new_n651_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n652_), .B1(new_n883_), .B2(new_n876_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n877_), .ZN(new_n885_));
  AOI211_X1 g684(.A(new_n661_), .B(new_n882_), .C1(new_n884_), .C2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n868_), .B1(new_n881_), .B2(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n864_), .B1(new_n888_), .B2(new_n706_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(KEYINPUT58), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n528_), .A2(new_n662_), .A3(new_n867_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n892_), .B1(new_n878_), .B2(KEYINPUT56), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n661_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT56), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n891_), .B1(new_n893_), .B2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n878_), .A2(KEYINPUT56), .ZN(new_n898_));
  INV_X1    g697(.A(new_n891_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n894_), .A2(new_n895_), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n898_), .A2(new_n899_), .A3(new_n900_), .A4(new_n892_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n897_), .A2(new_n901_), .A3(new_n718_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n663_), .A2(new_n528_), .A3(new_n867_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n662_), .A2(new_n879_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n777_), .B1(new_n894_), .B2(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n903_), .B1(new_n905_), .B2(new_n886_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n906_), .A2(KEYINPUT57), .A3(new_n630_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n889_), .A2(new_n902_), .A3(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n863_), .B1(new_n908_), .B2(new_n581_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n386_), .A2(new_n430_), .A3(new_n734_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(G113gat), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n911_), .A2(new_n912_), .A3(new_n777_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n910_), .ZN(new_n914_));
  AND3_X1   g713(.A1(new_n906_), .A2(KEYINPUT57), .A3(new_n630_), .ZN(new_n915_));
  AOI21_X1  g714(.A(KEYINPUT57), .B1(new_n906_), .B2(new_n630_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n711_), .B1(new_n917_), .B2(new_n902_), .ZN(new_n918_));
  OAI211_X1 g717(.A(KEYINPUT59), .B(new_n914_), .C1(new_n918_), .C2(new_n863_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT59), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n920_), .B1(new_n909_), .B2(new_n910_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n533_), .B1(new_n919_), .B2(new_n921_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n913_), .B1(new_n922_), .B2(new_n912_), .ZN(G1340gat));
  INV_X1    g722(.A(G120gat), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n924_), .B1(new_n826_), .B2(KEYINPUT60), .ZN(new_n925_));
  OAI211_X1 g724(.A(new_n911_), .B(new_n925_), .C1(KEYINPUT60), .C2(new_n924_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n826_), .B1(new_n919_), .B2(new_n921_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n927_), .B2(new_n924_), .ZN(G1341gat));
  AOI21_X1  g727(.A(G127gat), .B1(new_n911_), .B2(new_n711_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n919_), .A2(new_n921_), .ZN(new_n930_));
  XOR2_X1   g729(.A(KEYINPUT121), .B(G127gat), .Z(new_n931_));
  NAND2_X1  g730(.A1(new_n711_), .A2(new_n931_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(KEYINPUT122), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n929_), .B1(new_n930_), .B2(new_n933_), .ZN(G1342gat));
  NOR2_X1   g733(.A1(new_n717_), .A2(new_n405_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n908_), .A2(new_n581_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n863_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(KEYINPUT59), .B1(new_n938_), .B2(new_n914_), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n909_), .A2(new_n920_), .A3(new_n910_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n935_), .B1(new_n939_), .B2(new_n940_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n911_), .A2(new_n706_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n942_), .A2(new_n405_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n941_), .A2(KEYINPUT123), .A3(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT123), .ZN(new_n945_));
  INV_X1    g744(.A(new_n935_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n946_), .B1(new_n919_), .B2(new_n921_), .ZN(new_n947_));
  AOI21_X1  g746(.A(G134gat), .B1(new_n911_), .B2(new_n706_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n945_), .B1(new_n947_), .B2(new_n948_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n944_), .A2(new_n949_), .ZN(G1343gat));
  NOR3_X1   g749(.A1(new_n325_), .A2(new_n488_), .A3(new_n457_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n462_), .A2(new_n951_), .ZN(new_n952_));
  INV_X1    g751(.A(new_n952_), .ZN(new_n953_));
  AOI21_X1  g752(.A(KEYINPUT124), .B1(new_n938_), .B2(new_n953_), .ZN(new_n954_));
  INV_X1    g753(.A(KEYINPUT124), .ZN(new_n955_));
  NOR3_X1   g754(.A1(new_n909_), .A2(new_n955_), .A3(new_n952_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n777_), .B1(new_n954_), .B2(new_n956_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n957_), .A2(G141gat), .ZN(new_n958_));
  OAI211_X1 g757(.A(new_n328_), .B(new_n777_), .C1(new_n954_), .C2(new_n956_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n958_), .A2(new_n959_), .ZN(G1344gat));
  OAI21_X1  g759(.A(new_n667_), .B1(new_n954_), .B2(new_n956_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(KEYINPUT125), .B(G148gat), .ZN(new_n962_));
  INV_X1    g761(.A(new_n962_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n961_), .A2(new_n963_), .ZN(new_n964_));
  OAI211_X1 g763(.A(new_n667_), .B(new_n962_), .C1(new_n954_), .C2(new_n956_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n964_), .A2(new_n965_), .ZN(G1345gat));
  OAI21_X1  g765(.A(new_n711_), .B1(new_n954_), .B2(new_n956_), .ZN(new_n967_));
  XNOR2_X1  g766(.A(KEYINPUT61), .B(G155gat), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n967_), .A2(new_n968_), .ZN(new_n969_));
  INV_X1    g768(.A(new_n968_), .ZN(new_n970_));
  OAI211_X1 g769(.A(new_n711_), .B(new_n970_), .C1(new_n954_), .C2(new_n956_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n969_), .A2(new_n971_), .ZN(G1346gat));
  OR2_X1    g771(.A1(new_n954_), .A2(new_n956_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n718_), .A2(G162gat), .ZN(new_n974_));
  XNOR2_X1  g773(.A(new_n974_), .B(KEYINPUT126), .ZN(new_n975_));
  OAI21_X1  g774(.A(new_n706_), .B1(new_n954_), .B2(new_n956_), .ZN(new_n976_));
  AOI22_X1  g775(.A1(new_n973_), .A2(new_n975_), .B1(new_n976_), .B2(new_n340_), .ZN(G1347gat));
  INV_X1    g776(.A(KEYINPUT62), .ZN(new_n978_));
  NOR2_X1   g777(.A1(new_n909_), .A2(new_n468_), .ZN(new_n979_));
  NOR3_X1   g778(.A1(new_n462_), .A2(new_n734_), .A3(new_n385_), .ZN(new_n980_));
  AND3_X1   g779(.A1(new_n979_), .A2(new_n777_), .A3(new_n980_), .ZN(new_n981_));
  OAI21_X1  g780(.A(new_n978_), .B1(new_n981_), .B2(new_n212_), .ZN(new_n982_));
  NAND3_X1  g781(.A1(new_n981_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n983_));
  NAND2_X1  g782(.A1(new_n979_), .A2(new_n980_), .ZN(new_n984_));
  OAI211_X1 g783(.A(KEYINPUT62), .B(G169gat), .C1(new_n984_), .C2(new_n533_), .ZN(new_n985_));
  NAND3_X1  g784(.A1(new_n982_), .A2(new_n983_), .A3(new_n985_), .ZN(G1348gat));
  NAND3_X1  g785(.A1(new_n979_), .A2(new_n667_), .A3(new_n980_), .ZN(new_n987_));
  NOR2_X1   g786(.A1(new_n987_), .A2(new_n208_), .ZN(new_n988_));
  AOI21_X1  g787(.A(new_n988_), .B1(new_n219_), .B2(new_n987_), .ZN(G1349gat));
  NAND3_X1  g788(.A1(new_n979_), .A2(new_n711_), .A3(new_n980_), .ZN(new_n990_));
  AND2_X1   g789(.A1(new_n265_), .A2(new_n267_), .ZN(new_n991_));
  NOR2_X1   g790(.A1(new_n990_), .A2(new_n991_), .ZN(new_n992_));
  AOI21_X1  g791(.A(new_n992_), .B1(new_n229_), .B2(new_n990_), .ZN(G1350gat));
  OAI21_X1  g792(.A(G190gat), .B1(new_n984_), .B2(new_n717_), .ZN(new_n994_));
  NAND3_X1  g793(.A1(new_n706_), .A2(new_n268_), .A3(new_n270_), .ZN(new_n995_));
  OAI21_X1  g794(.A(new_n994_), .B1(new_n984_), .B2(new_n995_), .ZN(G1351gat));
  NOR2_X1   g795(.A1(new_n675_), .A2(new_n471_), .ZN(new_n997_));
  NAND2_X1  g796(.A1(new_n979_), .A2(new_n997_), .ZN(new_n998_));
  OAI21_X1  g797(.A(new_n251_), .B1(new_n998_), .B2(new_n533_), .ZN(new_n999_));
  NAND4_X1  g798(.A1(new_n979_), .A2(G197gat), .A3(new_n777_), .A4(new_n997_), .ZN(new_n1000_));
  NAND2_X1  g799(.A1(new_n1000_), .A2(KEYINPUT127), .ZN(new_n1001_));
  NOR4_X1   g800(.A1(new_n909_), .A2(new_n675_), .A3(new_n471_), .A4(new_n468_), .ZN(new_n1002_));
  INV_X1    g801(.A(KEYINPUT127), .ZN(new_n1003_));
  NAND4_X1  g802(.A1(new_n1002_), .A2(new_n1003_), .A3(G197gat), .A4(new_n777_), .ZN(new_n1004_));
  AND3_X1   g803(.A1(new_n999_), .A2(new_n1001_), .A3(new_n1004_), .ZN(G1352gat));
  AOI21_X1  g804(.A(G204gat), .B1(new_n1002_), .B2(new_n667_), .ZN(new_n1006_));
  NAND2_X1  g805(.A1(new_n246_), .A2(new_n247_), .ZN(new_n1007_));
  NOR2_X1   g806(.A1(new_n998_), .A2(new_n826_), .ZN(new_n1008_));
  AOI21_X1  g807(.A(new_n1006_), .B1(new_n1007_), .B2(new_n1008_), .ZN(G1353gat));
  NAND3_X1  g808(.A1(new_n979_), .A2(new_n711_), .A3(new_n997_), .ZN(new_n1010_));
  XNOR2_X1  g809(.A(KEYINPUT63), .B(G211gat), .ZN(new_n1011_));
  NOR2_X1   g810(.A1(new_n1010_), .A2(new_n1011_), .ZN(new_n1012_));
  NOR2_X1   g811(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1013_));
  AOI21_X1  g812(.A(new_n1012_), .B1(new_n1010_), .B2(new_n1013_), .ZN(G1354gat));
  OAI21_X1  g813(.A(G218gat), .B1(new_n998_), .B2(new_n717_), .ZN(new_n1015_));
  NAND3_X1  g814(.A1(new_n1002_), .A2(new_n239_), .A3(new_n706_), .ZN(new_n1016_));
  NAND2_X1  g815(.A1(new_n1015_), .A2(new_n1016_), .ZN(G1355gat));
endmodule


