//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n626_, new_n627_, new_n628_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n634_, new_n635_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n831_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n837_, new_n839_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n877_, new_n878_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(KEYINPUT88), .Z(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT31), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G71gat), .B(G99gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT84), .B(KEYINPUT23), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT23), .ZN(new_n210_));
  INV_X1    g009(.A(G183gat), .ZN(new_n211_));
  INV_X1    g010(.A(G190gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  MUX2_X1   g012(.A(new_n209_), .B(new_n210_), .S(new_n213_), .Z(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT25), .B(G183gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT26), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT83), .B1(new_n216_), .B2(G190gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT26), .B(G190gat), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n215_), .B(new_n217_), .C1(new_n218_), .C2(KEYINPUT83), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT24), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222_));
  MUX2_X1   g021(.A(new_n221_), .B(KEYINPUT24), .S(new_n222_), .Z(new_n223_));
  NAND3_X1  g022(.A1(new_n214_), .A2(new_n219_), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n209_), .A2(new_n213_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n211_), .A2(new_n212_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n210_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  XOR2_X1   g027(.A(KEYINPUT86), .B(G176gat), .Z(new_n229_));
  INV_X1    g028(.A(KEYINPUT85), .ZN(new_n230_));
  INV_X1    g029(.A(G169gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n230_), .B1(new_n231_), .B2(KEYINPUT22), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT22), .B(G169gat), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n229_), .B(new_n232_), .C1(new_n230_), .C2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n228_), .A2(new_n234_), .A3(new_n220_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n224_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G227gat), .A2(G233gat), .ZN(new_n237_));
  INV_X1    g036(.A(G15gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT30), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n236_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT87), .B(G43gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n208_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n208_), .A2(new_n243_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G141gat), .A2(G148gat), .ZN(new_n248_));
  OR2_X1    g047(.A1(G141gat), .A2(G148gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G155gat), .A2(G162gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT1), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n251_), .B(KEYINPUT90), .Z(new_n252_));
  OR3_X1    g051(.A1(KEYINPUT89), .A2(G155gat), .A3(G162gat), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT89), .B1(G155gat), .B2(G162gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n255_), .B1(KEYINPUT1), .B2(new_n250_), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n248_), .B(new_n249_), .C1(new_n252_), .C2(new_n256_), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n255_), .A2(new_n250_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT92), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT2), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n249_), .A2(KEYINPUT3), .B1(new_n260_), .B2(new_n248_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n261_), .B1(KEYINPUT3), .B2(new_n249_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n263_));
  XOR2_X1   g062(.A(new_n263_), .B(KEYINPUT91), .Z(new_n264_));
  OAI22_X1  g063(.A1(new_n258_), .A2(new_n259_), .B1(new_n262_), .B2(new_n264_), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n258_), .A2(new_n259_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n257_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n205_), .A2(new_n267_), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n204_), .B(new_n257_), .C1(new_n265_), .C2(new_n266_), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT4), .ZN(new_n271_));
  AND2_X1   g070(.A1(G225gat), .A2(G233gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT104), .B(KEYINPUT4), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n205_), .A2(new_n267_), .A3(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n271_), .A2(new_n272_), .A3(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n268_), .A2(new_n269_), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT105), .B1(new_n276_), .B2(new_n272_), .ZN(new_n277_));
  OR3_X1    g076(.A1(new_n276_), .A2(KEYINPUT105), .A3(new_n272_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n275_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G1gat), .B(G29gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(G85gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT0), .B(G57gat), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n281_), .B(new_n282_), .Z(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n279_), .A2(new_n284_), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n275_), .A2(new_n283_), .A3(new_n277_), .A4(new_n278_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(G204gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n288_), .A2(KEYINPUT95), .A3(G197gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G197gat), .B(G204gat), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  OAI211_X1 g090(.A(KEYINPUT21), .B(new_n289_), .C1(new_n291_), .C2(KEYINPUT95), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT96), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT21), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n290_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT97), .ZN(new_n297_));
  XOR2_X1   g096(.A(G211gat), .B(G218gat), .Z(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n294_), .A2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n291_), .A2(KEYINPUT21), .A3(new_n298_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(new_n236_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT101), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n302_), .A2(KEYINPUT101), .A3(new_n236_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G226gat), .A2(G233gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT19), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT20), .ZN(new_n311_));
  INV_X1    g110(.A(new_n302_), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n220_), .B(KEYINPUT99), .Z(new_n313_));
  AOI21_X1  g112(.A(new_n313_), .B1(new_n214_), .B2(new_n226_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n233_), .B(KEYINPUT100), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n229_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n225_), .A2(new_n227_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n317_), .B1(new_n218_), .B2(new_n215_), .ZN(new_n318_));
  AOI22_X1  g117(.A1(new_n314_), .A2(new_n316_), .B1(new_n318_), .B2(new_n223_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n311_), .B1(new_n312_), .B2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n307_), .A2(new_n310_), .A3(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT20), .B1(new_n312_), .B2(new_n319_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n302_), .A2(new_n236_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n309_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(G64gat), .B(G92gat), .Z(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT103), .ZN(new_n326_));
  XOR2_X1   g125(.A(KEYINPUT102), .B(KEYINPUT18), .Z(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G8gat), .B(G36gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT32), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n321_), .A2(new_n324_), .A3(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n310_), .B1(new_n307_), .B2(new_n320_), .ZN(new_n333_));
  NOR3_X1   g132(.A1(new_n322_), .A2(new_n309_), .A3(new_n323_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n287_), .B(new_n332_), .C1(new_n331_), .C2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT33), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n286_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT106), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n321_), .A2(new_n330_), .A3(new_n324_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n330_), .B1(new_n321_), .B2(new_n324_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n286_), .A2(new_n337_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n283_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n271_), .A2(new_n274_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n344_), .B1(new_n345_), .B2(new_n272_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n342_), .A2(new_n343_), .A3(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n336_), .B1(new_n339_), .B2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n267_), .A2(KEYINPUT29), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT28), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G22gat), .B(G50gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT94), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n267_), .A2(KEYINPUT29), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n302_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G78gat), .B(G106gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT98), .ZN(new_n357_));
  INV_X1    g156(.A(G228gat), .ZN(new_n358_));
  INV_X1    g157(.A(G233gat), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n359_), .A2(KEYINPUT93), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(KEYINPUT93), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n358_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n357_), .B(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n355_), .B(new_n363_), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n352_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n352_), .A2(new_n364_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n348_), .A2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n287_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT27), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n370_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n330_), .B(KEYINPUT107), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n372_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n321_), .A2(new_n330_), .A3(new_n324_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(KEYINPUT27), .A3(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n369_), .A2(new_n371_), .A3(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n247_), .B1(new_n368_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT109), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT108), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n371_), .A2(new_n379_), .A3(new_n375_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n379_), .B1(new_n371_), .B2(new_n375_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n367_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n378_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  OAI211_X1 g183(.A(KEYINPUT109), .B(new_n367_), .C1(new_n380_), .C2(new_n381_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n287_), .A2(new_n246_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n377_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G29gat), .B(G36gat), .ZN(new_n389_));
  OR2_X1    g188(.A1(new_n389_), .A2(KEYINPUT74), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(KEYINPUT74), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G43gat), .B(G50gat), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n390_), .A2(new_n391_), .A3(new_n393_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT15), .ZN(new_n398_));
  XOR2_X1   g197(.A(G15gat), .B(G22gat), .Z(new_n399_));
  NAND2_X1  g198(.A1(G1gat), .A2(G8gat), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n399_), .B1(KEYINPUT14), .B2(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT79), .ZN(new_n402_));
  XOR2_X1   g201(.A(G1gat), .B(G8gat), .Z(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT79), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n401_), .B(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n403_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n404_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n398_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n404_), .A2(new_n408_), .A3(new_n397_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G229gat), .A2(G233gat), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n410_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n409_), .B(new_n397_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n413_), .B1(new_n414_), .B2(new_n412_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G113gat), .B(G141gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G169gat), .B(G197gat), .ZN(new_n417_));
  XOR2_X1   g216(.A(new_n416_), .B(new_n417_), .Z(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n415_), .A2(new_n419_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n413_), .B(new_n418_), .C1(new_n414_), .C2(new_n412_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n388_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G230gat), .A2(G233gat), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT65), .ZN(new_n426_));
  AND2_X1   g225(.A1(G85gat), .A2(G92gat), .ZN(new_n427_));
  NOR2_X1   g226(.A1(G85gat), .A2(G92gat), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT9), .ZN(new_n429_));
  NOR3_X1   g228(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n429_), .A2(G85gat), .A3(G92gat), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n426_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n428_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G85gat), .A2(G92gat), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n434_), .A2(KEYINPUT9), .A3(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(KEYINPUT65), .A3(new_n431_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n433_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT66), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT6), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n440_), .B1(G99gat), .B2(G106gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G99gat), .A2(G106gat), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n442_), .A2(KEYINPUT6), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n439_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n444_));
  OR2_X1    g243(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n445_));
  OR2_X1    g244(.A1(KEYINPUT64), .A2(G106gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(KEYINPUT64), .A2(G106gat), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .A4(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n442_), .A2(KEYINPUT6), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n440_), .A2(G99gat), .A3(G106gat), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n450_), .A2(new_n451_), .A3(KEYINPUT66), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n444_), .A2(new_n449_), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT67), .ZN(new_n454_));
  AND3_X1   g253(.A1(new_n438_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n454_), .B1(new_n438_), .B2(new_n453_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT8), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT7), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT68), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n459_), .A2(G99gat), .ZN(new_n460_));
  INV_X1    g259(.A(G106gat), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n458_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(G99gat), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n458_), .A2(new_n463_), .A3(new_n461_), .A4(KEYINPUT68), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT69), .B1(new_n462_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n450_), .A2(new_n451_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n463_), .A2(new_n461_), .A3(KEYINPUT68), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT7), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT69), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n469_), .A2(new_n470_), .A3(new_n464_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n466_), .A2(new_n467_), .A3(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n427_), .A2(new_n428_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n457_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n457_), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n450_), .A2(new_n451_), .A3(KEYINPUT66), .ZN(new_n476_));
  AOI21_X1  g275(.A(KEYINPUT66), .B1(new_n450_), .B2(new_n451_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n469_), .A2(new_n464_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n475_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n481_));
  OAI22_X1  g280(.A1(new_n455_), .A2(new_n456_), .B1(new_n474_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT70), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G57gat), .B(G64gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G71gat), .B(G78gat), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n484_), .A2(new_n485_), .A3(KEYINPUT11), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(KEYINPUT11), .ZN(new_n487_));
  INV_X1    g286(.A(new_n485_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n484_), .A2(KEYINPUT11), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n483_), .B(new_n486_), .C1(new_n489_), .C2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  OR2_X1    g291(.A1(new_n484_), .A2(KEYINPUT11), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n493_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n483_), .B1(new_n494_), .B2(new_n486_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n492_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n482_), .A2(new_n497_), .ZN(new_n498_));
  NOR3_X1   g297(.A1(new_n430_), .A2(new_n426_), .A3(new_n432_), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT65), .B1(new_n436_), .B2(new_n431_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n478_), .A2(new_n449_), .ZN(new_n502_));
  OAI21_X1  g301(.A(KEYINPUT67), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n438_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n481_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n473_), .ZN(new_n507_));
  AOI22_X1  g306(.A1(new_n479_), .A2(KEYINPUT69), .B1(new_n450_), .B2(new_n451_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n507_), .B1(new_n508_), .B2(new_n471_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n506_), .B1(new_n509_), .B2(new_n457_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n505_), .A2(new_n510_), .A3(new_n496_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n425_), .B1(new_n498_), .B2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n494_), .A2(KEYINPUT12), .A3(new_n486_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n455_), .A2(new_n456_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n472_), .A2(new_n473_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n481_), .B1(new_n516_), .B2(KEYINPUT8), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n514_), .B1(new_n515_), .B2(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n496_), .B1(new_n505_), .B2(new_n510_), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n518_), .B(new_n511_), .C1(new_n519_), .C2(KEYINPUT12), .ZN(new_n520_));
  INV_X1    g319(.A(new_n425_), .ZN(new_n521_));
  OAI21_X1  g320(.A(KEYINPUT71), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  AND3_X1   g321(.A1(new_n505_), .A2(new_n510_), .A3(new_n496_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n513_), .B1(new_n505_), .B2(new_n510_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT12), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n498_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT71), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n525_), .A2(new_n527_), .A3(new_n528_), .A4(new_n425_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n512_), .B1(new_n522_), .B2(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n530_), .A2(KEYINPUT72), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G120gat), .B(G148gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT5), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G176gat), .B(G204gat), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n533_), .B(new_n534_), .Z(new_n535_));
  OAI21_X1  g334(.A(new_n535_), .B1(new_n530_), .B2(KEYINPUT72), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT73), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n522_), .A2(new_n529_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n512_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n535_), .ZN(new_n540_));
  AND4_X1   g339(.A1(new_n537_), .A2(new_n538_), .A3(new_n539_), .A4(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n537_), .B1(new_n530_), .B2(new_n540_), .ZN(new_n542_));
  OAI22_X1  g341(.A1(new_n531_), .A2(new_n536_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n544_), .A2(KEYINPUT13), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(KEYINPUT13), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n398_), .A2(new_n482_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n516_), .A2(KEYINPUT8), .ZN(new_n550_));
  AOI22_X1  g349(.A1(new_n550_), .A2(new_n506_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n397_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G232gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT34), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n554_), .A2(KEYINPUT35), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n549_), .A2(new_n552_), .A3(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n556_), .A2(KEYINPUT35), .A3(new_n554_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n554_), .A2(KEYINPUT35), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n549_), .A2(new_n552_), .A3(new_n558_), .A4(new_n555_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G190gat), .B(G218gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G134gat), .B(G162gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n563_), .B(KEYINPUT36), .Z(new_n564_));
  XOR2_X1   g363(.A(new_n564_), .B(KEYINPUT76), .Z(new_n565_));
  NAND2_X1  g364(.A1(new_n560_), .A2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT75), .B(KEYINPUT36), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n563_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n557_), .A2(new_n559_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n566_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(KEYINPUT37), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT77), .ZN(new_n572_));
  INV_X1    g371(.A(new_n569_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n564_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT78), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n574_), .B1(new_n560_), .B2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n557_), .A2(KEYINPUT78), .A3(new_n559_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n573_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT37), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT77), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n570_), .A2(new_n581_), .A3(KEYINPUT37), .ZN(new_n582_));
  AND3_X1   g381(.A1(new_n572_), .A2(new_n580_), .A3(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(KEYINPUT82), .B(KEYINPUT17), .Z(new_n584_));
  XOR2_X1   g383(.A(G127gat), .B(G155gat), .Z(new_n585_));
  XNOR2_X1  g384(.A(G183gat), .B(G211gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n587_), .B(new_n588_), .Z(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(G231gat), .A2(G233gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n409_), .B(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n494_), .A2(new_n486_), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n593_), .B(KEYINPUT80), .Z(new_n594_));
  AOI211_X1 g393(.A(new_n584_), .B(new_n590_), .C1(new_n592_), .C2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n595_), .B1(new_n592_), .B2(new_n594_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n589_), .B(KEYINPUT17), .ZN(new_n597_));
  INV_X1    g396(.A(new_n592_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n597_), .B1(new_n598_), .B2(new_n497_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n599_), .B1(new_n497_), .B2(new_n598_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n596_), .A2(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n583_), .A2(new_n601_), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n424_), .A2(new_n548_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(G1gat), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n603_), .A2(new_n604_), .A3(new_n287_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT38), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n388_), .A2(new_n578_), .ZN(new_n608_));
  NOR3_X1   g407(.A1(new_n547_), .A2(new_n423_), .A3(new_n601_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n604_), .B1(new_n610_), .B2(new_n287_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n607_), .A2(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n612_), .B1(new_n606_), .B2(new_n605_), .ZN(G1324gat));
  INV_X1    g412(.A(G8gat), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n603_), .A2(new_n614_), .A3(new_n382_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT39), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n610_), .A2(new_n382_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n616_), .B1(new_n617_), .B2(G8gat), .ZN(new_n618_));
  AOI211_X1 g417(.A(KEYINPUT39), .B(new_n614_), .C1(new_n610_), .C2(new_n382_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n615_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(KEYINPUT110), .B(KEYINPUT40), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n615_), .B(new_n621_), .C1(new_n618_), .C2(new_n619_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1325gat));
  AOI21_X1  g424(.A(new_n238_), .B1(new_n610_), .B2(new_n247_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT41), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n603_), .A2(new_n238_), .A3(new_n247_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(G1326gat));
  INV_X1    g428(.A(G22gat), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n603_), .A2(new_n630_), .A3(new_n383_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n630_), .B1(new_n610_), .B2(new_n383_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(KEYINPUT111), .B(KEYINPUT42), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n632_), .A2(new_n633_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n631_), .B1(new_n634_), .B2(new_n635_), .ZN(G1327gat));
  INV_X1    g435(.A(new_n601_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n578_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n547_), .A2(new_n637_), .A3(new_n638_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n424_), .A2(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(G29gat), .B1(new_n640_), .B2(new_n287_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n583_), .ZN(new_n642_));
  OAI21_X1  g441(.A(KEYINPUT43), .B1(new_n388_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT43), .ZN(new_n644_));
  INV_X1    g443(.A(new_n387_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n645_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n646_));
  OAI211_X1 g445(.A(new_n644_), .B(new_n583_), .C1(new_n646_), .C2(new_n377_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n643_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n548_), .A2(new_n422_), .A3(new_n601_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(KEYINPUT44), .B1(new_n648_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT44), .ZN(new_n652_));
  AOI211_X1 g451(.A(new_n652_), .B(new_n649_), .C1(new_n643_), .C2(new_n647_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n287_), .A2(G29gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n641_), .B1(new_n654_), .B2(new_n655_), .ZN(G1328gat));
  INV_X1    g455(.A(KEYINPUT46), .ZN(new_n657_));
  INV_X1    g456(.A(G36gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n658_), .B1(new_n654_), .B2(new_n382_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n424_), .A2(new_n658_), .A3(new_n382_), .A4(new_n639_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n660_), .B(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n657_), .B1(new_n659_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n662_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n382_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n651_), .A2(new_n653_), .A3(new_n665_), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n664_), .B(KEYINPUT46), .C1(new_n666_), .C2(new_n658_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n663_), .A2(new_n667_), .ZN(G1329gat));
  NAND2_X1  g467(.A1(new_n648_), .A2(new_n650_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(new_n652_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n648_), .A2(KEYINPUT44), .A3(new_n650_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n247_), .A2(G43gat), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n670_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(G43gat), .B1(new_n640_), .B2(new_n247_), .ZN(new_n674_));
  OAI21_X1  g473(.A(KEYINPUT47), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n654_), .B2(new_n672_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT47), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n675_), .A2(new_n678_), .ZN(G1330gat));
  INV_X1    g478(.A(G50gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n640_), .A2(new_n680_), .A3(new_n383_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n670_), .A2(new_n383_), .A3(new_n671_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n682_), .A2(KEYINPUT113), .A3(G50gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT113), .B1(new_n682_), .B2(G50gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n681_), .B1(new_n683_), .B2(new_n684_), .ZN(G1331gat));
  NOR3_X1   g484(.A1(new_n388_), .A2(new_n422_), .A3(new_n548_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n686_), .A2(new_n602_), .ZN(new_n687_));
  INV_X1    g486(.A(G57gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(new_n688_), .A3(new_n287_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n548_), .A2(new_n422_), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n608_), .A2(new_n637_), .A3(new_n690_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n691_), .A2(new_n287_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n689_), .B1(new_n692_), .B2(new_n688_), .ZN(G1332gat));
  INV_X1    g492(.A(G64gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n694_), .B1(new_n691_), .B2(new_n382_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT48), .Z(new_n696_));
  NAND3_X1  g495(.A1(new_n687_), .A2(new_n694_), .A3(new_n382_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1333gat));
  INV_X1    g497(.A(G71gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n699_), .B1(new_n691_), .B2(new_n247_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT49), .Z(new_n701_));
  NAND3_X1  g500(.A1(new_n687_), .A2(new_n699_), .A3(new_n247_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1334gat));
  INV_X1    g502(.A(G78gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n704_), .B1(new_n691_), .B2(new_n383_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT50), .Z(new_n706_));
  NAND3_X1  g505(.A1(new_n687_), .A2(new_n704_), .A3(new_n383_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1335gat));
  NOR2_X1   g507(.A1(new_n638_), .A2(new_n637_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n686_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(G85gat), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n710_), .A2(new_n711_), .A3(new_n287_), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n648_), .A2(new_n601_), .A3(new_n690_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n713_), .A2(new_n287_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n712_), .B1(new_n714_), .B2(new_n711_), .ZN(G1336gat));
  AOI21_X1  g514(.A(G92gat), .B1(new_n710_), .B2(new_n382_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n382_), .A2(G92gat), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT114), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n716_), .B1(new_n713_), .B2(new_n718_), .ZN(G1337gat));
  NAND4_X1  g518(.A1(new_n648_), .A2(new_n247_), .A3(new_n601_), .A4(new_n690_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(G99gat), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n247_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n722_));
  AOI22_X1  g521(.A1(new_n710_), .A2(new_n722_), .B1(KEYINPUT115), .B2(KEYINPUT51), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n724_), .B(new_n725_), .Z(G1338gat));
  NAND4_X1  g525(.A1(new_n710_), .A2(new_n383_), .A3(new_n446_), .A4(new_n448_), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n648_), .A2(new_n383_), .A3(new_n601_), .A4(new_n690_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT52), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n728_), .A2(new_n729_), .A3(G106gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n728_), .B2(G106gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT53), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT53), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n734_), .B(new_n727_), .C1(new_n730_), .C2(new_n731_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1339gat));
  NAND3_X1  g535(.A1(new_n386_), .A2(new_n287_), .A3(new_n247_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT120), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT118), .ZN(new_n740_));
  AOI21_X1  g539(.A(KEYINPUT55), .B1(new_n522_), .B2(new_n529_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n511_), .B1(new_n551_), .B2(new_n513_), .ZN(new_n742_));
  AOI21_X1  g541(.A(KEYINPUT12), .B1(new_n482_), .B2(new_n497_), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n425_), .A2(KEYINPUT116), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n742_), .A2(new_n743_), .A3(new_n744_), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n521_), .A2(KEYINPUT55), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n525_), .A2(new_n527_), .A3(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n745_), .B1(new_n744_), .B2(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n535_), .B1(new_n741_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT56), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT117), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n751_), .ZN(new_n753_));
  OAI211_X1 g552(.A(new_n535_), .B(new_n753_), .C1(new_n741_), .C2(new_n748_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n422_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n740_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n538_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT73), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n530_), .A2(new_n537_), .A3(new_n540_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n423_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n761_), .A2(KEYINPUT118), .A3(new_n752_), .A4(new_n754_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n412_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n410_), .A2(new_n411_), .A3(new_n763_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n764_), .B(new_n419_), .C1(new_n414_), .C2(new_n763_), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n421_), .A2(new_n765_), .A3(KEYINPUT119), .ZN(new_n766_));
  AOI21_X1  g565(.A(KEYINPUT119), .B1(new_n421_), .B2(new_n765_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n543_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n757_), .A2(new_n762_), .A3(new_n770_), .ZN(new_n771_));
  AOI211_X1 g570(.A(new_n739_), .B(KEYINPUT57), .C1(new_n771_), .C2(new_n638_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(KEYINPUT57), .A3(new_n638_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT58), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n749_), .B(KEYINPUT56), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n759_), .A2(new_n760_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n769_), .A2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n774_), .B1(new_n775_), .B2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n768_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n749_), .A2(KEYINPUT56), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n749_), .A2(KEYINPUT56), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n779_), .A2(KEYINPUT58), .A3(new_n780_), .A4(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n778_), .A2(new_n782_), .A3(new_n583_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n773_), .A2(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n772_), .A2(new_n784_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n776_), .A2(new_n752_), .A3(new_n422_), .A4(new_n754_), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n786_), .A2(new_n740_), .B1(new_n543_), .B2(new_n769_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n578_), .B1(new_n787_), .B2(new_n762_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n739_), .B1(new_n788_), .B2(KEYINPUT57), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n637_), .B1(new_n785_), .B2(new_n789_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n602_), .A2(new_n423_), .A3(new_n545_), .A4(new_n546_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n791_), .B(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n738_), .B1(new_n790_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(G113gat), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n796_), .A3(new_n422_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT57), .B1(new_n771_), .B2(new_n638_), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n778_), .A2(new_n583_), .A3(new_n782_), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT121), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT121), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n801_), .B(new_n783_), .C1(new_n788_), .C2(KEYINPUT57), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n800_), .A2(new_n802_), .A3(new_n773_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n601_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n793_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n737_), .A2(KEYINPUT59), .ZN(new_n807_));
  AOI22_X1  g606(.A1(new_n794_), .A2(KEYINPUT59), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n808_), .A2(new_n422_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n797_), .B1(new_n809_), .B2(new_n796_), .ZN(G1340gat));
  INV_X1    g609(.A(G120gat), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n548_), .B2(KEYINPUT60), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n795_), .B(new_n812_), .C1(KEYINPUT60), .C2(new_n811_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n808_), .A2(new_n547_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(new_n811_), .ZN(G1341gat));
  INV_X1    g614(.A(G127gat), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n816_), .B1(new_n808_), .B2(new_n637_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n794_), .A2(G127gat), .A3(new_n601_), .ZN(new_n818_));
  OAI21_X1  g617(.A(KEYINPUT122), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n798_), .A2(KEYINPUT120), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n789_), .A2(new_n820_), .A3(new_n773_), .A4(new_n783_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n793_), .B1(new_n821_), .B2(new_n601_), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT59), .B1(new_n822_), .B2(new_n737_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n806_), .A2(new_n807_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n637_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(G127gat), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT122), .ZN(new_n827_));
  INV_X1    g626(.A(new_n818_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n826_), .A2(new_n827_), .A3(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n819_), .A2(new_n829_), .ZN(G1342gat));
  INV_X1    g629(.A(G134gat), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n795_), .A2(new_n831_), .A3(new_n578_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n808_), .A2(new_n583_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n832_), .B1(new_n833_), .B2(new_n831_), .ZN(G1343gat));
  NAND4_X1  g633(.A1(new_n665_), .A2(new_n287_), .A3(new_n383_), .A4(new_n246_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n822_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n422_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n547_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g639(.A1(new_n836_), .A2(new_n637_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(KEYINPUT61), .B(G155gat), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n841_), .B(new_n842_), .ZN(G1346gat));
  INV_X1    g642(.A(G162gat), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n844_), .B1(new_n836_), .B2(new_n583_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT123), .ZN(new_n847_));
  INV_X1    g646(.A(new_n836_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n578_), .A2(new_n844_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n846_), .B(new_n847_), .C1(new_n848_), .C2(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n848_), .A2(new_n849_), .ZN(new_n851_));
  OAI21_X1  g650(.A(KEYINPUT123), .B1(new_n851_), .B2(new_n845_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(G1347gat));
  NOR3_X1   g652(.A1(new_n665_), .A2(new_n383_), .A3(new_n645_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n806_), .A2(new_n422_), .A3(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n855_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n806_), .A2(new_n315_), .A3(new_n422_), .A4(new_n854_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(KEYINPUT62), .B1(new_n855_), .B2(G169gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(KEYINPUT124), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n855_), .A2(G169gat), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT62), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT124), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n863_), .A2(new_n864_), .A3(new_n857_), .A4(new_n856_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n860_), .A2(new_n865_), .ZN(G1348gat));
  NAND2_X1  g665(.A1(new_n806_), .A2(new_n854_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n547_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n822_), .A2(new_n383_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n665_), .A2(new_n645_), .ZN(new_n871_));
  AND3_X1   g670(.A1(new_n871_), .A2(new_n547_), .A3(G176gat), .ZN(new_n872_));
  AOI22_X1  g671(.A1(new_n869_), .A2(new_n229_), .B1(new_n870_), .B2(new_n872_), .ZN(G1349gat));
  NOR3_X1   g672(.A1(new_n867_), .A2(new_n215_), .A3(new_n601_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n870_), .A2(new_n637_), .A3(new_n871_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n211_), .B2(new_n875_), .ZN(G1350gat));
  OAI21_X1  g675(.A(G190gat), .B1(new_n867_), .B2(new_n642_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n578_), .A2(new_n218_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n867_), .B2(new_n878_), .ZN(G1351gat));
  NAND2_X1  g678(.A1(new_n369_), .A2(new_n246_), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n880_), .A2(KEYINPUT125), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(KEYINPUT125), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n881_), .A2(new_n382_), .A3(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n822_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n422_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g685(.A(new_n884_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n548_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT126), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n889_), .B2(new_n288_), .ZN(new_n890_));
  XOR2_X1   g689(.A(KEYINPUT126), .B(G204gat), .Z(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n888_), .B2(new_n891_), .ZN(G1353gat));
  INV_X1    g691(.A(KEYINPUT127), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT63), .B(G211gat), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n884_), .A2(new_n637_), .A3(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n887_), .A2(new_n601_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n893_), .B(new_n895_), .C1(new_n896_), .C2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n895_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n897_), .B1(new_n884_), .B2(new_n637_), .ZN(new_n900_));
  OAI21_X1  g699(.A(KEYINPUT127), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n898_), .A2(new_n901_), .ZN(G1354gat));
  OR3_X1    g701(.A1(new_n887_), .A2(G218gat), .A3(new_n638_), .ZN(new_n903_));
  OAI21_X1  g702(.A(G218gat), .B1(new_n887_), .B2(new_n642_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1355gat));
endmodule


