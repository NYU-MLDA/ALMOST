//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 1 1 1 0 1 1 0 1 1 0 1 0 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 1 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n794_, new_n795_, new_n797_,
    new_n798_, new_n799_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n945_, new_n946_, new_n947_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n954_, new_n955_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n962_, new_n963_;
  NOR2_X1   g000(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT64), .ZN(new_n204_));
  NAND2_X1  g003(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n205_), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT64), .B1(new_n207_), .B2(new_n202_), .ZN(new_n208_));
  AOI21_X1  g007(.A(G106gat), .B1(new_n206_), .B2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  AND2_X1   g010(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(G85gat), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n211_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT66), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G99gat), .A2(G106gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT6), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NOR4_X1   g021(.A1(new_n209_), .A2(new_n216_), .A3(new_n217_), .A4(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n214_), .A2(new_n215_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n222_), .B1(new_n224_), .B2(new_n210_), .ZN(new_n225_));
  INV_X1    g024(.A(G106gat), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n204_), .B1(new_n203_), .B2(new_n205_), .ZN(new_n227_));
  NOR3_X1   g026(.A1(new_n207_), .A2(new_n202_), .A3(KEYINPUT64), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n226_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(KEYINPUT66), .B1(new_n225_), .B2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT8), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT7), .ZN(new_n232_));
  INV_X1    g031(.A(G99gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(new_n233_), .A3(new_n226_), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n222_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n234_), .A2(KEYINPUT68), .A3(new_n235_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n238_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  XOR2_X1   g040(.A(G85gat), .B(G92gat), .Z(new_n242_));
  AOI21_X1  g041(.A(new_n231_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n231_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n236_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(new_n239_), .A3(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT67), .B1(new_n236_), .B2(new_n222_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n244_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  OAI22_X1  g048(.A1(new_n223_), .A2(new_n230_), .B1(new_n243_), .B2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G29gat), .B(G36gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G43gat), .B(G50gat), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n251_), .A2(new_n252_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT73), .B(KEYINPUT15), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT35), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G232gat), .A2(G233gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT34), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  AOI22_X1  g061(.A1(new_n250_), .A2(new_n258_), .B1(new_n259_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT74), .ZN(new_n264_));
  INV_X1    g063(.A(new_n256_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n264_), .B1(new_n250_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n244_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n246_), .B1(new_n245_), .B2(new_n239_), .ZN(new_n268_));
  NOR3_X1   g067(.A1(new_n236_), .A2(new_n222_), .A3(KEYINPUT67), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n267_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n242_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n222_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n271_), .B1(new_n272_), .B2(new_n240_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n270_), .B1(new_n231_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n215_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT65), .B(G92gat), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n275_), .B1(new_n276_), .B2(G85gat), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n239_), .B1(new_n277_), .B2(new_n211_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n217_), .B1(new_n278_), .B2(new_n209_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n225_), .A2(KEYINPUT66), .A3(new_n229_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n274_), .A2(new_n281_), .A3(KEYINPUT74), .A4(new_n256_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n263_), .A2(new_n266_), .A3(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n262_), .A2(new_n259_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(G190gat), .B(G218gat), .Z(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT75), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G134gat), .B(G162gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n289_), .A2(KEYINPUT36), .ZN(new_n290_));
  INV_X1    g089(.A(new_n284_), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n263_), .A2(new_n266_), .A3(new_n291_), .A4(new_n282_), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n285_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n289_), .B(KEYINPUT36), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n285_), .A2(new_n292_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n294_), .B1(new_n295_), .B2(KEYINPUT77), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT77), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n285_), .A2(new_n297_), .A3(new_n292_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n293_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n300_), .A2(KEYINPUT100), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n300_), .A2(KEYINPUT100), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G127gat), .B(G134gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G113gat), .B(G120gat), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n305_), .A2(KEYINPUT87), .ZN(new_n306_));
  INV_X1    g105(.A(G120gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(G113gat), .ZN(new_n308_));
  INV_X1    g107(.A(G113gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(G120gat), .ZN(new_n310_));
  AND3_X1   g109(.A1(new_n308_), .A2(new_n310_), .A3(KEYINPUT87), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n304_), .B1(new_n306_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n308_), .A2(new_n310_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT87), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n305_), .A2(KEYINPUT87), .ZN(new_n316_));
  INV_X1    g115(.A(new_n304_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(KEYINPUT88), .B1(new_n312_), .B2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n317_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT88), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n319_), .A2(new_n322_), .ZN(new_n323_));
  XOR2_X1   g122(.A(KEYINPUT89), .B(KEYINPUT31), .Z(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G71gat), .B(G99gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(G43gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G227gat), .A2(G233gat), .ZN(new_n329_));
  INV_X1    g128(.A(G15gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n328_), .B(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(G190gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT26), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT82), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT25), .B(G183gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT83), .B(KEYINPUT26), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n336_), .B(new_n337_), .C1(new_n333_), .C2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G183gat), .A2(G190gat), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT23), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(G169gat), .ZN(new_n345_));
  INV_X1    g144(.A(G176gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  OR2_X1    g146(.A1(new_n347_), .A2(KEYINPUT24), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G169gat), .A2(G176gat), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n347_), .A2(KEYINPUT24), .A3(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n344_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n339_), .A2(new_n352_), .ZN(new_n353_));
  OR2_X1    g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n342_), .A2(new_n354_), .A3(new_n343_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT85), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT85), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n342_), .A2(new_n354_), .A3(new_n357_), .A4(new_n343_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n345_), .A2(KEYINPUT22), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT22), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(G169gat), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n359_), .A2(new_n361_), .A3(new_n346_), .ZN(new_n362_));
  AND3_X1   g161(.A1(new_n362_), .A2(KEYINPUT84), .A3(new_n349_), .ZN(new_n363_));
  AOI21_X1  g162(.A(KEYINPUT84), .B1(new_n362_), .B2(new_n349_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n356_), .B(new_n358_), .C1(new_n363_), .C2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n353_), .A2(KEYINPUT30), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(KEYINPUT30), .B1(new_n353_), .B2(new_n365_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT86), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n353_), .A2(new_n365_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT30), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT86), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(new_n373_), .A3(new_n366_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n332_), .B1(new_n369_), .B2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n373_), .B1(new_n372_), .B2(new_n366_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n332_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n326_), .B1(new_n375_), .B2(new_n378_), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n367_), .A2(KEYINPUT86), .A3(new_n368_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n377_), .B1(new_n380_), .B2(new_n376_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n369_), .A2(new_n332_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n381_), .A2(new_n382_), .A3(new_n325_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n379_), .A2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G22gat), .B(G50gat), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT28), .ZN(new_n387_));
  XOR2_X1   g186(.A(G155gat), .B(G162gat), .Z(new_n388_));
  NAND3_X1  g187(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT90), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT3), .ZN(new_n391_));
  INV_X1    g190(.A(G141gat), .ZN(new_n392_));
  INV_X1    g191(.A(G148gat), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n391_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G141gat), .A2(G148gat), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT2), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n394_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n388_), .B1(new_n390_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n392_), .A2(new_n393_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT1), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n402_), .B1(G155gat), .B2(G162gat), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(G155gat), .A3(G162gat), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n404_), .B1(G155gat), .B2(G162gat), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n401_), .B(new_n395_), .C1(new_n403_), .C2(new_n405_), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n400_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT29), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n387_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n400_), .A2(new_n406_), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n411_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n386_), .B1(new_n410_), .B2(new_n413_), .ZN(new_n414_));
  NOR3_X1   g213(.A1(new_n409_), .A2(new_n412_), .A3(new_n385_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(G228gat), .ZN(new_n417_));
  INV_X1    g216(.A(G233gat), .ZN(new_n418_));
  NOR3_X1   g217(.A1(new_n417_), .A2(new_n418_), .A3(KEYINPUT92), .ZN(new_n419_));
  OAI21_X1  g218(.A(KEYINPUT92), .B1(new_n417_), .B2(new_n418_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n408_), .B1(new_n400_), .B2(new_n406_), .ZN(new_n421_));
  OR2_X1    g220(.A1(G197gat), .A2(G204gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G197gat), .A2(G204gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT21), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n422_), .A2(KEYINPUT21), .A3(new_n423_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G211gat), .B(G218gat), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n426_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n427_), .A2(new_n428_), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n420_), .B1(new_n421_), .B2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G78gat), .B(G106gat), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n420_), .B(new_n433_), .C1(new_n421_), .C2(new_n431_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n419_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n435_), .A2(new_n419_), .A3(new_n436_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n416_), .A2(new_n438_), .A3(KEYINPUT91), .A4(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(KEYINPUT91), .ZN(new_n441_));
  OAI22_X1  g240(.A1(new_n441_), .A2(new_n437_), .B1(new_n415_), .B2(new_n414_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n440_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n384_), .A2(new_n443_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n440_), .A2(new_n379_), .A3(new_n383_), .A4(new_n442_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n431_), .B1(new_n353_), .B2(new_n365_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G226gat), .A2(G233gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT19), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n349_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT22), .B(G169gat), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n451_), .B1(new_n452_), .B2(new_n346_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n355_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(KEYINPUT26), .B(G190gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n337_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n454_), .B1(new_n351_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n429_), .A2(new_n430_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n450_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT20), .ZN(new_n461_));
  OR3_X1    g260(.A1(new_n447_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n449_), .B(KEYINPUT93), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n353_), .A2(new_n365_), .A3(new_n431_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n461_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n464_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G8gat), .B(G36gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G64gat), .B(G92gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n462_), .A2(new_n468_), .A3(new_n473_), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n465_), .A2(new_n466_), .A3(new_n464_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n447_), .A2(new_n461_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n459_), .B1(new_n458_), .B2(KEYINPUT98), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n477_), .B1(KEYINPUT98), .B2(new_n458_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n475_), .B1(new_n479_), .B2(new_n449_), .ZN(new_n480_));
  OAI211_X1 g279(.A(KEYINPUT27), .B(new_n474_), .C1(new_n480_), .C2(new_n473_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n473_), .ZN(new_n482_));
  NOR3_X1   g281(.A1(new_n447_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n482_), .B1(new_n483_), .B2(new_n467_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n474_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT27), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n481_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G225gat), .A2(G233gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT96), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT4), .ZN(new_n491_));
  NOR3_X1   g290(.A1(new_n306_), .A2(new_n311_), .A3(new_n304_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n321_), .B1(new_n492_), .B2(new_n320_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n493_), .B(new_n411_), .C1(new_n321_), .C2(new_n320_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT95), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n495_), .B1(new_n492_), .B2(new_n320_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n312_), .A2(KEYINPUT95), .A3(new_n318_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(new_n407_), .A3(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n491_), .B1(new_n494_), .B2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(KEYINPUT4), .B1(new_n323_), .B2(new_n411_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n490_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n494_), .A2(new_n489_), .A3(new_n498_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G1gat), .B(G29gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(G85gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(KEYINPUT0), .B(G57gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n503_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n507_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n501_), .A2(new_n502_), .A3(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n488_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n446_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n443_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n489_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n494_), .A2(new_n498_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT4), .ZN(new_n517_));
  INV_X1    g316(.A(new_n500_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n515_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n490_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n507_), .B1(new_n516_), .B2(new_n520_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n474_), .B(new_n484_), .C1(new_n519_), .C2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n510_), .A2(KEYINPUT33), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT33), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n501_), .A2(new_n524_), .A3(new_n502_), .A4(new_n509_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n522_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n473_), .A2(KEYINPUT32), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT97), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n462_), .A2(new_n468_), .A3(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n480_), .A2(new_n528_), .A3(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n462_), .A2(new_n468_), .A3(KEYINPUT97), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n527_), .ZN(new_n533_));
  AOI22_X1  g332(.A1(new_n508_), .A2(new_n510_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n384_), .B(new_n514_), .C1(new_n526_), .C2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n513_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n303_), .A2(KEYINPUT101), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(KEYINPUT101), .B1(new_n303_), .B2(new_n536_), .ZN(new_n539_));
  OR2_X1    g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G57gat), .B(G64gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT11), .ZN(new_n542_));
  XOR2_X1   g341(.A(G71gat), .B(G78gat), .Z(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n542_), .A2(new_n543_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n541_), .A2(KEYINPUT11), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n544_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n250_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(KEYINPUT69), .B(KEYINPUT12), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(G230gat), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n552_), .A2(new_n418_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n243_), .ZN(new_n554_));
  AOI22_X1  g353(.A1(new_n554_), .A2(new_n270_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n548_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n553_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n250_), .A2(KEYINPUT12), .A3(new_n548_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n551_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n274_), .A2(new_n281_), .A3(new_n556_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n549_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(new_n553_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G176gat), .B(G204gat), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT71), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(G120gat), .B(G148gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n568_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n559_), .A2(new_n562_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT72), .ZN(new_n574_));
  INV_X1    g373(.A(new_n570_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n567_), .A2(new_n568_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n574_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n569_), .A2(KEYINPUT72), .A3(new_n570_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n579_), .B1(new_n559_), .B2(new_n562_), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT13), .B1(new_n573_), .B2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n559_), .A2(new_n562_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n579_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT13), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(new_n585_), .A3(new_n572_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n581_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G127gat), .B(G155gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G183gat), .B(G211gat), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n591_), .A2(new_n592_), .ZN(new_n594_));
  OR3_X1    g393(.A1(new_n593_), .A2(new_n594_), .A3(KEYINPUT17), .ZN(new_n595_));
  OAI21_X1  g394(.A(KEYINPUT17), .B1(new_n593_), .B2(new_n594_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(G1gat), .ZN(new_n598_));
  INV_X1    g397(.A(G8gat), .ZN(new_n599_));
  OAI21_X1  g398(.A(KEYINPUT14), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  OR2_X1    g399(.A1(KEYINPUT78), .A2(G15gat), .ZN(new_n601_));
  NAND2_X1  g400(.A1(KEYINPUT78), .A2(G15gat), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n601_), .A2(G22gat), .A3(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(G22gat), .B1(new_n601_), .B2(new_n602_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n600_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  XOR2_X1   g404(.A(G1gat), .B(G8gat), .Z(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n606_), .B(new_n600_), .C1(new_n603_), .C2(new_n604_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(G231gat), .A3(G233gat), .ZN(new_n611_));
  INV_X1    g410(.A(G231gat), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n608_), .B(new_n609_), .C1(new_n612_), .C2(new_n418_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n556_), .B1(new_n611_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n611_), .A2(new_n613_), .A3(new_n556_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n597_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n616_), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n618_), .A2(new_n614_), .A3(new_n596_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT81), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n254_), .A2(KEYINPUT80), .A3(new_n255_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT80), .ZN(new_n624_));
  INV_X1    g423(.A(new_n255_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n624_), .B1(new_n625_), .B2(new_n253_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n623_), .A2(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n627_), .A2(new_n610_), .ZN(new_n628_));
  AOI22_X1  g427(.A1(new_n623_), .A2(new_n626_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n622_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(G229gat), .A2(G233gat), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n627_), .A2(new_n610_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n608_), .A2(new_n623_), .A3(new_n626_), .A4(new_n609_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n633_), .A2(new_n634_), .A3(KEYINPUT81), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n630_), .A2(new_n632_), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n258_), .A2(new_n610_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n637_), .A2(new_n631_), .A3(new_n634_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G113gat), .B(G141gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(G169gat), .B(G197gat), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n639_), .B(new_n640_), .Z(new_n641_));
  NAND3_X1  g440(.A1(new_n636_), .A2(new_n638_), .A3(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n641_), .B1(new_n636_), .B2(new_n638_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n588_), .A2(new_n621_), .A3(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n540_), .A2(new_n511_), .A3(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(G1gat), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n588_), .A2(new_n645_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n649_), .A2(new_n536_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n294_), .B1(new_n285_), .B2(new_n292_), .ZN(new_n651_));
  OAI21_X1  g450(.A(KEYINPUT37), .B1(new_n293_), .B2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT76), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT76), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n654_), .B(KEYINPUT37), .C1(new_n293_), .C2(new_n651_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT37), .ZN(new_n656_));
  AOI22_X1  g455(.A1(new_n653_), .A2(new_n655_), .B1(new_n299_), .B2(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n657_), .A2(new_n621_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n650_), .A2(new_n658_), .ZN(new_n659_));
  XOR2_X1   g458(.A(new_n511_), .B(KEYINPUT99), .Z(new_n660_));
  NAND3_X1  g459(.A1(new_n659_), .A2(new_n598_), .A3(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT38), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n648_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n648_), .A2(KEYINPUT102), .A3(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1324gat));
  NAND3_X1  g466(.A1(new_n659_), .A2(new_n599_), .A3(new_n488_), .ZN(new_n668_));
  OAI211_X1 g467(.A(new_n488_), .B(new_n646_), .C1(new_n538_), .C2(new_n539_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT39), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n669_), .A2(new_n670_), .A3(G8gat), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n669_), .B2(G8gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n668_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT40), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  OAI211_X1 g474(.A(KEYINPUT40), .B(new_n668_), .C1(new_n671_), .C2(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1325gat));
  INV_X1    g476(.A(new_n384_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n659_), .A2(new_n330_), .A3(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n540_), .A2(new_n678_), .A3(new_n646_), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n680_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT41), .B1(new_n680_), .B2(G15gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n679_), .B1(new_n681_), .B2(new_n682_), .ZN(G1326gat));
  INV_X1    g482(.A(G22gat), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n659_), .A2(new_n684_), .A3(new_n443_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n540_), .A2(new_n443_), .A3(new_n646_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n686_), .A2(G22gat), .A3(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n686_), .B2(G22gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n685_), .B1(new_n688_), .B2(new_n689_), .ZN(G1327gat));
  NOR2_X1   g489(.A1(new_n300_), .A2(new_n620_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n650_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(G29gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n692_), .A2(new_n693_), .A3(new_n511_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n660_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n649_), .A2(new_n621_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n657_), .A2(new_n536_), .A3(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n657_), .B2(new_n536_), .ZN(new_n700_));
  OAI211_X1 g499(.A(KEYINPUT44), .B(new_n697_), .C1(new_n699_), .C2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n653_), .A2(new_n655_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n299_), .A2(new_n656_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n531_), .A2(new_n533_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n511_), .A2(new_n707_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n523_), .A2(new_n525_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n708_), .B1(new_n709_), .B2(new_n522_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n678_), .A2(new_n443_), .ZN(new_n711_));
  AOI22_X1  g510(.A1(new_n710_), .A2(new_n711_), .B1(new_n446_), .B2(new_n512_), .ZN(new_n712_));
  OAI21_X1  g511(.A(KEYINPUT43), .B1(new_n706_), .B2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n657_), .A2(new_n536_), .A3(new_n698_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n696_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n703_), .B1(new_n715_), .B2(KEYINPUT44), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n697_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n717_), .A2(KEYINPUT104), .A3(new_n718_), .ZN(new_n719_));
  AOI211_X1 g518(.A(new_n695_), .B(new_n702_), .C1(new_n716_), .C2(new_n719_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n720_), .A2(KEYINPUT105), .ZN(new_n721_));
  OAI21_X1  g520(.A(G29gat), .B1(new_n720_), .B2(KEYINPUT105), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n694_), .B1(new_n721_), .B2(new_n722_), .ZN(G1328gat));
  INV_X1    g522(.A(KEYINPUT46), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n724_), .A2(KEYINPUT107), .ZN(new_n725_));
  INV_X1    g524(.A(G36gat), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n716_), .A2(new_n719_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n488_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n702_), .A2(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n726_), .B1(new_n727_), .B2(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n692_), .A2(new_n726_), .A3(new_n488_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n731_), .B(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n725_), .B1(new_n730_), .B2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n724_), .A2(KEYINPUT107), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n734_), .B(new_n735_), .ZN(G1329gat));
  AND4_X1   g535(.A1(G43gat), .A2(new_n727_), .A3(new_n678_), .A4(new_n701_), .ZN(new_n737_));
  AOI21_X1  g536(.A(G43gat), .B1(new_n692_), .B2(new_n678_), .ZN(new_n738_));
  OR3_X1    g537(.A1(new_n737_), .A2(KEYINPUT47), .A3(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(KEYINPUT47), .B1(new_n737_), .B2(new_n738_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1330gat));
  INV_X1    g540(.A(G50gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n692_), .A2(new_n742_), .A3(new_n443_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n514_), .B1(new_n715_), .B2(KEYINPUT44), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n715_), .A2(new_n703_), .A3(KEYINPUT44), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT104), .B1(new_n717_), .B2(new_n718_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n744_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n742_), .B1(new_n747_), .B2(KEYINPUT108), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n727_), .A2(new_n749_), .A3(new_n744_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n748_), .A2(KEYINPUT109), .A3(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(KEYINPUT109), .B1(new_n748_), .B2(new_n750_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n743_), .B1(new_n751_), .B2(new_n752_), .ZN(G1331gat));
  INV_X1    g552(.A(new_n645_), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n587_), .A2(new_n621_), .A3(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n755_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT110), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  OAI211_X1 g557(.A(KEYINPUT110), .B(new_n755_), .C1(new_n538_), .C2(new_n539_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n758_), .A2(G57gat), .A3(new_n511_), .A4(new_n759_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n760_), .A2(KEYINPUT111), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n760_), .A2(KEYINPUT111), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n587_), .A2(new_n754_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n536_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n658_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(G57gat), .B1(new_n766_), .B2(new_n660_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n761_), .A2(new_n762_), .A3(new_n767_), .ZN(G1332gat));
  OR3_X1    g567(.A1(new_n765_), .A2(G64gat), .A3(new_n728_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n758_), .A2(new_n488_), .A3(new_n759_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n770_), .A2(G64gat), .A3(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n770_), .B2(G64gat), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n772_), .B2(new_n773_), .ZN(G1333gat));
  OR3_X1    g573(.A1(new_n765_), .A2(G71gat), .A3(new_n384_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n758_), .A2(new_n678_), .A3(new_n759_), .ZN(new_n776_));
  XOR2_X1   g575(.A(KEYINPUT113), .B(KEYINPUT49), .Z(new_n777_));
  AND3_X1   g576(.A1(new_n776_), .A2(G71gat), .A3(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n776_), .B2(G71gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(G1334gat));
  OR3_X1    g579(.A1(new_n765_), .A2(G78gat), .A3(new_n514_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n758_), .A2(new_n443_), .A3(new_n759_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n782_), .A2(new_n783_), .A3(G78gat), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n782_), .B2(G78gat), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n781_), .B1(new_n784_), .B2(new_n785_), .ZN(G1335gat));
  AND2_X1   g585(.A1(new_n764_), .A2(new_n691_), .ZN(new_n787_));
  AOI21_X1  g586(.A(G85gat), .B1(new_n787_), .B2(new_n660_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n763_), .A2(new_n621_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n511_), .A2(G85gat), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n791_), .B(KEYINPUT114), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n788_), .B1(new_n790_), .B2(new_n792_), .ZN(G1336gat));
  AOI21_X1  g592(.A(G92gat), .B1(new_n787_), .B2(new_n488_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n488_), .A2(new_n276_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(new_n790_), .B2(new_n795_), .ZN(G1337gat));
  AOI21_X1  g595(.A(new_n233_), .B1(new_n790_), .B2(new_n678_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n384_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n797_), .B1(new_n787_), .B2(new_n798_), .ZN(new_n799_));
  XOR2_X1   g598(.A(new_n799_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g599(.A(KEYINPUT115), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802_));
  OAI21_X1  g601(.A(G106gat), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n803_), .B1(new_n790_), .B2(new_n443_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n801_), .A2(new_n802_), .ZN(new_n805_));
  OR2_X1    g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n805_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n787_), .A2(new_n226_), .A3(new_n443_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n806_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g609(.A1(new_n660_), .A2(new_n728_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n811_), .A2(KEYINPUT59), .A3(new_n445_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT58), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n556_), .B1(new_n274_), .B2(new_n281_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n550_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n558_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n560_), .B1(new_n552_), .B2(new_n418_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n814_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n558_), .B(new_n560_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n553_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n551_), .A2(new_n557_), .A3(KEYINPUT55), .A4(new_n558_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n819_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT56), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n583_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n630_), .A2(new_n631_), .A3(new_n635_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n628_), .A2(new_n631_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n641_), .B1(new_n827_), .B2(new_n637_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n572_), .A2(new_n642_), .A3(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n825_), .A2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n824_), .B1(new_n823_), .B2(new_n583_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n813_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n832_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n834_), .A2(KEYINPUT58), .A3(new_n825_), .A4(new_n830_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n704_), .A2(new_n833_), .A3(new_n835_), .A4(new_n705_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n642_), .B(new_n829_), .C1(new_n573_), .C2(new_n580_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n824_), .A2(KEYINPUT117), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n823_), .A2(new_n583_), .A3(new_n838_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n559_), .A2(new_n562_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n636_), .A2(new_n638_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n641_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n840_), .A2(new_n571_), .B1(new_n843_), .B2(new_n642_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n839_), .A2(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n838_), .B1(new_n823_), .B2(new_n583_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n837_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n847_), .A2(new_n848_), .A3(new_n300_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n848_), .B1(new_n847_), .B2(new_n300_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n836_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n851_), .A2(new_n621_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n621_), .A2(new_n643_), .A3(new_n644_), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n573_), .A2(new_n580_), .A3(KEYINPUT13), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n585_), .B1(new_n584_), .B2(new_n572_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n853_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n587_), .A2(KEYINPUT116), .A3(new_n853_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n860_), .A2(new_n861_), .A3(new_n706_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n861_), .B1(new_n860_), .B2(new_n706_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n812_), .B1(new_n852_), .B2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n620_), .B1(new_n851_), .B2(KEYINPUT118), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n867_), .B(new_n836_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n864_), .B1(new_n866_), .B2(new_n868_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n869_), .A2(new_n445_), .A3(new_n811_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT59), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n865_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(G113gat), .B1(new_n872_), .B2(new_n645_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n870_), .A2(new_n309_), .A3(new_n754_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1340gat));
  OAI21_X1  g674(.A(G120gat), .B1(new_n872_), .B2(new_n587_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n307_), .B1(new_n587_), .B2(KEYINPUT60), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n870_), .B(new_n877_), .C1(KEYINPUT60), .C2(new_n307_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(G1341gat));
  OAI21_X1  g678(.A(G127gat), .B1(new_n872_), .B2(new_n621_), .ZN(new_n880_));
  INV_X1    g679(.A(G127gat), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n870_), .A2(new_n881_), .A3(new_n620_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(G1342gat));
  NAND2_X1  g682(.A1(new_n657_), .A2(G134gat), .ZN(new_n884_));
  XOR2_X1   g683(.A(new_n884_), .B(KEYINPUT119), .Z(new_n885_));
  OAI211_X1 g684(.A(new_n865_), .B(new_n885_), .C1(new_n870_), .C2(new_n871_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n303_), .ZN(new_n888_));
  AOI21_X1  g687(.A(G134gat), .B1(new_n870_), .B2(new_n888_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n887_), .A2(new_n889_), .ZN(G1343gat));
  NAND2_X1  g689(.A1(new_n851_), .A2(KEYINPUT118), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n891_), .A2(new_n621_), .A3(new_n868_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n864_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n811_), .A2(new_n444_), .ZN(new_n895_));
  XOR2_X1   g694(.A(new_n895_), .B(KEYINPUT120), .Z(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n645_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(new_n392_), .ZN(G1344gat));
  NOR2_X1   g698(.A1(new_n897_), .A2(new_n587_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(new_n393_), .ZN(G1345gat));
  NOR2_X1   g700(.A1(new_n897_), .A2(new_n621_), .ZN(new_n902_));
  XOR2_X1   g701(.A(KEYINPUT61), .B(G155gat), .Z(new_n903_));
  XNOR2_X1  g702(.A(new_n902_), .B(new_n903_), .ZN(G1346gat));
  INV_X1    g703(.A(G162gat), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n894_), .A2(new_n896_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n905_), .B1(new_n906_), .B2(new_n657_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n888_), .A2(new_n905_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n897_), .A2(new_n908_), .ZN(new_n909_));
  OAI21_X1  g708(.A(KEYINPUT121), .B1(new_n907_), .B2(new_n909_), .ZN(new_n910_));
  OAI21_X1  g709(.A(G162gat), .B1(new_n897_), .B2(new_n706_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n911_), .B(new_n912_), .C1(new_n897_), .C2(new_n908_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n910_), .A2(new_n913_), .ZN(G1347gat));
  INV_X1    g713(.A(KEYINPUT62), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n728_), .A2(new_n384_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n695_), .A2(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  OAI211_X1 g717(.A(new_n514_), .B(new_n918_), .C1(new_n852_), .C2(new_n864_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n919_), .A2(new_n645_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n915_), .B1(new_n920_), .B2(new_n345_), .ZN(new_n921_));
  OAI211_X1 g720(.A(KEYINPUT62), .B(G169gat), .C1(new_n919_), .C2(new_n645_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n920_), .A2(new_n452_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n921_), .A2(new_n922_), .A3(new_n923_), .ZN(G1348gat));
  OAI21_X1  g723(.A(new_n346_), .B1(new_n919_), .B2(new_n587_), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n443_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n917_), .A2(new_n346_), .A3(new_n587_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n926_), .B1(new_n927_), .B2(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n928_), .ZN(new_n930_));
  NOR4_X1   g729(.A1(new_n869_), .A2(KEYINPUT122), .A3(new_n443_), .A4(new_n930_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n925_), .B1(new_n929_), .B2(new_n931_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  OAI211_X1 g733(.A(KEYINPUT123), .B(new_n925_), .C1(new_n929_), .C2(new_n931_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n934_), .A2(new_n935_), .ZN(G1349gat));
  OAI21_X1  g735(.A(new_n514_), .B1(new_n852_), .B2(new_n864_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n917_), .A2(new_n621_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n938_), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n937_), .A2(new_n337_), .A3(new_n939_), .ZN(new_n940_));
  AOI21_X1  g739(.A(KEYINPUT124), .B1(new_n927_), .B2(new_n938_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n941_), .A2(G183gat), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n927_), .A2(KEYINPUT124), .A3(new_n938_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n940_), .B1(new_n942_), .B2(new_n943_), .ZN(G1350gat));
  OAI21_X1  g743(.A(G190gat), .B1(new_n919_), .B2(new_n706_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n888_), .A2(new_n455_), .ZN(new_n946_));
  XOR2_X1   g745(.A(new_n946_), .B(KEYINPUT125), .Z(new_n947_));
  OAI21_X1  g746(.A(new_n945_), .B1(new_n947_), .B2(new_n919_), .ZN(G1351gat));
  NOR3_X1   g747(.A1(new_n728_), .A2(new_n444_), .A3(new_n511_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n894_), .A2(new_n949_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n950_), .A2(new_n645_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(KEYINPUT126), .B(G197gat), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n951_), .B(new_n952_), .ZN(G1352gat));
  INV_X1    g752(.A(new_n950_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n954_), .A2(new_n588_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n955_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g755(.A(new_n621_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n957_));
  XNOR2_X1  g756(.A(new_n957_), .B(KEYINPUT127), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n954_), .A2(new_n958_), .ZN(new_n959_));
  OR2_X1    g758(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n959_), .B(new_n960_), .ZN(G1354gat));
  OR3_X1    g760(.A1(new_n950_), .A2(G218gat), .A3(new_n303_), .ZN(new_n962_));
  OAI21_X1  g761(.A(G218gat), .B1(new_n950_), .B2(new_n706_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n962_), .A2(new_n963_), .ZN(G1355gat));
endmodule


