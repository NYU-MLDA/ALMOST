//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 1 1 1 1 0 1 0 0 1 1 0 1 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n646_, new_n647_,
    new_n648_, new_n650_, new_n651_, new_n652_, new_n653_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n865_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n888_, new_n890_, new_n891_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n203_), .A2(KEYINPUT89), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT29), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT81), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT81), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n208_), .A2(G155gat), .A3(G162gat), .ZN(new_n209_));
  INV_X1    g008(.A(G155gat), .ZN(new_n210_));
  INV_X1    g009(.A(G162gat), .ZN(new_n211_));
  AOI22_X1  g010(.A1(new_n207_), .A2(new_n209_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G141gat), .ZN(new_n213_));
  INV_X1    g012(.A(G148gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n213_), .A2(new_n214_), .A3(KEYINPUT3), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n216_), .B1(G141gat), .B2(G148gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT83), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n222_), .B1(new_n219_), .B2(KEYINPUT83), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n212_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT84), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G141gat), .A2(G148gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT2), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT83), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n218_), .A2(new_n230_), .A3(new_n222_), .A4(new_n220_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT84), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(new_n232_), .A3(new_n212_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n225_), .A2(new_n233_), .ZN(new_n234_));
  XOR2_X1   g033(.A(G141gat), .B(G148gat), .Z(new_n235_));
  NAND2_X1  g034(.A1(new_n210_), .A2(new_n211_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT1), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n207_), .A2(new_n209_), .A3(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n237_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT82), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n236_), .B(new_n238_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n239_), .A2(new_n240_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n235_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n205_), .B1(new_n234_), .B2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G228gat), .A2(G233gat), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  OR2_X1    g045(.A1(G197gat), .A2(G204gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G197gat), .A2(G204gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT21), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT87), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT87), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n249_), .A2(new_n253_), .A3(new_n250_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n247_), .A2(KEYINPUT21), .A3(new_n248_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G211gat), .B(G218gat), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n252_), .A2(new_n254_), .A3(new_n255_), .A4(new_n256_), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n255_), .A2(new_n256_), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NOR3_X1   g058(.A1(new_n244_), .A2(new_n246_), .A3(new_n259_), .ZN(new_n260_));
  AND3_X1   g059(.A1(new_n231_), .A2(new_n232_), .A3(new_n212_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n232_), .B1(new_n231_), .B2(new_n212_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n243_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT29), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n257_), .A2(new_n258_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n245_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n204_), .B1(new_n260_), .B2(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n246_), .B1(new_n244_), .B2(new_n259_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n264_), .A2(new_n245_), .A3(new_n265_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n268_), .B(new_n269_), .C1(KEYINPUT89), .C2(new_n203_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n243_), .B(new_n205_), .C1(new_n262_), .C2(new_n261_), .ZN(new_n271_));
  XOR2_X1   g070(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(G22gat), .B(G50gat), .Z(new_n274_));
  INV_X1    g073(.A(new_n272_), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n234_), .A2(new_n205_), .A3(new_n243_), .A4(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n273_), .A2(new_n274_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n274_), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n207_), .A2(new_n209_), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT82), .B1(new_n279_), .B2(new_n237_), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n238_), .A2(new_n236_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n239_), .A2(new_n240_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  AOI22_X1  g082(.A1(new_n225_), .A2(new_n233_), .B1(new_n283_), .B2(new_n235_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n275_), .B1(new_n284_), .B2(new_n205_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n271_), .A2(new_n272_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n278_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n267_), .A2(new_n270_), .A3(new_n277_), .A4(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT86), .ZN(new_n289_));
  AND3_X1   g088(.A1(new_n273_), .A2(new_n274_), .A3(new_n276_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n274_), .B1(new_n273_), .B2(new_n276_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n289_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n287_), .A2(KEYINPUT86), .A3(new_n277_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT88), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n294_), .B(new_n202_), .C1(new_n260_), .C2(new_n266_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n292_), .A2(new_n293_), .A3(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n268_), .A2(new_n269_), .A3(new_n203_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT88), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n203_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n288_), .B1(new_n296_), .B2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G1gat), .B(G29gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(G85gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT0), .B(G57gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(G134gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(G127gat), .ZN(new_n307_));
  INV_X1    g106(.A(G127gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(G134gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(G120gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(G113gat), .ZN(new_n312_));
  INV_X1    g111(.A(G113gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(G120gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n310_), .A2(new_n315_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n307_), .A2(new_n309_), .A3(new_n312_), .A4(new_n314_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT80), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT4), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n263_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G225gat), .A2(G233gat), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  AND3_X1   g124(.A1(new_n316_), .A2(KEYINPUT91), .A3(new_n317_), .ZN(new_n326_));
  AOI21_X1  g125(.A(KEYINPUT91), .B1(new_n316_), .B2(new_n317_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n328_), .B(new_n243_), .C1(new_n262_), .C2(new_n261_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n318_), .B(KEYINPUT80), .ZN(new_n330_));
  OAI211_X1 g129(.A(new_n329_), .B(KEYINPUT4), .C1(new_n284_), .C2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT92), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n263_), .A2(new_n320_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT92), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n333_), .A2(new_n334_), .A3(KEYINPUT4), .A4(new_n329_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n325_), .B1(new_n332_), .B2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n333_), .A2(new_n329_), .A3(new_n323_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n305_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n332_), .A2(new_n335_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n325_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n305_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n337_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n342_), .A2(KEYINPUT95), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT95), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n347_), .B1(new_n336_), .B2(new_n344_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  XOR2_X1   g148(.A(G8gat), .B(G36gat), .Z(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G64gat), .B(G92gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n354_), .B(KEYINPUT97), .Z(new_n355_));
  INV_X1    g154(.A(KEYINPUT94), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G226gat), .A2(G233gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT19), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G183gat), .A2(G190gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT23), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n360_), .B1(G183gat), .B2(G190gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G169gat), .A2(G176gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT22), .B(G169gat), .ZN(new_n363_));
  INV_X1    g162(.A(G176gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n361_), .A2(new_n362_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n362_), .A2(KEYINPUT24), .ZN(new_n367_));
  NOR2_X1   g166(.A1(G169gat), .A2(G176gat), .ZN(new_n368_));
  MUX2_X1   g167(.A(new_n367_), .B(KEYINPUT24), .S(new_n368_), .Z(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT26), .B(G190gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT25), .B(G183gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n369_), .A2(new_n360_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n366_), .A2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT20), .B1(new_n265_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT78), .ZN(new_n376_));
  AND3_X1   g175(.A1(new_n365_), .A2(new_n376_), .A3(new_n362_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n376_), .B1(new_n365_), .B2(new_n362_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n361_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT77), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n370_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(G190gat), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n380_), .B1(new_n382_), .B2(KEYINPUT26), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n371_), .A2(new_n383_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n369_), .B(new_n360_), .C1(new_n381_), .C2(new_n384_), .ZN(new_n385_));
  AOI22_X1  g184(.A1(new_n379_), .A2(new_n385_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n358_), .B1(new_n375_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT20), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n388_), .B1(new_n265_), .B2(new_n374_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n358_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n379_), .A2(new_n385_), .A3(new_n257_), .A4(new_n258_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n389_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n356_), .B1(new_n387_), .B2(new_n392_), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n392_), .A2(new_n356_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n355_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT27), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n375_), .A2(new_n386_), .A3(new_n358_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n390_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n354_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n396_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n389_), .A2(new_n391_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n358_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n374_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n388_), .B1(new_n404_), .B2(new_n259_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n386_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(new_n406_), .A3(new_n390_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n403_), .A2(new_n407_), .A3(new_n400_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n354_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n395_), .A2(new_n401_), .B1(new_n410_), .B2(new_n396_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n301_), .A2(new_n339_), .A3(new_n349_), .A4(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT98), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n343_), .B1(new_n342_), .B2(new_n337_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n414_), .B1(new_n348_), .B2(new_n346_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT98), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n415_), .A2(new_n416_), .A3(new_n301_), .A4(new_n411_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n413_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n301_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n342_), .A2(KEYINPUT33), .A3(new_n345_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT33), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n421_), .B1(new_n336_), .B2(new_n344_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n420_), .A2(new_n422_), .A3(new_n408_), .A4(new_n409_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n322_), .A2(new_n323_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n424_), .B1(new_n332_), .B2(new_n335_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT93), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n333_), .A2(new_n329_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n343_), .B1(new_n428_), .B2(new_n324_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n429_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n423_), .A2(new_n431_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n400_), .A2(KEYINPUT32), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n399_), .A2(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n393_), .A2(new_n394_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n434_), .B1(new_n433_), .B2(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n436_), .B1(new_n349_), .B2(new_n339_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n419_), .B1(new_n432_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT96), .ZN(new_n439_));
  OAI22_X1  g238(.A1(new_n415_), .A2(new_n436_), .B1(new_n423_), .B2(new_n431_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT96), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(new_n441_), .A3(new_n419_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n418_), .A2(new_n439_), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n379_), .A2(new_n385_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT30), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT79), .B(G43gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G227gat), .A2(G233gat), .ZN(new_n448_));
  INV_X1    g247(.A(G15gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(G71gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n447_), .A2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n320_), .B(KEYINPUT31), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(G99gat), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n445_), .A2(new_n446_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n445_), .A2(new_n446_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n451_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n452_), .A2(new_n454_), .A3(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n454_), .B1(new_n452_), .B2(new_n458_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n292_), .A2(new_n293_), .A3(new_n295_), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n298_), .A2(new_n299_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n464_), .A2(new_n288_), .A3(new_n411_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT99), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n459_), .A2(new_n460_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT99), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n464_), .A2(new_n468_), .A3(new_n288_), .A4(new_n411_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n466_), .A2(new_n467_), .A3(new_n415_), .A4(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT100), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n461_), .B1(KEYINPUT99), .B2(new_n465_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n473_), .A2(KEYINPUT100), .A3(new_n415_), .A4(new_n469_), .ZN(new_n474_));
  AOI22_X1  g273(.A1(new_n443_), .A2(new_n461_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G99gat), .A2(G106gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT6), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT6), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n479_), .A2(G99gat), .A3(G106gat), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT65), .ZN(new_n482_));
  INV_X1    g281(.A(G85gat), .ZN(new_n483_));
  INV_X1    g282(.A(G92gat), .ZN(new_n484_));
  NOR3_X1   g283(.A1(new_n483_), .A2(new_n484_), .A3(KEYINPUT9), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G85gat), .B(G92gat), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n485_), .B1(new_n487_), .B2(KEYINPUT9), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT10), .B(G99gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT64), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n482_), .B(new_n488_), .C1(G106gat), .C2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT8), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n478_), .A2(new_n480_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT66), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n493_), .A2(new_n494_), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT67), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n481_), .A2(KEYINPUT66), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT67), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n499_), .A2(new_n495_), .A3(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(G99gat), .A2(G106gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT7), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n498_), .A2(new_n501_), .A3(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n492_), .B1(new_n504_), .B2(new_n487_), .ZN(new_n505_));
  AOI211_X1 g304(.A(KEYINPUT8), .B(new_n486_), .C1(new_n482_), .C2(new_n503_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n491_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT68), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  OAI211_X1 g308(.A(KEYINPUT68), .B(new_n491_), .C1(new_n505_), .C2(new_n506_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G57gat), .B(G64gat), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n511_), .A2(KEYINPUT11), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(KEYINPUT11), .ZN(new_n513_));
  XOR2_X1   g312(.A(G71gat), .B(G78gat), .Z(new_n514_));
  NAND3_X1  g313(.A1(new_n512_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n513_), .A2(new_n514_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n509_), .A2(KEYINPUT12), .A3(new_n510_), .A4(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G230gat), .A2(G233gat), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n491_), .B(new_n517_), .C1(new_n505_), .C2(new_n506_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT12), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n507_), .A2(new_n518_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n519_), .A2(new_n520_), .A3(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n521_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n520_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(G120gat), .B(G148gat), .Z(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G176gat), .B(G204gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n525_), .A2(new_n528_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n533_), .B1(new_n525_), .B2(new_n528_), .ZN(new_n536_));
  NOR3_X1   g335(.A1(new_n535_), .A2(KEYINPUT70), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT70), .ZN(new_n538_));
  AOI211_X1 g337(.A(new_n538_), .B(new_n533_), .C1(new_n525_), .C2(new_n528_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n476_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n536_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n541_), .A2(new_n538_), .A3(new_n534_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n539_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT71), .B(KEYINPUT13), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n540_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT76), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G113gat), .B(G141gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G169gat), .B(G197gat), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n548_), .B(new_n549_), .Z(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G229gat), .A2(G233gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G15gat), .B(G22gat), .ZN(new_n553_));
  INV_X1    g352(.A(G1gat), .ZN(new_n554_));
  INV_X1    g353(.A(G8gat), .ZN(new_n555_));
  OAI21_X1  g354(.A(KEYINPUT14), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n553_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G1gat), .B(G8gat), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n557_), .B(new_n558_), .Z(new_n559_));
  XNOR2_X1  g358(.A(G29gat), .B(G36gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G43gat), .B(G50gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n559_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT75), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n563_), .A2(KEYINPUT74), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n564_), .B1(new_n563_), .B2(KEYINPUT74), .ZN(new_n567_));
  OAI22_X1  g366(.A1(new_n566_), .A2(new_n567_), .B1(new_n562_), .B2(new_n559_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n563_), .A2(KEYINPUT74), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT75), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n559_), .A2(new_n562_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n570_), .A2(new_n571_), .A3(new_n565_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n552_), .B1(new_n568_), .B2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n562_), .B(KEYINPUT15), .ZN(new_n574_));
  INV_X1    g373(.A(new_n559_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n576_), .A2(new_n552_), .A3(new_n563_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n551_), .B1(new_n573_), .B2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NOR3_X1   g379(.A1(new_n573_), .A2(new_n578_), .A3(new_n551_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n547_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  OR3_X1    g381(.A1(new_n573_), .A2(new_n578_), .A3(new_n551_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n583_), .A2(KEYINPUT76), .A3(new_n579_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n546_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G190gat), .B(G218gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G134gat), .B(G162gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n589_), .B(KEYINPUT36), .Z(new_n590_));
  OAI211_X1 g389(.A(new_n562_), .B(new_n491_), .C1(new_n505_), .C2(new_n506_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT35), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G232gat), .A2(G233gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT34), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n592_), .B1(new_n593_), .B2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n593_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n509_), .A2(new_n574_), .A3(new_n510_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n597_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n599_), .B1(new_n597_), .B2(new_n600_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n590_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n603_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n589_), .A2(KEYINPUT36), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n605_), .A2(new_n606_), .A3(new_n601_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(KEYINPUT72), .B(KEYINPUT37), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n604_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n608_), .B1(new_n604_), .B2(new_n607_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n559_), .B(new_n517_), .Z(new_n612_));
  NAND2_X1  g411(.A1(G231gat), .A2(G233gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(G127gat), .B(G155gat), .Z(new_n615_));
  XNOR2_X1  g414(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G183gat), .B(G211gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT17), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n614_), .A2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n619_), .B(KEYINPUT17), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n623_), .B1(new_n614_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n611_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n475_), .A2(new_n586_), .A3(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n415_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(new_n554_), .A3(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT38), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT101), .ZN(new_n633_));
  AND3_X1   g432(.A1(new_n604_), .A2(new_n607_), .A3(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n633_), .B1(new_n604_), .B2(new_n607_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NOR4_X1   g435(.A1(new_n475_), .A2(new_n636_), .A3(new_n626_), .A4(new_n586_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n637_), .A2(new_n630_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n632_), .B1(new_n554_), .B2(new_n638_), .ZN(G1324gat));
  INV_X1    g438(.A(new_n411_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n555_), .B1(new_n637_), .B2(new_n640_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT39), .Z(new_n642_));
  NAND3_X1  g441(.A1(new_n629_), .A2(new_n555_), .A3(new_n640_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT40), .Z(G1325gat));
  AOI21_X1  g444(.A(new_n449_), .B1(new_n637_), .B2(new_n467_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT41), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n629_), .A2(new_n449_), .A3(new_n467_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(G1326gat));
  INV_X1    g448(.A(G22gat), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n650_), .B1(new_n637_), .B2(new_n301_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT42), .Z(new_n652_));
  NAND3_X1  g451(.A1(new_n629_), .A2(new_n650_), .A3(new_n301_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1327gat));
  NOR3_X1   g453(.A1(new_n634_), .A2(new_n635_), .A3(new_n625_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n655_), .A2(new_n546_), .A3(new_n585_), .ZN(new_n656_));
  OAI21_X1  g455(.A(KEYINPUT102), .B1(new_n475_), .B2(new_n656_), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n655_), .A2(new_n546_), .A3(new_n585_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n441_), .B1(new_n440_), .B2(new_n419_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n413_), .A2(new_n417_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n467_), .B1(new_n662_), .B2(new_n442_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n470_), .B(KEYINPUT100), .ZN(new_n664_));
  OAI211_X1 g463(.A(new_n658_), .B(new_n659_), .C1(new_n663_), .C2(new_n664_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n657_), .A2(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(G29gat), .B1(new_n666_), .B2(new_n630_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n611_), .ZN(new_n668_));
  OAI21_X1  g467(.A(KEYINPUT43), .B1(new_n475_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT43), .ZN(new_n670_));
  OAI211_X1 g469(.A(new_n670_), .B(new_n611_), .C1(new_n663_), .C2(new_n664_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n546_), .A2(new_n626_), .A3(new_n585_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(KEYINPUT44), .B1(new_n672_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n676_));
  AOI211_X1 g475(.A(new_n676_), .B(new_n673_), .C1(new_n669_), .C2(new_n671_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n630_), .A2(G29gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n667_), .B1(new_n678_), .B2(new_n679_), .ZN(G1328gat));
  INV_X1    g479(.A(KEYINPUT105), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n411_), .A2(G36gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n657_), .A2(new_n665_), .A3(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT103), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT103), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n657_), .A2(new_n665_), .A3(new_n685_), .A4(new_n682_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n684_), .A2(KEYINPUT45), .A3(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n684_), .A2(new_n686_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT45), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n675_), .A2(new_n677_), .A3(new_n411_), .ZN(new_n691_));
  INV_X1    g490(.A(G36gat), .ZN(new_n692_));
  OAI211_X1 g491(.A(new_n687_), .B(new_n690_), .C1(new_n691_), .C2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT46), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n681_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n672_), .A2(new_n674_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(new_n676_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n672_), .A2(KEYINPUT44), .A3(new_n674_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n697_), .A2(new_n640_), .A3(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(G36gat), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n700_), .A2(new_n701_), .A3(new_n687_), .A4(new_n690_), .ZN(new_n702_));
  AOI21_X1  g501(.A(KEYINPUT46), .B1(new_n693_), .B2(KEYINPUT104), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n695_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n692_), .B1(new_n678_), .B2(new_n640_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n690_), .A2(new_n687_), .ZN(new_n706_));
  OAI21_X1  g505(.A(KEYINPUT104), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  AND4_X1   g506(.A1(KEYINPUT105), .A2(new_n707_), .A3(new_n694_), .A4(new_n702_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n704_), .A2(new_n708_), .ZN(G1329gat));
  NAND3_X1  g508(.A1(new_n678_), .A2(G43gat), .A3(new_n467_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n666_), .A2(new_n467_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n710_), .B1(G43gat), .B2(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g512(.A(G50gat), .B1(new_n666_), .B2(new_n301_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n301_), .A2(G50gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n678_), .B2(new_n715_), .ZN(G1331gat));
  NOR2_X1   g515(.A1(new_n475_), .A2(new_n636_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n585_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n546_), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n717_), .A2(new_n625_), .A3(new_n718_), .A4(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(G57gat), .B1(new_n720_), .B2(new_n415_), .ZN(new_n721_));
  NOR4_X1   g520(.A1(new_n475_), .A2(new_n585_), .A3(new_n628_), .A4(new_n546_), .ZN(new_n722_));
  INV_X1    g521(.A(G57gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n722_), .A2(new_n723_), .A3(new_n630_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n721_), .A2(new_n724_), .ZN(G1332gat));
  OAI21_X1  g524(.A(G64gat), .B1(new_n720_), .B2(new_n411_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT48), .ZN(new_n727_));
  INV_X1    g526(.A(G64gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n722_), .A2(new_n728_), .A3(new_n640_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(G1333gat));
  OAI21_X1  g529(.A(G71gat), .B1(new_n720_), .B2(new_n461_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(KEYINPUT106), .B(KEYINPUT49), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n731_), .B(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(G71gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n722_), .A2(new_n734_), .A3(new_n467_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(G1334gat));
  OAI21_X1  g535(.A(G78gat), .B1(new_n720_), .B2(new_n419_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT50), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n419_), .A2(G78gat), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT107), .Z(new_n740_));
  NAND2_X1  g539(.A1(new_n722_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n738_), .A2(new_n741_), .ZN(G1335gat));
  NOR2_X1   g541(.A1(new_n475_), .A2(new_n585_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n636_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n744_), .A2(new_n546_), .A3(new_n625_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n747_), .A2(new_n483_), .A3(new_n630_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n546_), .A2(new_n625_), .A3(new_n585_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT108), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n750_), .B1(new_n669_), .B2(new_n671_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT109), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n752_), .A2(new_n630_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n748_), .B1(new_n753_), .B2(new_n483_), .ZN(G1336gat));
  NAND3_X1  g553(.A1(new_n747_), .A2(new_n484_), .A3(new_n640_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n752_), .A2(new_n640_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(new_n484_), .ZN(G1337gat));
  AND2_X1   g556(.A1(new_n751_), .A2(new_n467_), .ZN(new_n758_));
  INV_X1    g557(.A(G99gat), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n461_), .A2(new_n490_), .ZN(new_n760_));
  OAI22_X1  g559(.A1(new_n758_), .A2(new_n759_), .B1(new_n746_), .B2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(KEYINPUT110), .A2(KEYINPUT51), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n761_), .B(new_n762_), .Z(G1338gat));
  NOR3_X1   g562(.A1(new_n746_), .A2(G106gat), .A3(new_n419_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765_));
  OAI21_X1  g564(.A(G106gat), .B1(new_n765_), .B2(KEYINPUT111), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n751_), .B2(new_n301_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n765_), .A2(KEYINPUT111), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n768_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n764_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n772_));
  XOR2_X1   g571(.A(new_n771_), .B(new_n772_), .Z(G1339gat));
  INV_X1    g572(.A(new_n552_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n774_), .B1(new_n568_), .B2(new_n572_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n576_), .A2(new_n774_), .A3(new_n563_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n551_), .ZN(new_n777_));
  OR3_X1    g576(.A1(new_n775_), .A2(KEYINPUT119), .A3(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT119), .B1(new_n775_), .B2(new_n777_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n778_), .A2(new_n583_), .A3(new_n779_), .ZN(new_n780_));
  XOR2_X1   g579(.A(new_n780_), .B(KEYINPUT120), .Z(new_n781_));
  NAND2_X1  g580(.A1(new_n542_), .A2(new_n543_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n784_));
  OR2_X1    g583(.A1(new_n525_), .A2(new_n784_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT117), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n525_), .A2(new_n784_), .ZN(new_n787_));
  AOI211_X1 g586(.A(KEYINPUT116), .B(new_n520_), .C1(new_n519_), .C2(new_n524_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT116), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n519_), .A2(new_n524_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n790_), .B2(new_n527_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n787_), .B1(new_n788_), .B2(new_n791_), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n786_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT56), .ZN(new_n794_));
  INV_X1    g593(.A(new_n533_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n793_), .A2(KEYINPUT118), .A3(new_n794_), .A4(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n585_), .A2(new_n534_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n795_), .B1(new_n786_), .B2(new_n792_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n794_), .A2(KEYINPUT118), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n797_), .B1(new_n798_), .B2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n783_), .B1(new_n796_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n803_), .A2(KEYINPUT57), .A3(new_n744_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n793_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n798_), .A2(KEYINPUT56), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n781_), .A2(new_n535_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n805_), .A2(new_n806_), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT58), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n805_), .A2(new_n806_), .A3(KEYINPUT58), .A4(new_n807_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n810_), .A2(new_n611_), .A3(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n802_), .B2(new_n636_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n804_), .A2(new_n812_), .A3(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n626_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n817_));
  OAI21_X1  g616(.A(KEYINPUT113), .B1(new_n585_), .B2(new_n626_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n582_), .A2(new_n819_), .A3(new_n584_), .A4(new_n625_), .ZN(new_n820_));
  AOI22_X1  g619(.A1(new_n818_), .A2(new_n820_), .B1(KEYINPUT114), .B2(KEYINPUT54), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n821_), .A2(new_n668_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n817_), .B1(new_n822_), .B2(new_n546_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n668_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n824_), .A2(KEYINPUT115), .A3(new_n719_), .ZN(new_n825_));
  OAI22_X1  g624(.A1(new_n823_), .A2(new_n825_), .B1(KEYINPUT114), .B2(KEYINPUT54), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n822_), .A2(new_n817_), .A3(new_n546_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(KEYINPUT114), .A2(KEYINPUT54), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT115), .B1(new_n824_), .B2(new_n719_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n827_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n826_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n816_), .A2(new_n832_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n473_), .A2(new_n469_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n630_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n833_), .A2(KEYINPUT59), .A3(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT59), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n831_), .B1(new_n815_), .B2(new_n626_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n839_), .B2(new_n835_), .ZN(new_n840_));
  AND2_X1   g639(.A1(new_n837_), .A2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(G113gat), .B1(new_n841_), .B2(new_n718_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n839_), .A2(new_n835_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n843_), .A2(new_n313_), .A3(new_n585_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n844_), .ZN(G1340gat));
  OAI21_X1  g644(.A(new_n311_), .B1(new_n546_), .B2(KEYINPUT60), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n843_), .B(new_n846_), .C1(KEYINPUT60), .C2(new_n311_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n546_), .B1(new_n837_), .B2(new_n840_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n847_), .B1(new_n848_), .B2(new_n311_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT121), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  OAI211_X1 g650(.A(KEYINPUT121), .B(new_n847_), .C1(new_n848_), .C2(new_n311_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1341gat));
  OAI21_X1  g652(.A(G127gat), .B1(new_n841_), .B2(new_n626_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n843_), .A2(new_n308_), .A3(new_n625_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(G1342gat));
  OAI21_X1  g655(.A(G134gat), .B1(new_n841_), .B2(new_n668_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n843_), .A2(new_n306_), .A3(new_n636_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(G1343gat));
  NAND3_X1  g658(.A1(new_n461_), .A2(new_n630_), .A3(new_n411_), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n839_), .A2(new_n419_), .A3(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n585_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n719_), .ZN(new_n864_));
  XOR2_X1   g663(.A(KEYINPUT122), .B(G148gat), .Z(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1345gat));
  NAND2_X1  g665(.A1(new_n861_), .A2(new_n625_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT61), .B(G155gat), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(G1346gat));
  AOI21_X1  g668(.A(G162gat), .B1(new_n861_), .B2(new_n636_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n611_), .A2(G162gat), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(KEYINPUT123), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n870_), .B1(new_n861_), .B2(new_n872_), .ZN(G1347gat));
  NOR4_X1   g672(.A1(new_n630_), .A2(new_n461_), .A3(new_n301_), .A4(new_n411_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n833_), .A2(new_n585_), .A3(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n875_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n833_), .A2(new_n363_), .A3(new_n585_), .A4(new_n874_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(KEYINPUT62), .B1(new_n875_), .B2(G169gat), .ZN(new_n879_));
  OAI21_X1  g678(.A(KEYINPUT124), .B1(new_n878_), .B2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n879_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT124), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n881_), .A2(new_n882_), .A3(new_n877_), .A4(new_n876_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n880_), .A2(new_n883_), .ZN(G1348gat));
  NAND2_X1  g683(.A1(new_n833_), .A2(new_n874_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n546_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(new_n364_), .ZN(G1349gat));
  NOR2_X1   g686(.A1(new_n885_), .A2(new_n626_), .ZN(new_n888_));
  MUX2_X1   g687(.A(G183gat), .B(new_n371_), .S(new_n888_), .Z(G1350gat));
  OAI21_X1  g688(.A(G190gat), .B1(new_n885_), .B2(new_n668_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n636_), .A2(new_n370_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n885_), .B2(new_n891_), .ZN(G1351gat));
  NAND4_X1  g691(.A1(new_n461_), .A2(new_n415_), .A3(new_n301_), .A4(new_n640_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n839_), .A2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n585_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n719_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g697(.A1(new_n894_), .A2(new_n625_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(KEYINPUT63), .B(G211gat), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT63), .ZN(new_n902_));
  INV_X1    g701(.A(G211gat), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n899_), .A2(new_n902_), .A3(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT125), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n899_), .A2(KEYINPUT125), .A3(new_n902_), .A4(new_n903_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n901_), .B1(new_n906_), .B2(new_n907_), .ZN(G1354gat));
  NAND2_X1  g707(.A1(new_n894_), .A2(new_n636_), .ZN(new_n909_));
  XOR2_X1   g708(.A(KEYINPUT126), .B(G218gat), .Z(new_n910_));
  NOR2_X1   g709(.A1(new_n668_), .A2(new_n910_), .ZN(new_n911_));
  AOI22_X1  g710(.A1(new_n909_), .A2(new_n910_), .B1(new_n894_), .B2(new_n911_), .ZN(G1355gat));
endmodule


