//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 1 0 0 1 1 1 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n805_, new_n806_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n937_, new_n939_, new_n940_, new_n942_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n966_, new_n967_, new_n969_, new_n970_, new_n972_, new_n973_,
    new_n974_, new_n976_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n983_, new_n984_;
  XNOR2_X1  g000(.A(G22gat), .B(G50gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(G155gat), .ZN(new_n204_));
  INV_X1    g003(.A(G162gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n204_), .A2(new_n205_), .A3(KEYINPUT84), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT84), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n207_), .B1(G155gat), .B2(G162gat), .ZN(new_n208_));
  AOI22_X1  g007(.A1(new_n206_), .A2(new_n208_), .B1(G155gat), .B2(G162gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n210_));
  INV_X1    g009(.A(G141gat), .ZN(new_n211_));
  INV_X1    g010(.A(G148gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT85), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G141gat), .A2(G148gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT85), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(new_n216_), .A3(new_n210_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n214_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G141gat), .A2(G148gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT2), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n221_), .B(new_n222_), .C1(new_n210_), .C2(new_n215_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n209_), .B1(new_n218_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n206_), .A2(new_n208_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT1), .B1(new_n204_), .B2(new_n205_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT1), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(G155gat), .A3(G162gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n225_), .A2(new_n226_), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n211_), .A2(new_n212_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n230_), .A2(new_n219_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n224_), .A2(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n233_), .A2(KEYINPUT29), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT28), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  AOI22_X1  g035(.A1(new_n230_), .A2(KEYINPUT3), .B1(new_n220_), .B2(new_n219_), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n237_), .A2(new_n214_), .A3(new_n222_), .A4(new_n217_), .ZN(new_n238_));
  AOI22_X1  g037(.A1(new_n238_), .A2(new_n209_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT29), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n241_), .A2(KEYINPUT28), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n203_), .B1(new_n236_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n234_), .A2(new_n235_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n241_), .A2(KEYINPUT28), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(new_n245_), .A3(new_n202_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n240_), .B1(new_n224_), .B2(new_n232_), .ZN(new_n248_));
  INV_X1    g047(.A(G197gat), .ZN(new_n249_));
  INV_X1    g048(.A(G204gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G197gat), .A2(G204gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT21), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n251_), .A2(KEYINPUT21), .A3(new_n252_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G211gat), .B(G218gat), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n256_), .A2(new_n257_), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT86), .B1(new_n248_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT86), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n258_), .A2(new_n259_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n262_), .B(new_n263_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n261_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G228gat), .A2(G233gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n266_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n261_), .A2(new_n268_), .A3(new_n264_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G78gat), .B(G106gat), .ZN(new_n271_));
  XOR2_X1   g070(.A(new_n271_), .B(KEYINPUT87), .Z(new_n272_));
  AOI21_X1  g071(.A(new_n247_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT88), .ZN(new_n274_));
  AND3_X1   g073(.A1(new_n261_), .A2(new_n268_), .A3(new_n264_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n268_), .B1(new_n261_), .B2(new_n264_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n274_), .B1(new_n277_), .B2(new_n271_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n271_), .ZN(new_n279_));
  NOR4_X1   g078(.A1(new_n275_), .A2(new_n276_), .A3(KEYINPUT88), .A4(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n273_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n272_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n272_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n267_), .A2(new_n283_), .A3(new_n269_), .ZN(new_n284_));
  AOI22_X1  g083(.A1(new_n282_), .A2(new_n284_), .B1(new_n246_), .B2(new_n243_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n281_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(G134gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(G127gat), .ZN(new_n289_));
  INV_X1    g088(.A(G127gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(G134gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(G120gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(G113gat), .ZN(new_n294_));
  INV_X1    g093(.A(G113gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G120gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n292_), .A2(new_n297_), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n289_), .A2(new_n291_), .A3(new_n294_), .A4(new_n296_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n224_), .A2(new_n300_), .A3(new_n232_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT83), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n302_), .B1(new_n292_), .B2(new_n297_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  OAI211_X1 g105(.A(KEYINPUT4), .B(new_n301_), .C1(new_n306_), .C2(new_n239_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G225gat), .A2(G233gat), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(KEYINPUT83), .B1(new_n298_), .B2(new_n299_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n310_), .A2(new_n304_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT4), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n233_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n307_), .A2(new_n309_), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n233_), .A2(new_n311_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n315_), .A2(new_n301_), .A3(new_n308_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G1gat), .B(G29gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(G85gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT0), .B(G57gat), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n319_), .B(new_n320_), .Z(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n317_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n314_), .A2(new_n316_), .A3(new_n321_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(G8gat), .B(G36gat), .Z(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT18), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G64gat), .B(G92gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT20), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT79), .ZN(new_n333_));
  INV_X1    g132(.A(G190gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(KEYINPUT79), .A2(G190gat), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(KEYINPUT26), .A3(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT80), .ZN(new_n338_));
  INV_X1    g137(.A(G183gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT25), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT25), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(G183gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT26), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(G190gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n340_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT80), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n335_), .A2(new_n347_), .A3(KEYINPUT26), .A4(new_n336_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n338_), .A2(new_n346_), .A3(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(G169gat), .ZN(new_n354_));
  INV_X1    g153(.A(G176gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G169gat), .A2(G176gat), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n356_), .A2(KEYINPUT24), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT24), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n359_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n353_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n354_), .A2(KEYINPUT22), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT22), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(G169gat), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n362_), .A2(new_n364_), .A3(new_n355_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT22), .B(G169gat), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n368_), .A2(KEYINPUT81), .A3(new_n355_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n357_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n335_), .A2(new_n339_), .A3(new_n336_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n371_), .B1(new_n353_), .B2(new_n372_), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n349_), .A2(new_n361_), .B1(new_n370_), .B2(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n332_), .B1(new_n374_), .B2(new_n260_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n334_), .A2(KEYINPUT26), .ZN(new_n376_));
  NAND4_X1  g175(.A1(new_n340_), .A2(new_n342_), .A3(new_n344_), .A4(new_n376_), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n377_), .A2(KEYINPUT91), .A3(new_n358_), .ZN(new_n378_));
  AOI21_X1  g177(.A(KEYINPUT91), .B1(new_n377_), .B2(new_n358_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n353_), .A2(new_n360_), .ZN(new_n380_));
  NOR3_X1   g179(.A1(new_n378_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n353_), .B1(G183gat), .B2(G190gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n357_), .B(KEYINPUT92), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(new_n365_), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n263_), .B1(new_n381_), .B2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT90), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n375_), .A2(new_n386_), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n349_), .A2(new_n361_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n370_), .A2(new_n373_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n332_), .B1(new_n394_), .B2(new_n263_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n377_), .A2(new_n358_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT91), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n377_), .A2(KEYINPUT91), .A3(new_n358_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n380_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n398_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n401_), .A2(new_n260_), .A3(new_n384_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n389_), .B1(new_n395_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT95), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n391_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  AOI211_X1 g204(.A(KEYINPUT95), .B(new_n389_), .C1(new_n395_), .C2(new_n402_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n331_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n390_), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT20), .B1(new_n394_), .B2(new_n263_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n260_), .B1(new_n401_), .B2(new_n384_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n408_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n395_), .A2(new_n389_), .A3(new_n402_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(new_n330_), .A3(new_n412_), .ZN(new_n413_));
  AND2_X1   g212(.A1(new_n413_), .A2(KEYINPUT27), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n370_), .A2(new_n373_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n353_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n345_), .B1(KEYINPUT80), .B2(new_n337_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n416_), .B1(new_n417_), .B2(new_n348_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n263_), .B1(new_n415_), .B2(new_n418_), .ZN(new_n419_));
  AND4_X1   g218(.A1(KEYINPUT20), .A2(new_n419_), .A3(new_n402_), .A4(new_n389_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n390_), .B1(new_n375_), .B2(new_n386_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n331_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n413_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT27), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n407_), .A2(new_n414_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n287_), .A2(new_n326_), .A3(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n330_), .A2(KEYINPUT32), .ZN(new_n427_));
  INV_X1    g226(.A(new_n389_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n402_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT20), .B1(new_n374_), .B2(new_n260_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n428_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n409_), .A2(new_n410_), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n431_), .A2(KEYINPUT95), .B1(new_n432_), .B2(new_n390_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n406_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n427_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n324_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n321_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n427_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n411_), .A2(new_n412_), .ZN(new_n439_));
  OAI22_X1  g238(.A1(new_n436_), .A2(new_n437_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n435_), .A2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n436_), .A2(KEYINPUT94), .A3(KEYINPUT33), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT94), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT33), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n443_), .B1(new_n324_), .B2(new_n444_), .ZN(new_n445_));
  AND3_X1   g244(.A1(new_n307_), .A2(new_n308_), .A3(new_n313_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n315_), .A2(new_n301_), .A3(new_n309_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n322_), .A2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT33), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(new_n324_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n442_), .A2(new_n445_), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT93), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n453_), .B1(new_n422_), .B2(new_n413_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n422_), .A2(new_n453_), .A3(new_n413_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n441_), .B1(new_n452_), .B2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n426_), .B1(new_n458_), .B2(new_n287_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT31), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n460_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n461_));
  NOR3_X1   g260(.A1(new_n310_), .A2(KEYINPUT31), .A3(new_n304_), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT82), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G227gat), .A2(G233gat), .ZN(new_n464_));
  INV_X1    g263(.A(G15gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT30), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n374_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n467_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n394_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n463_), .A2(new_n468_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT82), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n303_), .A2(new_n460_), .A3(new_n305_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT31), .B1(new_n310_), .B2(new_n304_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n472_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n394_), .A2(new_n469_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n374_), .A2(new_n467_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n475_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G71gat), .B(G99gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(G43gat), .ZN(new_n480_));
  AND3_X1   g279(.A1(new_n471_), .A2(new_n478_), .A3(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n480_), .B1(new_n471_), .B2(new_n478_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n483_), .A2(new_n325_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n425_), .A2(new_n281_), .A3(new_n286_), .A4(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT96), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT88), .B1(new_n270_), .B2(new_n279_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n277_), .A2(new_n274_), .A3(new_n271_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n285_), .B1(new_n490_), .B2(new_n273_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n491_), .A2(KEYINPUT96), .A3(new_n425_), .A4(new_n484_), .ZN(new_n492_));
  AOI22_X1  g291(.A1(new_n459_), .A2(new_n483_), .B1(new_n487_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G229gat), .A2(G233gat), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(G29gat), .B(G36gat), .Z(new_n496_));
  INV_X1    g295(.A(KEYINPUT67), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G29gat), .B(G36gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n499_), .A2(KEYINPUT67), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT68), .B1(new_n498_), .B2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G43gat), .B(G50gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n496_), .A2(new_n497_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT68), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n499_), .A2(KEYINPUT67), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  AND3_X1   g305(.A1(new_n501_), .A2(new_n502_), .A3(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n502_), .B1(new_n501_), .B2(new_n506_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT73), .B(G8gat), .ZN(new_n510_));
  INV_X1    g309(.A(G1gat), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT14), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G15gat), .B(G22gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT74), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G1gat), .B(G8gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT74), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n514_), .B(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n516_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n509_), .A2(new_n517_), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n509_), .B1(new_n517_), .B2(new_n521_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n495_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n517_), .A2(new_n521_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n502_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n506_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n504_), .B1(new_n503_), .B2(new_n505_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n527_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n501_), .A2(new_n502_), .A3(new_n506_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n526_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT15), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n534_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n530_), .A2(KEYINPUT15), .A3(new_n531_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n535_), .A2(new_n536_), .A3(new_n517_), .A4(new_n521_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n533_), .A2(new_n537_), .A3(new_n494_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G113gat), .B(G141gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G169gat), .B(G197gat), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n539_), .B(new_n540_), .Z(new_n541_));
  NAND3_X1  g340(.A1(new_n525_), .A2(new_n538_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n541_), .B1(new_n525_), .B2(new_n538_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(G230gat), .ZN(new_n546_));
  INV_X1    g345(.A(G233gat), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G57gat), .B(G64gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G71gat), .B(G78gat), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(new_n550_), .A3(KEYINPUT11), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(KEYINPUT11), .ZN(new_n552_));
  INV_X1    g351(.A(new_n550_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n549_), .A2(KEYINPUT11), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n551_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G99gat), .A2(G106gat), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT6), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  OR2_X1    g360(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n562_));
  INV_X1    g361(.A(G106gat), .ZN(new_n563_));
  NAND2_X1  g362(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n562_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G85gat), .A2(G92gat), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n566_), .A2(KEYINPUT9), .ZN(new_n567_));
  INV_X1    g366(.A(G85gat), .ZN(new_n568_));
  INV_X1    g367(.A(G92gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(KEYINPUT9), .A3(new_n566_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n561_), .A2(new_n565_), .A3(new_n567_), .A4(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT7), .ZN(new_n573_));
  INV_X1    g372(.A(G99gat), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n573_), .A2(new_n574_), .A3(new_n563_), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n575_), .A2(new_n559_), .A3(new_n560_), .A4(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT8), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n570_), .A2(new_n566_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n577_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n578_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n556_), .B(new_n572_), .C1(new_n581_), .C2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT64), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n572_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n556_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n548_), .B1(new_n585_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n572_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n582_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n591_), .B1(new_n592_), .B2(new_n580_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n548_), .B1(new_n593_), .B2(new_n556_), .ZN(new_n594_));
  AOI21_X1  g393(.A(KEYINPUT12), .B1(new_n588_), .B2(KEYINPUT65), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT65), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT12), .ZN(new_n597_));
  AOI211_X1 g396(.A(new_n596_), .B(new_n597_), .C1(new_n586_), .C2(new_n587_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n594_), .B1(new_n595_), .B2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n590_), .A2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G120gat), .B(G148gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT5), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G176gat), .B(G204gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT66), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n600_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT13), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n590_), .A2(new_n599_), .A3(new_n604_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n606_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n607_), .B1(new_n606_), .B2(new_n608_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n493_), .A2(new_n545_), .A3(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(G127gat), .B(G155gat), .Z(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT16), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G183gat), .B(G211gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G231gat), .A2(G233gat), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT75), .Z(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n517_), .A2(new_n521_), .A3(new_n556_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n556_), .B1(new_n517_), .B2(new_n521_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n622_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n526_), .A2(new_n587_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n627_), .A2(new_n621_), .A3(new_n623_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n619_), .B1(new_n626_), .B2(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n616_), .B(KEYINPUT17), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n626_), .A2(new_n628_), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT77), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n626_), .A2(new_n628_), .A3(KEYINPUT77), .A4(new_n630_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n629_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(G190gat), .B(G218gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT69), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G134gat), .B(G162gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT36), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n535_), .A2(new_n536_), .A3(new_n586_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT35), .ZN(new_n643_));
  NAND2_X1  g442(.A1(G232gat), .A2(G233gat), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT34), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  AOI22_X1  g445(.A1(new_n532_), .A2(new_n593_), .B1(new_n643_), .B2(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n646_), .A2(new_n643_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n642_), .A2(new_n647_), .A3(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n642_), .B2(new_n647_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n641_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n642_), .A2(new_n647_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(new_n648_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n642_), .A2(new_n647_), .A3(new_n649_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT36), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n640_), .A2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT70), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n654_), .A2(new_n655_), .A3(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n652_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n636_), .A2(new_n661_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n612_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G1gat), .B1(new_n664_), .B2(new_n326_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT38), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT78), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n652_), .A2(KEYINPUT71), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT71), .ZN(new_n669_));
  OAI211_X1 g468(.A(new_n669_), .B(new_n641_), .C1(new_n650_), .C2(new_n651_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n668_), .A2(new_n670_), .A3(new_n659_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n671_), .A2(KEYINPUT72), .A3(KEYINPUT37), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(KEYINPUT72), .B1(new_n671_), .B2(KEYINPUT37), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n660_), .A2(KEYINPUT37), .ZN(new_n675_));
  NOR3_X1   g474(.A1(new_n673_), .A2(new_n674_), .A3(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n667_), .B1(new_n676_), .B2(new_n636_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n641_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n678_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n659_), .B1(new_n679_), .B2(new_n669_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n670_), .ZN(new_n681_));
  OAI21_X1  g480(.A(KEYINPUT37), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT72), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n675_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n684_), .A2(new_n672_), .A3(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n686_), .A2(KEYINPUT78), .A3(new_n635_), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n612_), .A2(new_n677_), .A3(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n688_), .A2(new_n511_), .A3(new_n325_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT97), .ZN(new_n690_));
  AND3_X1   g489(.A1(new_n689_), .A2(new_n690_), .A3(new_n666_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n689_), .B2(new_n666_), .ZN(new_n692_));
  OAI221_X1 g491(.A(new_n665_), .B1(new_n666_), .B2(new_n689_), .C1(new_n691_), .C2(new_n692_), .ZN(G1324gat));
  INV_X1    g492(.A(new_n425_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n688_), .A2(new_n510_), .A3(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n663_), .A2(new_n694_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT39), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n696_), .A2(new_n697_), .A3(G8gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n696_), .B2(G8gat), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n695_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g500(.A(new_n483_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n465_), .B1(new_n663_), .B2(new_n702_), .ZN(new_n703_));
  XOR2_X1   g502(.A(KEYINPUT98), .B(KEYINPUT41), .Z(new_n704_));
  OR2_X1    g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n688_), .A2(new_n465_), .A3(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n703_), .A2(new_n704_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n705_), .A2(new_n706_), .A3(new_n707_), .ZN(G1326gat));
  INV_X1    g507(.A(G22gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n663_), .B2(new_n287_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT42), .Z(new_n711_));
  NAND3_X1  g510(.A1(new_n688_), .A2(new_n709_), .A3(new_n287_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1327gat));
  NOR2_X1   g512(.A1(new_n635_), .A2(new_n660_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n612_), .A2(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(G29gat), .B1(new_n715_), .B2(new_n325_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT99), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT43), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n487_), .A2(new_n492_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n438_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n721_), .B(new_n325_), .C1(new_n438_), .C2(new_n439_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n456_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n723_), .A2(new_n454_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n722_), .B1(new_n724_), .B2(new_n451_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n325_), .B1(new_n281_), .B2(new_n286_), .ZN(new_n726_));
  AOI22_X1  g525(.A1(new_n725_), .A2(new_n491_), .B1(new_n726_), .B2(new_n425_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n720_), .B1(new_n727_), .B2(new_n702_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n676_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n717_), .A2(KEYINPUT43), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n719_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n720_), .B(KEYINPUT100), .C1(new_n727_), .C2(new_n702_), .ZN(new_n732_));
  AND2_X1   g531(.A1(KEYINPUT100), .A2(KEYINPUT43), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n732_), .B(new_n676_), .C1(new_n493_), .C2(new_n733_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n611_), .A2(new_n635_), .A3(new_n545_), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n731_), .A2(KEYINPUT44), .A3(new_n734_), .A4(new_n735_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n736_), .A2(G29gat), .A3(new_n325_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n730_), .B1(new_n493_), .B2(new_n686_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n734_), .A2(new_n718_), .A3(new_n738_), .A4(new_n735_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT44), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n716_), .B1(new_n737_), .B2(new_n741_), .ZN(G1328gat));
  INV_X1    g541(.A(G36gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n715_), .A2(new_n743_), .A3(new_n694_), .ZN(new_n744_));
  XOR2_X1   g543(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n745_));
  XNOR2_X1  g544(.A(new_n744_), .B(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n741_), .A2(new_n694_), .A3(new_n736_), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n747_), .A2(KEYINPUT101), .A3(G36gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(KEYINPUT101), .B1(new_n747_), .B2(G36gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n746_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT46), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  OAI211_X1 g551(.A(KEYINPUT46), .B(new_n746_), .C1(new_n748_), .C2(new_n749_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(G1329gat));
  NAND3_X1  g553(.A1(new_n736_), .A2(G43gat), .A3(new_n702_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n741_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n715_), .A2(new_n702_), .ZN(new_n757_));
  OAI22_X1  g556(.A1(new_n755_), .A2(new_n756_), .B1(new_n757_), .B2(G43gat), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g558(.A(G50gat), .B1(new_n715_), .B2(new_n287_), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n736_), .A2(G50gat), .A3(new_n287_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(new_n741_), .ZN(G1331gat));
  NAND3_X1  g561(.A1(new_n677_), .A2(new_n687_), .A3(new_n611_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT103), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n545_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n493_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n763_), .A2(new_n764_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n765_), .A2(new_n767_), .A3(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(G57gat), .B1(new_n769_), .B2(new_n325_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT104), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  AOI211_X1 g571(.A(KEYINPUT104), .B(G57gat), .C1(new_n769_), .C2(new_n325_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n611_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n635_), .A2(new_n545_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n774_), .A2(new_n775_), .A3(new_n661_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n728_), .A2(new_n776_), .ZN(new_n777_));
  XOR2_X1   g576(.A(new_n777_), .B(KEYINPUT105), .Z(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(G57gat), .A3(new_n325_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT106), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n772_), .A2(new_n773_), .A3(new_n780_), .ZN(G1332gat));
  INV_X1    g580(.A(G64gat), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n782_), .B1(new_n778_), .B2(new_n694_), .ZN(new_n783_));
  XOR2_X1   g582(.A(new_n783_), .B(KEYINPUT48), .Z(new_n784_));
  NAND3_X1  g583(.A1(new_n769_), .A2(new_n782_), .A3(new_n694_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(G1333gat));
  INV_X1    g585(.A(G71gat), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n787_), .B1(new_n778_), .B2(new_n702_), .ZN(new_n788_));
  XOR2_X1   g587(.A(new_n788_), .B(KEYINPUT49), .Z(new_n789_));
  NAND3_X1  g588(.A1(new_n769_), .A2(new_n787_), .A3(new_n702_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(G1334gat));
  INV_X1    g590(.A(G78gat), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n792_), .B1(new_n778_), .B2(new_n287_), .ZN(new_n793_));
  XOR2_X1   g592(.A(new_n793_), .B(KEYINPUT50), .Z(new_n794_));
  NOR2_X1   g593(.A1(new_n491_), .A2(G78gat), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT107), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n769_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n794_), .A2(new_n797_), .ZN(G1335gat));
  AND3_X1   g597(.A1(new_n767_), .A2(new_n611_), .A3(new_n714_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n799_), .A2(new_n568_), .A3(new_n325_), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n774_), .A2(new_n635_), .A3(new_n766_), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n731_), .A2(new_n734_), .A3(new_n801_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n802_), .A2(new_n325_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n800_), .B1(new_n803_), .B2(new_n568_), .ZN(G1336gat));
  NAND3_X1  g603(.A1(new_n799_), .A2(new_n569_), .A3(new_n694_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n802_), .A2(new_n694_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(new_n569_), .ZN(G1337gat));
  AND3_X1   g606(.A1(new_n702_), .A2(new_n562_), .A3(new_n564_), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT108), .B1(new_n799_), .B2(new_n808_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n802_), .A2(new_n702_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(new_n574_), .ZN(new_n811_));
  XOR2_X1   g610(.A(KEYINPUT109), .B(KEYINPUT51), .Z(new_n812_));
  XNOR2_X1  g611(.A(new_n811_), .B(new_n812_), .ZN(G1338gat));
  NAND3_X1  g612(.A1(new_n799_), .A2(new_n563_), .A3(new_n287_), .ZN(new_n814_));
  XOR2_X1   g613(.A(new_n814_), .B(KEYINPUT110), .Z(new_n815_));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n731_), .A2(new_n287_), .A3(new_n734_), .A4(new_n801_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT111), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(G106gat), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n817_), .A2(new_n818_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n816_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n802_), .A2(KEYINPUT111), .A3(new_n287_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n823_), .A2(KEYINPUT52), .A3(G106gat), .A4(new_n819_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n815_), .A2(new_n822_), .A3(new_n824_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n815_), .A2(new_n822_), .A3(new_n824_), .A4(new_n826_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(G1339gat));
  AOI21_X1  g629(.A(new_n495_), .B1(new_n533_), .B2(new_n522_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n832_));
  OR3_X1    g631(.A1(new_n831_), .A2(new_n832_), .A3(new_n541_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n533_), .A2(new_n537_), .A3(new_n495_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n832_), .B1(new_n831_), .B2(new_n541_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n833_), .A2(new_n834_), .A3(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n542_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n606_), .A2(new_n608_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n608_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n594_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT65), .B1(new_n593_), .B2(new_n556_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n597_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n588_), .A2(KEYINPUT65), .A3(KEYINPUT12), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n841_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(KEYINPUT115), .B1(new_n845_), .B2(KEYINPUT55), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT115), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT55), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n599_), .A2(new_n847_), .A3(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n595_), .A2(new_n598_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n548_), .B1(new_n850_), .B2(new_n585_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n845_), .A2(KEYINPUT55), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n846_), .A2(new_n849_), .A3(new_n851_), .A4(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n605_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT56), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n853_), .A2(KEYINPUT56), .A3(new_n605_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n840_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n839_), .A2(new_n858_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n859_), .A2(KEYINPUT57), .A3(new_n660_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n660_), .B1(new_n839_), .B2(new_n858_), .ZN(new_n861_));
  XOR2_X1   g660(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT118), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n857_), .A2(new_n865_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n853_), .A2(KEYINPUT118), .A3(KEYINPUT56), .A4(new_n605_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n866_), .A2(new_n856_), .A3(new_n867_), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n836_), .A2(new_n542_), .A3(new_n608_), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n676_), .B1(new_n870_), .B2(KEYINPUT58), .ZN(new_n871_));
  AND3_X1   g670(.A1(new_n868_), .A2(new_n869_), .A3(KEYINPUT58), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n860_), .B(new_n864_), .C1(new_n871_), .C2(new_n872_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n635_), .B(new_n545_), .C1(new_n610_), .C2(new_n609_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n675_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n877_));
  AOI211_X1 g676(.A(new_n875_), .B(new_n876_), .C1(new_n877_), .C2(new_n672_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n876_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT37), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n650_), .A2(new_n651_), .ZN(new_n881_));
  AOI22_X1  g680(.A1(new_n652_), .A2(KEYINPUT71), .B1(new_n881_), .B2(new_n658_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n880_), .B1(new_n882_), .B2(new_n670_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n685_), .B1(new_n883_), .B2(KEYINPUT72), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n879_), .B1(new_n884_), .B2(new_n673_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n875_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT114), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n878_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n885_), .A2(KEYINPUT114), .A3(new_n875_), .ZN(new_n889_));
  AOI22_X1  g688(.A1(new_n873_), .A2(new_n636_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n694_), .A2(new_n287_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n326_), .A2(new_n483_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(KEYINPUT59), .B1(new_n890_), .B2(new_n893_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n545_), .A2(new_n295_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(KEYINPUT121), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n888_), .A2(new_n889_), .ZN(new_n897_));
  AOI21_X1  g696(.A(KEYINPUT58), .B1(new_n868_), .B2(new_n869_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n872_), .A2(new_n898_), .A3(new_n686_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n864_), .ZN(new_n900_));
  OAI21_X1  g699(.A(KEYINPUT120), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT120), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n902_), .B(new_n864_), .C1(new_n871_), .C2(new_n872_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n901_), .A2(new_n903_), .A3(new_n860_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n897_), .B1(new_n904_), .B2(new_n636_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n893_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n894_), .B(new_n896_), .C1(new_n905_), .C2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n890_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n910_), .A2(new_n766_), .A3(new_n906_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n295_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n909_), .A2(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(KEYINPUT122), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n909_), .A2(new_n912_), .A3(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n916_), .ZN(G1340gat));
  OAI21_X1  g716(.A(new_n894_), .B1(new_n905_), .B2(new_n908_), .ZN(new_n918_));
  OAI21_X1  g717(.A(G120gat), .B1(new_n918_), .B2(new_n774_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n910_), .A2(new_n906_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n293_), .B1(new_n774_), .B2(KEYINPUT60), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n921_), .B1(KEYINPUT60), .B2(new_n293_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n919_), .B1(new_n920_), .B2(new_n922_), .ZN(G1341gat));
  INV_X1    g722(.A(new_n918_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n635_), .A2(G127gat), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(KEYINPUT123), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n910_), .A2(new_n635_), .A3(new_n906_), .ZN(new_n927_));
  AOI22_X1  g726(.A1(new_n924_), .A2(new_n926_), .B1(new_n290_), .B2(new_n927_), .ZN(G1342gat));
  OAI21_X1  g727(.A(G134gat), .B1(new_n918_), .B2(new_n686_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n661_), .A2(new_n288_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n920_), .B2(new_n930_), .ZN(G1343gat));
  NAND4_X1  g730(.A1(new_n287_), .A2(new_n325_), .A3(new_n425_), .A4(new_n483_), .ZN(new_n932_));
  XOR2_X1   g731(.A(new_n932_), .B(KEYINPUT124), .Z(new_n933_));
  NAND2_X1  g732(.A1(new_n910_), .A2(new_n933_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n934_), .A2(new_n545_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(new_n211_), .ZN(G1344gat));
  NOR2_X1   g735(.A1(new_n934_), .A2(new_n774_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(new_n212_), .ZN(G1345gat));
  NOR2_X1   g737(.A1(new_n934_), .A2(new_n636_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(KEYINPUT61), .B(G155gat), .ZN(new_n940_));
  XOR2_X1   g739(.A(new_n939_), .B(new_n940_), .Z(G1346gat));
  OAI21_X1  g740(.A(G162gat), .B1(new_n934_), .B2(new_n686_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n661_), .A2(new_n205_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n942_), .B1(new_n934_), .B2(new_n943_), .ZN(G1347gat));
  XOR2_X1   g743(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n945_));
  INV_X1    g744(.A(new_n945_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n354_), .B1(new_n946_), .B2(KEYINPUT126), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n946_), .A2(KEYINPUT126), .ZN(new_n948_));
  INV_X1    g747(.A(new_n948_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n694_), .A2(new_n491_), .A3(new_n484_), .ZN(new_n950_));
  INV_X1    g749(.A(new_n950_), .ZN(new_n951_));
  AND2_X1   g750(.A1(new_n904_), .A2(new_n636_), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n951_), .B1(new_n952_), .B2(new_n897_), .ZN(new_n953_));
  OAI211_X1 g752(.A(new_n947_), .B(new_n949_), .C1(new_n953_), .C2(new_n545_), .ZN(new_n954_));
  NOR3_X1   g753(.A1(new_n905_), .A2(new_n545_), .A3(new_n950_), .ZN(new_n955_));
  INV_X1    g754(.A(new_n947_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n948_), .B1(new_n955_), .B2(new_n956_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n955_), .A2(new_n368_), .ZN(new_n958_));
  NAND3_X1  g757(.A1(new_n954_), .A2(new_n957_), .A3(new_n958_), .ZN(G1348gat));
  NOR2_X1   g758(.A1(new_n905_), .A2(new_n950_), .ZN(new_n960_));
  AOI21_X1  g759(.A(G176gat), .B1(new_n960_), .B2(new_n611_), .ZN(new_n961_));
  NAND4_X1  g760(.A1(new_n910_), .A2(G176gat), .A3(new_n611_), .A4(new_n951_), .ZN(new_n962_));
  OR2_X1    g761(.A1(new_n962_), .A2(KEYINPUT127), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n962_), .A2(KEYINPUT127), .ZN(new_n964_));
  AOI21_X1  g763(.A(new_n961_), .B1(new_n963_), .B2(new_n964_), .ZN(G1349gat));
  AOI21_X1  g764(.A(new_n636_), .B1(new_n340_), .B2(new_n342_), .ZN(new_n966_));
  NAND3_X1  g765(.A1(new_n910_), .A2(new_n635_), .A3(new_n951_), .ZN(new_n967_));
  AOI22_X1  g766(.A1(new_n960_), .A2(new_n966_), .B1(new_n339_), .B2(new_n967_), .ZN(G1350gat));
  OAI21_X1  g767(.A(G190gat), .B1(new_n953_), .B2(new_n686_), .ZN(new_n969_));
  NAND3_X1  g768(.A1(new_n661_), .A2(new_n344_), .A3(new_n376_), .ZN(new_n970_));
  OAI21_X1  g769(.A(new_n969_), .B1(new_n953_), .B2(new_n970_), .ZN(G1351gat));
  NOR4_X1   g770(.A1(new_n491_), .A2(new_n425_), .A3(new_n325_), .A4(new_n702_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n910_), .A2(new_n972_), .ZN(new_n973_));
  NOR2_X1   g772(.A1(new_n973_), .A2(new_n545_), .ZN(new_n974_));
  XNOR2_X1  g773(.A(new_n974_), .B(new_n249_), .ZN(G1352gat));
  NOR2_X1   g774(.A1(new_n973_), .A2(new_n774_), .ZN(new_n976_));
  XNOR2_X1  g775(.A(new_n976_), .B(new_n250_), .ZN(G1353gat));
  NAND3_X1  g776(.A1(new_n910_), .A2(new_n635_), .A3(new_n972_), .ZN(new_n978_));
  NOR2_X1   g777(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n979_));
  AND2_X1   g778(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n980_));
  NOR3_X1   g779(.A1(new_n978_), .A2(new_n979_), .A3(new_n980_), .ZN(new_n981_));
  AOI21_X1  g780(.A(new_n981_), .B1(new_n978_), .B2(new_n979_), .ZN(G1354gat));
  OAI21_X1  g781(.A(G218gat), .B1(new_n973_), .B2(new_n686_), .ZN(new_n983_));
  OR2_X1    g782(.A1(new_n660_), .A2(G218gat), .ZN(new_n984_));
  OAI21_X1  g783(.A(new_n983_), .B1(new_n973_), .B2(new_n984_), .ZN(G1355gat));
endmodule


