//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0 0 0 1 0 1 1 0 0 1 0 1 1 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 1 0 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n903_, new_n904_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n944_, new_n945_, new_n947_, new_n948_, new_n949_,
    new_n951_, new_n952_, new_n953_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n960_, new_n961_, new_n962_, new_n963_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT36), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT10), .B(G99gat), .ZN(new_n210_));
  OAI211_X1 g009(.A(new_n208_), .B(new_n209_), .C1(new_n210_), .C2(G106gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G92gat), .ZN(new_n214_));
  INV_X1    g013(.A(G85gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n213_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n211_), .B1(new_n212_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT7), .ZN(new_n218_));
  INV_X1    g017(.A(G99gat), .ZN(new_n219_));
  INV_X1    g018(.A(G106gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n221_), .A2(new_n208_), .A3(new_n209_), .A4(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(G85gat), .B(G92gat), .Z(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n226_), .A2(KEYINPUT8), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n227_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n223_), .A2(new_n229_), .A3(new_n224_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n226_), .A2(KEYINPUT8), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n217_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G29gat), .B(G36gat), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(G43gat), .B(G50gat), .Z(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G43gat), .B(G50gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n234_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n233_), .A2(new_n240_), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n223_), .A2(new_n229_), .A3(new_n224_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n229_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n232_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n216_), .A2(new_n212_), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n210_), .A2(G106gat), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n245_), .A2(new_n246_), .A3(new_n208_), .A4(new_n209_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n244_), .A2(new_n247_), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n237_), .A2(KEYINPUT15), .A3(new_n239_), .ZN(new_n249_));
  AOI21_X1  g048(.A(KEYINPUT15), .B1(new_n237_), .B2(new_n239_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n248_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G232gat), .A2(G233gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT34), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n254_), .A2(KEYINPUT35), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n241_), .A2(new_n252_), .A3(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(KEYINPUT35), .A3(new_n254_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n204_), .A2(KEYINPUT36), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n254_), .A2(KEYINPUT35), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n241_), .A2(new_n252_), .A3(new_n259_), .A4(new_n255_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n257_), .A2(new_n258_), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n258_), .B1(new_n257_), .B2(new_n260_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n205_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT37), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT69), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n265_), .B1(new_n261_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n264_), .A2(new_n268_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n267_), .B(new_n205_), .C1(new_n262_), .C2(new_n263_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT72), .B(KEYINPUT16), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G127gat), .B(G155gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G183gat), .B(G211gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT17), .ZN(new_n277_));
  AND2_X1   g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n276_), .A2(new_n277_), .ZN(new_n279_));
  OR3_X1    g078(.A1(new_n278_), .A2(new_n279_), .A3(KEYINPUT73), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n281_));
  INV_X1    g080(.A(G64gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(G57gat), .ZN(new_n283_));
  INV_X1    g082(.A(G57gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(G64gat), .ZN(new_n285_));
  AND3_X1   g084(.A1(new_n283_), .A2(new_n285_), .A3(KEYINPUT11), .ZN(new_n286_));
  AOI21_X1  g085(.A(KEYINPUT11), .B1(new_n283_), .B2(new_n285_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G71gat), .B(G78gat), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n286_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G57gat), .B(G64gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n290_), .A2(new_n288_), .A3(KEYINPUT11), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n281_), .B1(new_n289_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n290_), .A2(KEYINPUT11), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT11), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n284_), .A2(G64gat), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n282_), .A2(G57gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n295_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n288_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n294_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n300_), .A2(KEYINPUT67), .A3(new_n291_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n293_), .A2(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(G1gat), .B(G8gat), .Z(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  AND2_X1   g103(.A1(G15gat), .A2(G22gat), .ZN(new_n305_));
  NOR2_X1   g104(.A1(G15gat), .A2(G22gat), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT14), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n308_), .B1(G1gat), .B2(G8gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT70), .B1(new_n307_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT71), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G15gat), .B(G22gat), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT70), .ZN(new_n313_));
  INV_X1    g112(.A(G1gat), .ZN(new_n314_));
  INV_X1    g113(.A(G8gat), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT14), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n312_), .A2(new_n313_), .A3(new_n316_), .ZN(new_n317_));
  AND3_X1   g116(.A1(new_n310_), .A2(new_n311_), .A3(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n311_), .B1(new_n310_), .B2(new_n317_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n304_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  NOR3_X1   g119(.A1(new_n307_), .A2(new_n309_), .A3(KEYINPUT70), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n313_), .B1(new_n312_), .B2(new_n316_), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT71), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n310_), .A2(new_n311_), .A3(new_n317_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n303_), .A3(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n320_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G231gat), .A2(G233gat), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n326_), .A2(new_n327_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n302_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT73), .B1(new_n278_), .B2(new_n279_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n280_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  NOR3_X1   g131(.A1(new_n328_), .A2(new_n329_), .A3(new_n302_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n300_), .A2(new_n291_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n335_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n279_), .ZN(new_n337_));
  NOR3_X1   g136(.A1(new_n328_), .A2(new_n329_), .A3(new_n335_), .ZN(new_n338_));
  OAI22_X1  g137(.A1(new_n332_), .A2(new_n333_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT74), .ZN(new_n340_));
  AOI22_X1  g139(.A1(new_n228_), .A2(new_n230_), .B1(new_n226_), .B2(KEYINPUT8), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n301_), .B(new_n293_), .C1(new_n341_), .C2(new_n217_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT12), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n334_), .A2(new_n343_), .ZN(new_n344_));
  AOI22_X1  g143(.A1(new_n342_), .A2(new_n343_), .B1(new_n248_), .B2(new_n344_), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n300_), .A2(KEYINPUT67), .A3(new_n291_), .ZN(new_n346_));
  AOI21_X1  g145(.A(KEYINPUT67), .B1(new_n300_), .B2(new_n291_), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n244_), .B(new_n247_), .C1(new_n346_), .C2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G230gat), .A2(G233gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT64), .ZN(new_n350_));
  AND3_X1   g149(.A1(new_n348_), .A2(KEYINPUT68), .A3(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT68), .B1(new_n348_), .B2(new_n350_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n345_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n342_), .A2(new_n348_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n350_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G120gat), .B(G148gat), .ZN(new_n357_));
  INV_X1    g156(.A(G204gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(KEYINPUT5), .B(G176gat), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n359_), .B(new_n360_), .Z(new_n361_));
  NAND3_X1  g160(.A1(new_n353_), .A2(new_n356_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n361_), .B1(new_n353_), .B2(new_n356_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  OR2_X1    g164(.A1(new_n365_), .A2(KEYINPUT13), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(KEYINPUT13), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n271_), .A2(new_n340_), .A3(new_n366_), .A4(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT27), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G226gat), .A2(G233gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT19), .ZN(new_n371_));
  XOR2_X1   g170(.A(new_n371_), .B(KEYINPUT90), .Z(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(G169gat), .ZN(new_n374_));
  INV_X1    g173(.A(G176gat), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT22), .B(G169gat), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n378_), .A2(KEYINPUT81), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT81), .B1(new_n374_), .B2(KEYINPUT22), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n375_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n377_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT82), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT82), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n384_), .B(new_n377_), .C1(new_n379_), .C2(new_n381_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT78), .B(G190gat), .ZN(new_n386_));
  INV_X1    g185(.A(G183gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G183gat), .A2(G190gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT23), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n383_), .A2(new_n385_), .A3(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(G169gat), .A2(G176gat), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT24), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n390_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT80), .ZN(new_n397_));
  NOR3_X1   g196(.A1(new_n376_), .A2(new_n394_), .A3(new_n393_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n390_), .A2(new_n395_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT80), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n398_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT25), .B(G183gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT77), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT77), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n404_), .A2(new_n387_), .A3(KEYINPUT25), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n386_), .A2(KEYINPUT26), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT26), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(G190gat), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT79), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n406_), .A2(new_n407_), .A3(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n397_), .A2(new_n401_), .A3(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n392_), .A2(new_n413_), .ZN(new_n414_));
  XOR2_X1   g213(.A(G211gat), .B(G218gat), .Z(new_n415_));
  XNOR2_X1  g214(.A(G197gat), .B(G204gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT87), .B(KEYINPUT21), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n415_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n358_), .A2(G197gat), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT86), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(G197gat), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n420_), .A2(new_n422_), .A3(G204gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n358_), .A2(G197gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT21), .B1(new_n421_), .B2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n418_), .A2(new_n426_), .A3(KEYINPUT88), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(KEYINPUT88), .B1(new_n418_), .B2(new_n426_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G211gat), .B(G218gat), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT89), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT21), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n416_), .A2(new_n433_), .ZN(new_n434_));
  OAI22_X1  g233(.A1(new_n428_), .A2(new_n429_), .B1(new_n432_), .B2(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(KEYINPUT20), .B1(new_n414_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT92), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n376_), .B1(new_n378_), .B2(new_n375_), .ZN(new_n438_));
  INV_X1    g237(.A(G190gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n387_), .A2(new_n439_), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n390_), .A2(KEYINPUT91), .A3(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(KEYINPUT91), .B1(new_n390_), .B2(new_n440_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n438_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n398_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n439_), .A2(KEYINPUT26), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n402_), .A2(new_n409_), .A3(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n396_), .A2(new_n444_), .A3(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n443_), .A2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n437_), .B1(new_n435_), .B2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n436_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n435_), .A2(new_n437_), .A3(new_n448_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n373_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NOR3_X1   g251(.A1(new_n432_), .A2(new_n433_), .A3(new_n416_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n429_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n453_), .B1(new_n454_), .B2(new_n427_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n448_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n414_), .A2(new_n435_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n371_), .ZN(new_n459_));
  AND4_X1   g258(.A1(KEYINPUT20), .A2(new_n457_), .A3(new_n458_), .A4(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(KEYINPUT93), .B(KEYINPUT18), .Z(new_n461_));
  XNOR2_X1  g260(.A(G8gat), .B(G36gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G64gat), .B(G92gat), .ZN(new_n464_));
  XOR2_X1   g263(.A(new_n463_), .B(new_n464_), .Z(new_n465_));
  NOR3_X1   g264(.A1(new_n452_), .A2(new_n460_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n465_), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT92), .B1(new_n455_), .B2(new_n456_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n455_), .A2(new_n413_), .A3(new_n392_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n468_), .A2(KEYINPUT20), .A3(new_n451_), .A4(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n372_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n460_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n467_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n369_), .B1(new_n466_), .B2(new_n473_), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n457_), .A2(new_n458_), .A3(KEYINPUT20), .ZN(new_n475_));
  OAI22_X1  g274(.A1(new_n470_), .A2(new_n372_), .B1(new_n475_), .B2(new_n459_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(new_n465_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n471_), .A2(new_n472_), .A3(new_n467_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(KEYINPUT27), .A3(new_n478_), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n474_), .A2(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(G127gat), .B(G134gat), .Z(new_n481_));
  XOR2_X1   g280(.A(G113gat), .B(G120gat), .Z(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT31), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT83), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT84), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n486_), .B1(KEYINPUT84), .B2(new_n484_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT30), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n414_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n392_), .A2(new_n413_), .A3(KEYINPUT30), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(G227gat), .ZN(new_n492_));
  INV_X1    g291(.A(G233gat), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n491_), .A2(new_n494_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n489_), .B(new_n490_), .C1(new_n492_), .C2(new_n493_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G15gat), .B(G43gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G71gat), .B(G99gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n495_), .A2(new_n496_), .A3(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n500_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n487_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n495_), .A2(new_n496_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n499_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n495_), .A2(new_n496_), .A3(new_n500_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(new_n506_), .A3(new_n486_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n503_), .A2(new_n507_), .ZN(new_n508_));
  XOR2_X1   g307(.A(G155gat), .B(G162gat), .Z(new_n509_));
  INV_X1    g308(.A(KEYINPUT1), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n512_));
  INV_X1    g311(.A(G141gat), .ZN(new_n513_));
  INV_X1    g312(.A(G148gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G141gat), .A2(G148gat), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n511_), .A2(KEYINPUT85), .A3(new_n512_), .A4(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT85), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G155gat), .B(G162gat), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n520_), .A2(KEYINPUT1), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n515_), .A2(new_n512_), .A3(new_n516_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n519_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n518_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n515_), .B(KEYINPUT3), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n516_), .B(KEYINPUT2), .Z(new_n526_));
  OAI21_X1  g325(.A(new_n509_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n483_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n524_), .A2(new_n527_), .A3(new_n483_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(KEYINPUT4), .A3(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G225gat), .A2(G233gat), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n483_), .B1(new_n524_), .B2(new_n527_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT4), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n533_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n524_), .A2(new_n527_), .A3(new_n483_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n537_), .A2(new_n534_), .ZN(new_n538_));
  AOI22_X1  g337(.A1(new_n532_), .A2(new_n536_), .B1(new_n538_), .B2(new_n533_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G57gat), .B(G85gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G1gat), .B(G29gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(KEYINPUT97), .B1(new_n539_), .B2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n530_), .A2(new_n531_), .A3(new_n533_), .ZN(new_n546_));
  NOR3_X1   g345(.A1(new_n537_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n534_), .A2(new_n535_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n533_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n546_), .B1(new_n547_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT97), .ZN(new_n552_));
  INV_X1    g351(.A(new_n544_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n546_), .B(new_n544_), .C1(new_n547_), .C2(new_n550_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n545_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(G228gat), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n557_), .A2(new_n493_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n528_), .A2(KEYINPUT29), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n559_), .B1(new_n560_), .B2(new_n435_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n560_), .A2(new_n435_), .A3(new_n559_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n528_), .A2(KEYINPUT29), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n562_), .A2(new_n563_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n563_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n564_), .B1(new_n567_), .B2(new_n561_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(G22gat), .B(G50gat), .Z(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT28), .ZN(new_n571_));
  XOR2_X1   g370(.A(G78gat), .B(G106gat), .Z(new_n572_));
  XOR2_X1   g371(.A(new_n571_), .B(new_n572_), .Z(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n569_), .A2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n566_), .A2(new_n568_), .A3(new_n573_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n508_), .A2(new_n556_), .A3(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n480_), .A2(new_n578_), .A3(KEYINPUT98), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT98), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n575_), .A2(new_n576_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n556_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n581_), .A2(new_n582_), .A3(new_n507_), .A4(new_n503_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n474_), .A2(new_n479_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n580_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n579_), .A2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n556_), .B1(new_n576_), .B2(new_n575_), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n587_), .A2(new_n474_), .A3(new_n479_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n465_), .B1(new_n452_), .B2(new_n460_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n532_), .A2(new_n533_), .A3(new_n548_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n538_), .A2(new_n549_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n590_), .A2(new_n553_), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(KEYINPUT95), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT95), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n590_), .A2(new_n594_), .A3(new_n553_), .A4(new_n591_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n555_), .A2(KEYINPUT33), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT33), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n539_), .A2(new_n598_), .A3(new_n544_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n589_), .A2(new_n596_), .A3(new_n478_), .A4(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT96), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  AOI22_X1  g402(.A1(new_n593_), .A2(new_n595_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n604_), .A2(KEYINPUT96), .A3(new_n478_), .A4(new_n589_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n467_), .A2(KEYINPUT32), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n476_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n471_), .A2(new_n472_), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n556_), .B(new_n607_), .C1(new_n608_), .C2(new_n606_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n603_), .A2(new_n605_), .A3(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n588_), .B1(new_n610_), .B2(new_n581_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n508_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n586_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n320_), .A2(new_n251_), .A3(new_n325_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G229gat), .A2(G233gat), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT75), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n617_), .B1(new_n326_), .B2(new_n240_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n240_), .ZN(new_n619_));
  AOI211_X1 g418(.A(KEYINPUT75), .B(new_n619_), .C1(new_n320_), .C2(new_n325_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n616_), .B1(new_n618_), .B2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT76), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n320_), .A2(new_n325_), .A3(new_n619_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n623_), .B1(new_n618_), .B2(new_n620_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n615_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT76), .ZN(new_n627_));
  OAI211_X1 g426(.A(new_n616_), .B(new_n627_), .C1(new_n618_), .C2(new_n620_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n622_), .A2(new_n626_), .A3(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G113gat), .B(G141gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(G169gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(new_n422_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n629_), .A2(new_n633_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n622_), .A2(new_n626_), .A3(new_n628_), .A4(new_n632_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n613_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT99), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n613_), .A2(KEYINPUT99), .A3(new_n636_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n368_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n641_), .A2(new_n314_), .A3(new_n556_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT38), .ZN(new_n643_));
  OR2_X1    g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n613_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n366_), .A2(new_n367_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(new_n636_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n264_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n340_), .A2(new_n648_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n645_), .A2(new_n647_), .A3(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(G1gat), .B1(new_n651_), .B2(new_n582_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n642_), .A2(new_n643_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n644_), .A2(new_n652_), .A3(new_n653_), .ZN(G1324gat));
  NAND3_X1  g453(.A1(new_n641_), .A2(new_n315_), .A3(new_n584_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n647_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n649_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n613_), .A2(new_n584_), .A3(new_n656_), .A4(new_n657_), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n658_), .A2(KEYINPUT100), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT39), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n315_), .B1(new_n658_), .B2(KEYINPUT100), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n659_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n660_), .B1(new_n659_), .B2(new_n661_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n655_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  XOR2_X1   g463(.A(KEYINPUT101), .B(KEYINPUT40), .Z(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(G1325gat));
  OAI21_X1  g465(.A(G15gat), .B1(new_n651_), .B2(new_n508_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(KEYINPUT102), .B(KEYINPUT41), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n668_), .ZN(new_n670_));
  INV_X1    g469(.A(G15gat), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n641_), .A2(new_n671_), .A3(new_n612_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n669_), .A2(new_n670_), .A3(new_n672_), .ZN(G1326gat));
  NOR2_X1   g472(.A1(new_n581_), .A2(G22gat), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT104), .Z(new_n675_));
  NAND2_X1  g474(.A1(new_n641_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n650_), .A2(new_n577_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G22gat), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n678_), .A2(KEYINPUT103), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(KEYINPUT103), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n679_), .A2(KEYINPUT42), .A3(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT42), .B1(new_n679_), .B2(new_n680_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n676_), .B1(new_n681_), .B2(new_n682_), .ZN(G1327gat));
  NAND2_X1  g482(.A1(new_n639_), .A2(new_n640_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n646_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n340_), .A2(new_n648_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n685_), .A2(new_n687_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n684_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(G29gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n689_), .A2(new_n690_), .A3(new_n556_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n647_), .A2(new_n340_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n271_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n613_), .A2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(KEYINPUT43), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n613_), .A2(new_n697_), .A3(new_n694_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n693_), .B1(new_n696_), .B2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n698_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n697_), .B1(new_n613_), .B2(new_n694_), .ZN(new_n704_));
  OAI211_X1 g503(.A(KEYINPUT44), .B(new_n692_), .C1(new_n703_), .C2(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n702_), .A2(new_n556_), .A3(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n706_), .A2(new_n707_), .A3(G29gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n706_), .B2(G29gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n691_), .B1(new_n708_), .B2(new_n709_), .ZN(G1328gat));
  OAI21_X1  g509(.A(new_n584_), .B1(new_n699_), .B2(KEYINPUT44), .ZN(new_n711_));
  INV_X1    g510(.A(new_n705_), .ZN(new_n712_));
  OAI21_X1  g511(.A(G36gat), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n480_), .A2(G36gat), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n613_), .A2(KEYINPUT99), .A3(new_n636_), .ZN(new_n715_));
  AOI21_X1  g514(.A(KEYINPUT99), .B1(new_n613_), .B2(new_n636_), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n688_), .B(new_n714_), .C1(new_n715_), .C2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT106), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n684_), .A2(new_n719_), .A3(new_n688_), .A4(new_n714_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT45), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n718_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n718_), .B2(new_n720_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n713_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT46), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n713_), .B(KEYINPUT46), .C1(new_n722_), .C2(new_n723_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(G1329gat));
  NAND4_X1  g527(.A1(new_n702_), .A2(G43gat), .A3(new_n612_), .A4(new_n705_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n689_), .A2(new_n612_), .ZN(new_n730_));
  INV_X1    g529(.A(G43gat), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT108), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n729_), .A2(new_n732_), .A3(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n729_), .B2(new_n732_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1330gat));
  AOI21_X1  g536(.A(G50gat), .B1(new_n689_), .B2(new_n577_), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n702_), .A2(G50gat), .A3(new_n577_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(new_n705_), .ZN(G1331gat));
  NOR2_X1   g539(.A1(new_n646_), .A2(new_n636_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n645_), .A2(new_n649_), .A3(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n743_), .A2(G57gat), .A3(new_n556_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT110), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n339_), .B(KEYINPUT74), .Z(new_n746_));
  NOR2_X1   g545(.A1(new_n694_), .A2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n613_), .A2(new_n747_), .A3(new_n741_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT109), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n582_), .B1(new_n748_), .B2(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(G57gat), .B1(new_n750_), .B2(new_n752_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n745_), .A2(new_n753_), .ZN(G1332gat));
  AOI21_X1  g553(.A(new_n282_), .B1(new_n743_), .B2(new_n584_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT48), .Z(new_n756_));
  NAND3_X1  g555(.A1(new_n749_), .A2(new_n282_), .A3(new_n584_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(G1333gat));
  INV_X1    g557(.A(G71gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n743_), .B2(new_n612_), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT49), .Z(new_n761_));
  NAND3_X1  g560(.A1(new_n749_), .A2(new_n759_), .A3(new_n612_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(G1334gat));
  INV_X1    g562(.A(G78gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n764_), .B1(new_n743_), .B2(new_n577_), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT50), .Z(new_n766_));
  NAND3_X1  g565(.A1(new_n749_), .A2(new_n764_), .A3(new_n577_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(G1335gat));
  NOR3_X1   g567(.A1(new_n645_), .A2(new_n687_), .A3(new_n742_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n769_), .A2(new_n215_), .A3(new_n556_), .ZN(new_n770_));
  AOI211_X1 g569(.A(new_n340_), .B(new_n742_), .C1(new_n696_), .C2(new_n698_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n556_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n770_), .B1(new_n773_), .B2(new_n215_), .ZN(G1336gat));
  AOI21_X1  g573(.A(G92gat), .B1(new_n769_), .B2(new_n584_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n480_), .A2(new_n214_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n771_), .B2(new_n776_), .ZN(G1337gat));
  INV_X1    g576(.A(new_n210_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n769_), .A2(new_n612_), .A3(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT51), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n779_), .B1(KEYINPUT111), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n771_), .A2(new_n612_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n782_), .B2(G99gat), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n780_), .A2(KEYINPUT111), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n783_), .B(new_n784_), .ZN(G1338gat));
  NOR2_X1   g584(.A1(new_n742_), .A2(new_n340_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n577_), .B(new_n786_), .C1(new_n703_), .C2(new_n704_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n220_), .B1(new_n788_), .B2(KEYINPUT52), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(KEYINPUT112), .A3(new_n791_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n787_), .B(new_n789_), .C1(new_n788_), .C2(KEYINPUT52), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n769_), .A2(new_n220_), .A3(new_n577_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n792_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n795_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g595(.A1(new_n584_), .A2(new_n582_), .A3(new_n508_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n624_), .A2(new_n615_), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n625_), .B(new_n614_), .C1(new_n618_), .C2(new_n620_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(new_n633_), .A3(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n635_), .A2(new_n362_), .A3(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n343_), .B1(new_n233_), .B2(new_n302_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n248_), .A2(new_n344_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n348_), .A3(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n802_), .A2(KEYINPUT113), .A3(new_n348_), .A4(new_n803_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n806_), .A2(new_n355_), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n353_), .A2(new_n809_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n345_), .B(KEYINPUT55), .C1(new_n351_), .C2(new_n352_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n808_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n361_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n812_), .A2(KEYINPUT56), .A3(new_n813_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n801_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT58), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n694_), .B1(new_n818_), .B2(KEYINPUT58), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n363_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n812_), .A2(KEYINPUT56), .A3(new_n813_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT56), .B1(new_n812_), .B2(new_n813_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n822_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n635_), .A2(new_n800_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n826_), .A2(new_n365_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n264_), .B1(new_n825_), .B2(new_n828_), .ZN(new_n829_));
  XOR2_X1   g628(.A(KEYINPUT114), .B(KEYINPUT57), .Z(new_n830_));
  OAI22_X1  g629(.A1(new_n820_), .A2(new_n821_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT115), .B1(new_n829_), .B2(KEYINPUT57), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n829_), .A2(KEYINPUT115), .A3(KEYINPUT57), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n340_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n836_));
  INV_X1    g635(.A(new_n636_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n747_), .A2(new_n646_), .A3(new_n836_), .A4(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(KEYINPUT54), .B1(new_n368_), .B2(new_n636_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n581_), .B(new_n797_), .C1(new_n835_), .C2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(G113gat), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n843_), .A3(new_n636_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n841_), .A2(KEYINPUT59), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n825_), .A2(new_n828_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n847_), .A2(KEYINPUT57), .A3(new_n648_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT115), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n830_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n816_), .A2(new_n817_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n827_), .B1(new_n852_), .B2(new_n822_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n851_), .B1(new_n853_), .B2(new_n264_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n823_), .A2(new_n824_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(new_n801_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n857_), .A2(new_n819_), .A3(new_n694_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n850_), .A2(new_n834_), .A3(new_n854_), .A4(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n746_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n840_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n577_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT59), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n862_), .A2(new_n863_), .A3(new_n797_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n846_), .A2(new_n865_), .A3(new_n837_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n844_), .B1(new_n866_), .B2(new_n843_), .ZN(G1340gat));
  INV_X1    g666(.A(G120gat), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(KEYINPUT60), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n646_), .B2(KEYINPUT60), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT116), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n869_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n842_), .B(new_n872_), .C1(new_n871_), .C2(new_n870_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n846_), .A2(new_n865_), .A3(new_n646_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n874_), .B2(new_n868_), .ZN(G1341gat));
  INV_X1    g674(.A(G127gat), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n746_), .A2(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n845_), .A2(new_n864_), .A3(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT57), .ZN(new_n879_));
  NOR4_X1   g678(.A1(new_n853_), .A2(new_n849_), .A3(new_n879_), .A4(new_n264_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n831_), .A2(new_n880_), .A3(new_n832_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n861_), .B1(new_n881_), .B2(new_n340_), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n882_), .A2(new_n581_), .A3(new_n340_), .A4(new_n797_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT117), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n883_), .A2(new_n884_), .A3(new_n876_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n883_), .B2(new_n876_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n878_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT118), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n878_), .B(KEYINPUT118), .C1(new_n885_), .C2(new_n886_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1342gat));
  AOI21_X1  g690(.A(G134gat), .B1(new_n842_), .B2(new_n264_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n846_), .A2(new_n865_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n694_), .A2(G134gat), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(KEYINPUT119), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n892_), .B1(new_n893_), .B2(new_n895_), .ZN(G1343gat));
  NOR3_X1   g695(.A1(new_n612_), .A2(new_n582_), .A3(new_n581_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n882_), .A2(new_n480_), .A3(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n837_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(new_n513_), .ZN(G1344gat));
  NOR2_X1   g699(.A1(new_n898_), .A2(new_n646_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(new_n514_), .ZN(G1345gat));
  NOR2_X1   g701(.A1(new_n898_), .A2(new_n746_), .ZN(new_n903_));
  XOR2_X1   g702(.A(KEYINPUT61), .B(G155gat), .Z(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1346gat));
  OAI21_X1  g704(.A(G162gat), .B1(new_n898_), .B2(new_n271_), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n648_), .A2(G162gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n898_), .B2(new_n907_), .ZN(G1347gat));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n840_), .B1(new_n859_), .B2(new_n746_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n508_), .A2(new_n556_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n584_), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n910_), .A2(new_n577_), .A3(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n636_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n909_), .B1(new_n914_), .B2(G169gat), .ZN(new_n915_));
  AOI211_X1 g714(.A(KEYINPUT62), .B(new_n374_), .C1(new_n913_), .C2(new_n636_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n912_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n862_), .A2(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT120), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n913_), .A2(KEYINPUT120), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n636_), .A2(new_n378_), .ZN(new_n923_));
  OAI22_X1  g722(.A1(new_n915_), .A2(new_n916_), .B1(new_n922_), .B2(new_n923_), .ZN(G1348gat));
  NOR3_X1   g723(.A1(new_n918_), .A2(new_n375_), .A3(new_n646_), .ZN(new_n925_));
  AOI21_X1  g724(.A(KEYINPUT120), .B1(new_n862_), .B2(new_n917_), .ZN(new_n926_));
  NOR4_X1   g725(.A1(new_n910_), .A2(new_n919_), .A3(new_n577_), .A4(new_n912_), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n926_), .A2(new_n927_), .A3(new_n646_), .ZN(new_n928_));
  OAI21_X1  g727(.A(KEYINPUT121), .B1(new_n928_), .B2(G176gat), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n920_), .A2(new_n685_), .A3(new_n921_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT121), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n930_), .A2(new_n931_), .A3(new_n375_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n925_), .B1(new_n929_), .B2(new_n932_), .ZN(G1349gat));
  NOR2_X1   g732(.A1(new_n746_), .A2(new_n402_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n920_), .A2(new_n921_), .A3(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT122), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  OAI21_X1  g736(.A(KEYINPUT123), .B1(new_n918_), .B2(new_n746_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT123), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n913_), .A2(new_n939_), .A3(new_n340_), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n938_), .A2(new_n387_), .A3(new_n940_), .ZN(new_n941_));
  NAND4_X1  g740(.A1(new_n920_), .A2(new_n921_), .A3(KEYINPUT122), .A4(new_n934_), .ZN(new_n942_));
  AND3_X1   g741(.A1(new_n937_), .A2(new_n941_), .A3(new_n942_), .ZN(G1350gat));
  OAI21_X1  g742(.A(G190gat), .B1(new_n922_), .B2(new_n271_), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n264_), .A2(new_n409_), .A3(new_n445_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n944_), .B1(new_n922_), .B2(new_n945_), .ZN(G1351gat));
  AND3_X1   g745(.A1(new_n584_), .A2(new_n587_), .A3(new_n508_), .ZN(new_n947_));
  AND2_X1   g746(.A1(new_n882_), .A2(new_n947_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n948_), .A2(new_n636_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n949_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g749(.A1(new_n948_), .A2(new_n685_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n952_));
  XOR2_X1   g751(.A(new_n952_), .B(KEYINPUT125), .Z(new_n953_));
  XNOR2_X1  g752(.A(new_n951_), .B(new_n953_), .ZN(G1353gat));
  NAND2_X1  g753(.A1(new_n948_), .A2(new_n340_), .ZN(new_n955_));
  NOR2_X1   g754(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n956_));
  AND2_X1   g755(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n957_));
  NOR3_X1   g756(.A1(new_n955_), .A2(new_n956_), .A3(new_n957_), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n958_), .B1(new_n955_), .B2(new_n956_), .ZN(G1354gat));
  NAND2_X1  g758(.A1(new_n948_), .A2(new_n264_), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n960_), .B(KEYINPUT126), .ZN(new_n961_));
  XNOR2_X1  g760(.A(KEYINPUT127), .B(G218gat), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n271_), .A2(new_n962_), .ZN(new_n963_));
  AOI22_X1  g762(.A1(new_n961_), .A2(new_n962_), .B1(new_n948_), .B2(new_n963_), .ZN(G1355gat));
endmodule


