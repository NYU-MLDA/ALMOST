//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 1 0 1 0 0 1 1 1 1 1 0 1 0 0 0 1 1 0 1 1 0 1 1 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 1 1 0 1 0 0 1 0 1 0 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n814_, new_n815_, new_n816_, new_n817_, new_n819_,
    new_n820_, new_n821_, new_n823_, new_n824_, new_n825_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n832_, new_n833_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n877_, new_n878_, new_n879_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_;
  XNOR2_X1  g000(.A(G120gat), .B(G148gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT5), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G176gat), .B(G204gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT73), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G230gat), .A2(G233gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G92gat), .ZN(new_n208_));
  AOI21_X1  g007(.A(KEYINPUT9), .B1(new_n208_), .B2(G85gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G85gat), .A2(G92gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n210_), .B1(new_n211_), .B2(KEYINPUT66), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n212_), .B1(KEYINPUT66), .B2(new_n210_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n209_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT67), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT6), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT68), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT10), .B(G99gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n220_), .A2(G106gat), .ZN(new_n221_));
  OR2_X1    g020(.A1(new_n221_), .A2(KEYINPUT64), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(KEYINPUT64), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n219_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n215_), .A2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G57gat), .B(G64gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT71), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT11), .ZN(new_n228_));
  XOR2_X1   g027(.A(G71gat), .B(G78gat), .Z(new_n229_));
  OR2_X1    g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n226_), .A2(KEYINPUT71), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n226_), .A2(KEYINPUT71), .ZN(new_n232_));
  OR3_X1    g031(.A1(new_n231_), .A2(new_n232_), .A3(KEYINPUT11), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n233_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n230_), .A2(new_n234_), .ZN(new_n235_));
  NOR3_X1   g034(.A1(KEYINPUT69), .A2(G99gat), .A3(G106gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n236_), .B(KEYINPUT7), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT70), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT70), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n237_), .A2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(new_n241_), .A3(new_n217_), .ZN(new_n242_));
  XOR2_X1   g041(.A(G85gat), .B(G92gat), .Z(new_n243_));
  NAND3_X1  g042(.A1(new_n242_), .A2(KEYINPUT8), .A3(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n243_), .B1(new_n219_), .B2(new_n238_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT8), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n225_), .A2(new_n235_), .A3(new_n244_), .A4(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT12), .ZN(new_n249_));
  AOI22_X1  g048(.A1(new_n215_), .A2(new_n224_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n235_), .B1(new_n250_), .B2(new_n244_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  AOI211_X1 g051(.A(KEYINPUT12), .B(new_n235_), .C1(new_n250_), .C2(new_n244_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n207_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n225_), .A2(new_n244_), .A3(new_n247_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n235_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT72), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(new_n258_), .A3(new_n248_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n207_), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n259_), .B(new_n260_), .C1(new_n258_), .C2(new_n257_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n206_), .B1(new_n254_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n254_), .A2(new_n261_), .A3(new_n206_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(KEYINPUT13), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT13), .ZN(new_n266_));
  INV_X1    g065(.A(new_n264_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n266_), .B1(new_n267_), .B2(new_n262_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT30), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT85), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT22), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n273_), .A2(G169gat), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT84), .ZN(new_n275_));
  AOI21_X1  g074(.A(G176gat), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(G169gat), .B1(new_n273_), .B2(KEYINPUT84), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n272_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(G169gat), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n275_), .A2(new_n279_), .A3(KEYINPUT22), .ZN(new_n280_));
  INV_X1    g079(.A(G176gat), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n277_), .A2(new_n280_), .A3(new_n272_), .A4(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT86), .B1(new_n278_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT83), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT23), .ZN(new_n288_));
  NOR2_X1   g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT23), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n286_), .A2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n288_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n277_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT85), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT86), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n295_), .A2(new_n296_), .A3(new_n283_), .A4(new_n282_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n285_), .A2(new_n293_), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT87), .ZN(new_n299_));
  MUX2_X1   g098(.A(new_n286_), .B(new_n287_), .S(new_n291_), .Z(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT25), .B(G183gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT26), .B(G190gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n279_), .A2(new_n281_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n304_), .A2(KEYINPUT24), .A3(new_n283_), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n304_), .A2(KEYINPUT24), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n300_), .A2(new_n303_), .A3(new_n305_), .A4(new_n306_), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n298_), .A2(new_n299_), .A3(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n299_), .B1(new_n298_), .B2(new_n307_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n271_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n298_), .A2(new_n307_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT87), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n298_), .A2(new_n299_), .A3(new_n307_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n312_), .A2(KEYINPUT30), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G227gat), .A2(G233gat), .ZN(new_n315_));
  INV_X1    g114(.A(G15gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(G71gat), .ZN(new_n318_));
  XOR2_X1   g117(.A(KEYINPUT88), .B(G43gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(G99gat), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n318_), .B(new_n320_), .Z(new_n321_));
  NAND4_X1  g120(.A1(new_n310_), .A2(new_n314_), .A3(KEYINPUT89), .A4(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n310_), .A2(new_n314_), .A3(KEYINPUT89), .ZN(new_n323_));
  INV_X1    g122(.A(new_n321_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(KEYINPUT89), .B1(new_n310_), .B2(new_n314_), .ZN(new_n326_));
  OAI211_X1 g125(.A(KEYINPUT90), .B(new_n322_), .C1(new_n325_), .C2(new_n326_), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n327_), .A2(KEYINPUT91), .ZN(new_n328_));
  XOR2_X1   g127(.A(G127gat), .B(G134gat), .Z(new_n329_));
  XOR2_X1   g128(.A(G113gat), .B(G120gat), .Z(new_n330_));
  XOR2_X1   g129(.A(new_n329_), .B(new_n330_), .Z(new_n331_));
  XOR2_X1   g130(.A(new_n331_), .B(KEYINPUT31), .Z(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n322_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT90), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n333_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n327_), .A2(KEYINPUT91), .ZN(new_n337_));
  AND3_X1   g136(.A1(new_n328_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n336_), .B1(new_n328_), .B2(new_n337_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(G197gat), .B(G204gat), .Z(new_n341_));
  OR2_X1    g140(.A1(new_n341_), .A2(KEYINPUT21), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(KEYINPUT21), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G211gat), .B(G218gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n343_), .A2(new_n344_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT94), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G141gat), .A2(G148gat), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT92), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(KEYINPUT92), .A2(G141gat), .A3(G148gat), .ZN(new_n353_));
  INV_X1    g152(.A(G141gat), .ZN(new_n354_));
  INV_X1    g153(.A(G148gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n352_), .A2(new_n353_), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G155gat), .A2(G162gat), .ZN(new_n358_));
  NOR2_X1   g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n358_), .B1(new_n359_), .B2(KEYINPUT1), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT93), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT1), .ZN(new_n362_));
  INV_X1    g161(.A(new_n358_), .ZN(new_n363_));
  AOI22_X1  g162(.A1(new_n360_), .A2(new_n361_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  OAI211_X1 g163(.A(KEYINPUT93), .B(new_n358_), .C1(new_n359_), .C2(KEYINPUT1), .ZN(new_n365_));
  AOI211_X1 g164(.A(new_n349_), .B(new_n357_), .C1(new_n364_), .C2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n360_), .A2(new_n361_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n363_), .A2(new_n362_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n367_), .A2(new_n365_), .A3(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n357_), .ZN(new_n370_));
  AOI21_X1  g169(.A(KEYINPUT94), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT3), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n373_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n374_));
  AOI21_X1  g173(.A(KEYINPUT2), .B1(new_n353_), .B2(KEYINPUT95), .ZN(new_n375_));
  NAND2_X1  g174(.A1(KEYINPUT95), .A2(KEYINPUT2), .ZN(new_n376_));
  AOI22_X1  g175(.A1(new_n376_), .A2(KEYINPUT92), .B1(G141gat), .B2(G148gat), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n372_), .B(new_n374_), .C1(new_n375_), .C2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n363_), .A2(new_n359_), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n378_), .A2(KEYINPUT96), .A3(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(KEYINPUT96), .B1(new_n378_), .B2(new_n379_), .ZN(new_n381_));
  OAI22_X1  g180(.A1(new_n366_), .A2(new_n371_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n348_), .B1(new_n382_), .B2(KEYINPUT29), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G228gat), .A2(G233gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT97), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT97), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n383_), .A2(new_n387_), .A3(new_n384_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n382_), .A2(KEYINPUT29), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n347_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n391_), .A2(KEYINPUT98), .A3(G228gat), .A4(G233gat), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT98), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n393_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n389_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G78gat), .B(G106gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n386_), .A2(new_n388_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n397_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT99), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n398_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n382_), .A2(KEYINPUT29), .ZN(new_n404_));
  XOR2_X1   g203(.A(new_n404_), .B(KEYINPUT28), .Z(new_n405_));
  XNOR2_X1  g204(.A(G22gat), .B(G50gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n396_), .A2(KEYINPUT99), .A3(new_n397_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n403_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n398_), .A2(KEYINPUT100), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT100), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n396_), .A2(new_n412_), .A3(new_n397_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n411_), .A2(new_n413_), .A3(new_n401_), .A4(new_n407_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G8gat), .B(G36gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT18), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G64gat), .B(G92gat), .ZN(new_n418_));
  XOR2_X1   g217(.A(new_n417_), .B(new_n418_), .Z(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G226gat), .A2(G233gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT19), .ZN(new_n422_));
  NOR3_X1   g221(.A1(new_n308_), .A2(new_n309_), .A3(new_n347_), .ZN(new_n423_));
  XOR2_X1   g222(.A(KEYINPUT22), .B(G169gat), .Z(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(new_n281_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(new_n283_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n427_), .B1(new_n300_), .B2(new_n290_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n303_), .A2(new_n305_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n288_), .A2(new_n292_), .A3(new_n306_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT101), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n429_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  OR2_X1    g231(.A1(new_n430_), .A2(new_n431_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n428_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT20), .B1(new_n434_), .B2(new_n348_), .ZN(new_n435_));
  OAI211_X1 g234(.A(KEYINPUT102), .B(new_n422_), .C1(new_n423_), .C2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n347_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT20), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n438_), .B1(new_n434_), .B2(new_n348_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n422_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n437_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n436_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n433_), .A2(new_n432_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n428_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n438_), .B1(new_n445_), .B2(new_n347_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n312_), .A2(new_n348_), .A3(new_n313_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT102), .B1(new_n448_), .B2(new_n422_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n420_), .B1(new_n442_), .B2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n422_), .B1(new_n423_), .B2(new_n435_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT102), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n453_), .A2(new_n419_), .A3(new_n441_), .A4(new_n436_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n450_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT27), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n446_), .A2(new_n447_), .A3(new_n440_), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n437_), .A2(new_n439_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n458_), .B1(new_n459_), .B2(new_n440_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n456_), .B1(new_n460_), .B2(new_n420_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n454_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n457_), .A2(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n415_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n382_), .A2(new_n331_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT96), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n374_), .A2(new_n372_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n377_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n353_), .A2(KEYINPUT95), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT2), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n467_), .B1(new_n468_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n379_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n466_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n378_), .A2(KEYINPUT96), .A3(new_n379_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n331_), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n476_), .B(new_n477_), .C1(new_n371_), .C2(new_n366_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n465_), .A2(KEYINPUT4), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT4), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n382_), .A2(new_n480_), .A3(new_n331_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G225gat), .A2(G233gat), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n482_), .A2(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(G1gat), .B(G29gat), .Z(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT103), .B(KEYINPUT0), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G57gat), .B(G85gat), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n488_), .B(new_n489_), .Z(new_n490_));
  AOI21_X1  g289(.A(new_n484_), .B1(new_n465_), .B2(new_n478_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n485_), .A2(new_n490_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT106), .ZN(new_n494_));
  INV_X1    g293(.A(new_n490_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n483_), .B1(new_n479_), .B2(new_n481_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n495_), .B1(new_n496_), .B2(new_n491_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n493_), .A2(new_n494_), .A3(new_n497_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n485_), .A2(KEYINPUT106), .A3(new_n490_), .A4(new_n492_), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n340_), .A2(new_n464_), .A3(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n442_), .A2(new_n449_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n419_), .A2(KEYINPUT32), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n503_), .A2(KEYINPUT105), .A3(new_n504_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n453_), .A2(new_n441_), .A3(new_n436_), .A4(new_n504_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT105), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n460_), .A2(KEYINPUT32), .A3(new_n419_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n500_), .A2(new_n505_), .A3(new_n508_), .A4(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n497_), .A2(KEYINPUT33), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT33), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n512_), .B(new_n495_), .C1(new_n496_), .C2(new_n491_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n482_), .A2(new_n484_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n465_), .A2(new_n484_), .A3(new_n478_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n490_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n514_), .A2(new_n450_), .A3(new_n454_), .A4(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT104), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n518_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n523_), .A2(KEYINPUT104), .A3(new_n454_), .A4(new_n450_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n510_), .A2(new_n522_), .A3(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n415_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n500_), .B1(new_n410_), .B2(new_n414_), .ZN(new_n527_));
  AOI22_X1  g326(.A1(new_n455_), .A2(new_n456_), .B1(new_n461_), .B2(new_n454_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n525_), .A2(new_n526_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n502_), .B1(new_n529_), .B2(new_n340_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G15gat), .B(G22gat), .ZN(new_n531_));
  INV_X1    g330(.A(G1gat), .ZN(new_n532_));
  INV_X1    g331(.A(G8gat), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT14), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n531_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G1gat), .B(G8gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G29gat), .B(G36gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G43gat), .B(G50gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n537_), .B(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G229gat), .A2(G233gat), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT78), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n540_), .B(KEYINPUT15), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n537_), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n537_), .A2(new_n541_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n548_), .A2(new_n543_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT79), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n551_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n546_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(G113gat), .B(G141gat), .Z(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT80), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n556_), .B(KEYINPUT81), .Z(new_n557_));
  XNOR2_X1  g356(.A(G169gat), .B(G197gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n554_), .A2(new_n560_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n546_), .A2(new_n552_), .A3(new_n553_), .A4(new_n559_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n561_), .A2(KEYINPUT82), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT82), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n554_), .A2(new_n564_), .A3(new_n560_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n530_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n537_), .B(new_n569_), .Z(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(new_n235_), .ZN(new_n571_));
  XOR2_X1   g370(.A(G127gat), .B(G155gat), .Z(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT16), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G183gat), .B(G211gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT76), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT17), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n575_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n571_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n575_), .A2(new_n577_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n578_), .A2(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n571_), .A2(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT77), .B1(new_n580_), .B2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT77), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n579_), .B(new_n585_), .C1(new_n571_), .C2(new_n582_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n255_), .A2(new_n547_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT35), .ZN(new_n592_));
  AOI21_X1  g391(.A(KEYINPUT75), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n588_), .B(new_n593_), .C1(new_n255_), .C2(new_n541_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n591_), .A2(new_n592_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G190gat), .B(G218gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G134gat), .B(G162gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n596_), .A2(KEYINPUT36), .A3(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n599_), .B(KEYINPUT36), .Z(new_n601_));
  AND2_X1   g400(.A1(new_n596_), .A2(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT37), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(KEYINPUT37), .B1(new_n600_), .B2(new_n602_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  AND4_X1   g406(.A1(new_n270_), .A2(new_n568_), .A3(new_n587_), .A4(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n608_), .A2(new_n532_), .A3(new_n500_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT38), .ZN(new_n610_));
  INV_X1    g409(.A(new_n603_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n530_), .A2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n580_), .A2(new_n583_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n269_), .A2(new_n614_), .A3(new_n566_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT107), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n617_), .A2(new_n500_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n610_), .B1(new_n618_), .B2(new_n532_), .ZN(G1324gat));
  NAND3_X1  g418(.A1(new_n608_), .A2(new_n533_), .A3(new_n463_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n612_), .A2(new_n463_), .A3(new_n615_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT39), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n621_), .A2(new_n622_), .A3(G8gat), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n622_), .B1(new_n621_), .B2(G8gat), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n620_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g425(.A1(new_n608_), .A2(new_n316_), .A3(new_n340_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n617_), .A2(new_n340_), .ZN(new_n628_));
  AOI21_X1  g427(.A(KEYINPUT41), .B1(new_n628_), .B2(G15gat), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT41), .ZN(new_n630_));
  AOI211_X1 g429(.A(new_n630_), .B(new_n316_), .C1(new_n617_), .C2(new_n340_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n627_), .B1(new_n629_), .B2(new_n631_), .ZN(G1326gat));
  INV_X1    g431(.A(G22gat), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n608_), .A2(new_n633_), .A3(new_n415_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT42), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n617_), .A2(new_n415_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n635_), .B1(new_n636_), .B2(G22gat), .ZN(new_n637_));
  AOI211_X1 g436(.A(KEYINPUT42), .B(new_n633_), .C1(new_n617_), .C2(new_n415_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n634_), .B1(new_n637_), .B2(new_n638_), .ZN(G1327gat));
  INV_X1    g438(.A(new_n587_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n603_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n568_), .A2(new_n270_), .A3(new_n642_), .ZN(new_n643_));
  OR3_X1    g442(.A1(new_n643_), .A2(G29gat), .A3(new_n501_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n269_), .A2(new_n566_), .A3(new_n587_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT43), .ZN(new_n646_));
  INV_X1    g445(.A(new_n607_), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n530_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n646_), .B1(new_n530_), .B2(new_n647_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n645_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT44), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  OAI211_X1 g451(.A(KEYINPUT44), .B(new_n645_), .C1(new_n648_), .C2(new_n649_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(KEYINPUT108), .B1(new_n654_), .B2(new_n500_), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n652_), .A2(KEYINPUT108), .A3(new_n500_), .A4(new_n653_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(G29gat), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n644_), .B1(new_n655_), .B2(new_n657_), .ZN(G1328gat));
  NAND3_X1  g457(.A1(new_n652_), .A2(new_n463_), .A3(new_n653_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(G36gat), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n528_), .A2(G36gat), .ZN(new_n661_));
  OR3_X1    g460(.A1(new_n643_), .A2(KEYINPUT45), .A3(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(KEYINPUT45), .B1(new_n643_), .B2(new_n661_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n660_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT46), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n660_), .A2(KEYINPUT46), .A3(new_n664_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1329gat));
  NAND3_X1  g468(.A1(new_n652_), .A2(new_n340_), .A3(new_n653_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(G43gat), .ZN(new_n671_));
  INV_X1    g470(.A(new_n340_), .ZN(new_n672_));
  OR3_X1    g471(.A1(new_n643_), .A2(G43gat), .A3(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n671_), .A2(new_n673_), .A3(new_n675_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1330gat));
  NAND3_X1  g478(.A1(new_n652_), .A2(new_n415_), .A3(new_n653_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT110), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n680_), .A2(new_n681_), .A3(G50gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n680_), .B2(G50gat), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n526_), .A2(G50gat), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT111), .ZN(new_n685_));
  OAI22_X1  g484(.A1(new_n682_), .A2(new_n683_), .B1(new_n643_), .B2(new_n685_), .ZN(G1331gat));
  AND2_X1   g485(.A1(new_n530_), .A2(new_n566_), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n647_), .A2(new_n270_), .A3(new_n640_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(G57gat), .B1(new_n689_), .B2(new_n500_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT112), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n566_), .A2(new_n587_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n270_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n612_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(G57gat), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n694_), .A2(new_n695_), .A3(new_n501_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n691_), .A2(new_n696_), .ZN(G1332gat));
  OAI21_X1  g496(.A(G64gat), .B1(new_n694_), .B2(new_n528_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT48), .ZN(new_n699_));
  INV_X1    g498(.A(new_n689_), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n528_), .A2(G64gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n699_), .B1(new_n700_), .B2(new_n701_), .ZN(G1333gat));
  OAI21_X1  g501(.A(G71gat), .B1(new_n694_), .B2(new_n672_), .ZN(new_n703_));
  XOR2_X1   g502(.A(KEYINPUT113), .B(KEYINPUT49), .Z(new_n704_));
  XNOR2_X1  g503(.A(new_n703_), .B(new_n704_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n672_), .A2(G71gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(new_n700_), .B2(new_n706_), .ZN(G1334gat));
  OAI21_X1  g506(.A(G78gat), .B1(new_n694_), .B2(new_n526_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT50), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n526_), .A2(G78gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n709_), .B1(new_n700_), .B2(new_n710_), .ZN(G1335gat));
  OR2_X1    g510(.A1(new_n648_), .A2(new_n649_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n270_), .A2(new_n567_), .A3(new_n587_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(G85gat), .B1(new_n714_), .B2(new_n501_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n687_), .A2(new_n269_), .A3(new_n642_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(KEYINPUT114), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT114), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n687_), .A2(new_n718_), .A3(new_n269_), .A4(new_n642_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n501_), .A2(G85gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n715_), .B1(new_n721_), .B2(new_n722_), .ZN(G1336gat));
  AOI21_X1  g522(.A(G92gat), .B1(new_n720_), .B2(new_n463_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n714_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n463_), .A2(new_n208_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT115), .Z(new_n727_));
  AOI21_X1  g526(.A(new_n724_), .B1(new_n725_), .B2(new_n727_), .ZN(G1337gat));
  OAI21_X1  g527(.A(G99gat), .B1(new_n714_), .B2(new_n672_), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n672_), .A2(new_n220_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(new_n721_), .B2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT51), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT51), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n729_), .B(new_n733_), .C1(new_n721_), .C2(new_n730_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(G1338gat));
  INV_X1    g534(.A(G106gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n720_), .A2(new_n736_), .A3(new_n415_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT52), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n415_), .B(new_n713_), .C1(new_n648_), .C2(new_n649_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(G106gat), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n739_), .A2(new_n738_), .A3(G106gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n737_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT53), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT53), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n737_), .B(new_n744_), .C1(new_n740_), .C2(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1339gat));
  NAND3_X1  g545(.A1(new_n548_), .A2(new_n544_), .A3(new_n549_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n542_), .A2(new_n543_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n560_), .A2(new_n747_), .A3(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n562_), .A2(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n750_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n751_));
  OAI211_X1 g550(.A(KEYINPUT55), .B(new_n207_), .C1(new_n252_), .C2(new_n253_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n249_), .A2(new_n251_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n257_), .A2(KEYINPUT12), .A3(new_n248_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n753_), .A2(new_n754_), .A3(new_n260_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n752_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT55), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT118), .B1(new_n254_), .B2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n260_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT118), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n760_), .A2(new_n761_), .A3(KEYINPUT55), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n757_), .B1(new_n759_), .B2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n763_), .A2(KEYINPUT56), .A3(new_n205_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT56), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n761_), .B1(new_n760_), .B2(KEYINPUT55), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n254_), .A2(KEYINPUT118), .A3(new_n758_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n756_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n205_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n765_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n764_), .A2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n254_), .A2(new_n261_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n772_), .A2(new_n205_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n566_), .A2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n751_), .B1(new_n771_), .B2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(KEYINPUT57), .B1(new_n775_), .B2(new_n603_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT57), .ZN(new_n777_));
  INV_X1    g576(.A(new_n774_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n778_), .B1(new_n770_), .B2(new_n764_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n777_), .B(new_n611_), .C1(new_n779_), .C2(new_n751_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n776_), .A2(new_n780_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n773_), .A2(new_n750_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT58), .B1(new_n771_), .B2(new_n782_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n783_), .A2(new_n607_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n771_), .A2(KEYINPUT58), .A3(new_n782_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n781_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n614_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT116), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n692_), .A2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n566_), .A2(KEYINPUT116), .A3(new_n587_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n790_), .A2(new_n265_), .A3(new_n268_), .A4(new_n791_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n792_), .A2(KEYINPUT117), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n607_), .B1(new_n792_), .B2(KEYINPUT117), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT54), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  OR2_X1    g594(.A1(new_n792_), .A2(KEYINPUT117), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n792_), .A2(KEYINPUT117), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT54), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n796_), .A2(new_n797_), .A3(new_n798_), .A4(new_n607_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n795_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n788_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n340_), .A2(new_n464_), .A3(new_n500_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(G113gat), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(new_n805_), .A3(new_n567_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT59), .ZN(new_n807_));
  INV_X1    g606(.A(new_n803_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n807_), .B1(new_n801_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n787_), .A2(new_n640_), .ZN(new_n810_));
  AOI211_X1 g609(.A(KEYINPUT59), .B(new_n803_), .C1(new_n810_), .C2(new_n800_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n809_), .A2(new_n811_), .A3(new_n566_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n806_), .B1(new_n812_), .B2(new_n805_), .ZN(G1340gat));
  INV_X1    g612(.A(G120gat), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n270_), .B2(KEYINPUT60), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n804_), .B(new_n815_), .C1(KEYINPUT60), .C2(new_n814_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n809_), .A2(new_n811_), .A3(new_n270_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n816_), .B1(new_n817_), .B2(new_n814_), .ZN(G1341gat));
  INV_X1    g617(.A(G127gat), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n804_), .A2(new_n819_), .A3(new_n587_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n809_), .A2(new_n811_), .A3(new_n614_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n820_), .B1(new_n821_), .B2(new_n819_), .ZN(G1342gat));
  INV_X1    g621(.A(G134gat), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n804_), .A2(new_n823_), .A3(new_n603_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n809_), .A2(new_n811_), .A3(new_n607_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n825_), .B2(new_n823_), .ZN(G1343gat));
  NOR4_X1   g625(.A1(new_n340_), .A2(new_n526_), .A3(new_n501_), .A4(new_n463_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n801_), .A2(new_n827_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n828_), .A2(new_n566_), .ZN(new_n829_));
  XOR2_X1   g628(.A(KEYINPUT119), .B(G141gat), .Z(new_n830_));
  XNOR2_X1  g629(.A(new_n829_), .B(new_n830_), .ZN(G1344gat));
  NOR2_X1   g630(.A1(new_n828_), .A2(new_n270_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(KEYINPUT120), .B(G148gat), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n832_), .B(new_n833_), .ZN(G1345gat));
  INV_X1    g633(.A(KEYINPUT121), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n801_), .A2(new_n835_), .A3(new_n587_), .A4(new_n827_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n613_), .B1(new_n781_), .B2(new_n786_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n795_), .A2(new_n799_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n587_), .B(new_n827_), .C1(new_n837_), .C2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT121), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n836_), .A2(new_n840_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(KEYINPUT61), .B(G155gat), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n841_), .B(new_n842_), .ZN(G1346gat));
  OAI211_X1 g642(.A(new_n603_), .B(new_n827_), .C1(new_n837_), .C2(new_n838_), .ZN(new_n844_));
  INV_X1    g643(.A(G162gat), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n647_), .A2(G162gat), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(KEYINPUT122), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n801_), .A2(new_n827_), .A3(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n846_), .A2(new_n849_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(KEYINPUT123), .ZN(G1347gat));
  NOR3_X1   g650(.A1(new_n672_), .A2(new_n500_), .A3(new_n528_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n852_), .A2(new_n526_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n587_), .B1(new_n781_), .B2(new_n786_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n567_), .B(new_n853_), .C1(new_n854_), .C2(new_n838_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n855_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n810_), .A2(new_n800_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n857_), .A2(new_n425_), .A3(new_n567_), .A4(new_n853_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(KEYINPUT62), .B1(new_n855_), .B2(G169gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(KEYINPUT124), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n855_), .A2(G169gat), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT62), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT124), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n864_), .A2(new_n865_), .A3(new_n858_), .A4(new_n856_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n861_), .A2(new_n866_), .ZN(G1348gat));
  AND2_X1   g666(.A1(new_n857_), .A2(new_n853_), .ZN(new_n868_));
  AOI21_X1  g667(.A(G176gat), .B1(new_n868_), .B2(new_n269_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n802_), .A2(new_n415_), .ZN(new_n870_));
  AND3_X1   g669(.A1(new_n852_), .A2(G176gat), .A3(new_n269_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n869_), .B1(new_n870_), .B2(new_n871_), .ZN(G1349gat));
  NAND3_X1  g671(.A1(new_n870_), .A2(new_n587_), .A3(new_n852_), .ZN(new_n873_));
  INV_X1    g672(.A(G183gat), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n614_), .A2(new_n301_), .ZN(new_n875_));
  AOI22_X1  g674(.A1(new_n873_), .A2(new_n874_), .B1(new_n868_), .B2(new_n875_), .ZN(G1350gat));
  NAND2_X1  g675(.A1(new_n868_), .A2(new_n647_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(G190gat), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n868_), .A2(new_n302_), .A3(new_n603_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1351gat));
  NOR3_X1   g679(.A1(new_n340_), .A2(new_n500_), .A3(new_n526_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT125), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n463_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n884_), .B1(new_n883_), .B2(new_n882_), .ZN(new_n885_));
  AND2_X1   g684(.A1(new_n801_), .A2(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(G197gat), .B1(new_n886_), .B2(new_n567_), .ZN(new_n887_));
  NAND4_X1  g686(.A1(new_n801_), .A2(G197gat), .A3(new_n567_), .A4(new_n885_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT126), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n888_), .A2(new_n889_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n887_), .A2(new_n890_), .A3(new_n891_), .ZN(G1352gat));
  NAND2_X1  g691(.A1(new_n886_), .A2(new_n269_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g693(.A1(new_n801_), .A2(new_n613_), .A3(new_n885_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n896_));
  AND2_X1   g695(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n895_), .A2(new_n896_), .A3(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n898_), .B1(new_n895_), .B2(new_n896_), .ZN(G1354gat));
  INV_X1    g698(.A(G218gat), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n886_), .A2(new_n900_), .A3(new_n603_), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n886_), .A2(new_n647_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n902_), .B2(new_n900_), .ZN(G1355gat));
endmodule


