//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 0 1 1 0 1 0 1 1 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 0 0 0 0 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n885_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n902_, new_n904_, new_n905_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n931_;
  XNOR2_X1  g000(.A(KEYINPUT25), .B(G183gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT26), .B(G190gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n206_), .A2(KEYINPUT24), .A3(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n204_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT92), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n206_), .A2(KEYINPUT24), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT23), .ZN(new_n213_));
  AND2_X1   g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n210_), .A2(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n213_), .B1(G183gat), .B2(G190gat), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n216_), .A2(new_n207_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT22), .B(G169gat), .ZN(new_n218_));
  XOR2_X1   g017(.A(new_n218_), .B(KEYINPUT93), .Z(new_n219_));
  OAI21_X1  g018(.A(new_n217_), .B1(new_n219_), .B2(G176gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n215_), .A2(new_n220_), .ZN(new_n221_));
  XOR2_X1   g020(.A(G197gat), .B(G204gat), .Z(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT21), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G197gat), .B(G204gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT21), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  OR2_X1    g025(.A1(G211gat), .A2(G218gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G211gat), .A2(G218gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(KEYINPUT86), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT86), .B1(new_n227_), .B2(new_n228_), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n223_), .B(new_n226_), .C1(new_n230_), .C2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n231_), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n233_), .A2(KEYINPUT21), .A3(new_n229_), .A4(new_n222_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT87), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n232_), .A2(KEYINPUT87), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n221_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(G190gat), .ZN(new_n241_));
  OR3_X1    g040(.A1(new_n241_), .A2(KEYINPUT80), .A3(KEYINPUT26), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT26), .B1(new_n241_), .B2(KEYINPUT80), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n242_), .A2(new_n202_), .A3(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n214_), .A2(new_n244_), .A3(new_n208_), .ZN(new_n245_));
  INV_X1    g044(.A(G176gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n218_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT81), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n217_), .A2(new_n249_), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n237_), .A2(new_n245_), .A3(new_n250_), .A4(new_n238_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n240_), .A2(new_n251_), .A3(KEYINPUT20), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G226gat), .A2(G233gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT19), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT20), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n250_), .A2(new_n245_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n256_), .B1(new_n239_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n254_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n215_), .A2(new_n237_), .A3(new_n238_), .A4(new_n220_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n258_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT94), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n258_), .A2(KEYINPUT94), .A3(new_n259_), .A4(new_n260_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n255_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G8gat), .B(G36gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT18), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(G64gat), .ZN(new_n268_));
  INV_X1    g067(.A(G92gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n265_), .B(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT27), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n258_), .A2(new_n260_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n254_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n276_), .B1(new_n254_), .B2(new_n252_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n271_), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n278_), .B(KEYINPUT27), .C1(new_n265_), .C2(new_n271_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n274_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT82), .ZN(new_n281_));
  OR2_X1    g080(.A1(G127gat), .A2(G134gat), .ZN(new_n282_));
  INV_X1    g081(.A(G113gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G127gat), .A2(G134gat), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(G120gat), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n283_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n286_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G127gat), .B(G134gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(G113gat), .ZN(new_n291_));
  AOI21_X1  g090(.A(G120gat), .B1(new_n291_), .B2(new_n285_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n281_), .B1(new_n289_), .B2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n287_), .B1(new_n286_), .B2(new_n288_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n291_), .A2(G120gat), .A3(new_n285_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(KEYINPUT82), .A3(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n293_), .A2(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n297_), .B(KEYINPUT31), .Z(new_n298_));
  INV_X1    g097(.A(KEYINPUT83), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G227gat), .A2(G233gat), .ZN(new_n300_));
  INV_X1    g099(.A(G15gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(G43gat), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G71gat), .B(G99gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT30), .ZN(new_n306_));
  AND3_X1   g105(.A1(new_n250_), .A2(new_n306_), .A3(new_n245_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n306_), .B1(new_n250_), .B2(new_n245_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n304_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NOR3_X1   g109(.A1(new_n307_), .A2(new_n308_), .A3(new_n304_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n299_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n311_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(new_n309_), .A3(KEYINPUT83), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n298_), .B1(new_n312_), .B2(new_n314_), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n314_), .A2(new_n298_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(G50gat), .ZN(new_n318_));
  NOR2_X1   g117(.A1(G141gat), .A2(G148gat), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G141gat), .A2(G148gat), .ZN(new_n321_));
  NOR2_X1   g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT84), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G155gat), .A2(G162gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT1), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n320_), .B(new_n321_), .C1(new_n323_), .C2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT84), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n322_), .B(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT3), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n319_), .B(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT2), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n321_), .B(new_n331_), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n328_), .B(new_n324_), .C1(new_n330_), .C2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n326_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT85), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT29), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n326_), .A2(new_n333_), .A3(KEYINPUT85), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n336_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT28), .ZN(new_n340_));
  INV_X1    g139(.A(G22gat), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT28), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n336_), .A2(new_n342_), .A3(new_n337_), .A4(new_n338_), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n340_), .A2(new_n341_), .A3(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n341_), .B1(new_n340_), .B2(new_n343_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n318_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n340_), .A2(new_n343_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(G22gat), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n340_), .A2(new_n341_), .A3(new_n343_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(G50gat), .A3(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n346_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT89), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n237_), .A2(new_n238_), .B1(KEYINPUT29), .B2(new_n334_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G228gat), .A2(G233gat), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n337_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n232_), .A2(KEYINPUT87), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT87), .B1(new_n232_), .B2(new_n234_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n354_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  OAI22_X1  g157(.A1(new_n353_), .A2(new_n354_), .B1(new_n355_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT88), .ZN(new_n360_));
  XOR2_X1   g159(.A(G78gat), .B(G106gat), .Z(new_n361_));
  NAND3_X1  g160(.A1(new_n359_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n326_), .A2(new_n333_), .ZN(new_n363_));
  OAI22_X1  g162(.A1(new_n356_), .A2(new_n357_), .B1(new_n363_), .B2(new_n337_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n364_), .A2(G228gat), .A3(G233gat), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n326_), .A2(new_n333_), .A3(KEYINPUT85), .ZN(new_n366_));
  AOI21_X1  g165(.A(KEYINPUT85), .B1(new_n326_), .B2(new_n333_), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT29), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n368_), .A2(new_n354_), .A3(new_n239_), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n361_), .A2(new_n360_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n361_), .A2(new_n360_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n365_), .A2(new_n369_), .A3(new_n370_), .A4(new_n371_), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n362_), .A2(new_n372_), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n351_), .A2(new_n352_), .A3(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n352_), .B1(new_n351_), .B2(new_n373_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n361_), .A2(KEYINPUT90), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n359_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n365_), .A2(new_n369_), .A3(new_n377_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n346_), .A2(new_n350_), .A3(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT91), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n346_), .A2(new_n350_), .A3(new_n381_), .A4(KEYINPUT91), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n317_), .B1(new_n376_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n351_), .A2(new_n373_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT89), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n351_), .A2(new_n352_), .A3(new_n373_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n317_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n384_), .A2(new_n385_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n391_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n280_), .B1(new_n387_), .B2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n297_), .B1(new_n367_), .B2(new_n366_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n363_), .A2(new_n295_), .A3(new_n294_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n396_), .A2(KEYINPUT4), .A3(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT95), .ZN(new_n399_));
  OR2_X1    g198(.A1(new_n396_), .A2(KEYINPUT4), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT95), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n396_), .A2(new_n401_), .A3(KEYINPUT4), .A4(new_n397_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n399_), .A2(new_n400_), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G225gat), .A2(G233gat), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(KEYINPUT96), .B(KEYINPUT0), .Z(new_n407_));
  XNOR2_X1  g206(.A(G1gat), .B(G29gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G57gat), .B(G85gat), .ZN(new_n410_));
  XOR2_X1   g209(.A(new_n409_), .B(new_n410_), .Z(new_n411_));
  AND2_X1   g210(.A1(new_n396_), .A2(new_n397_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n412_), .A2(new_n405_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n406_), .A2(new_n411_), .A3(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT99), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n406_), .A2(new_n414_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n411_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n413_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n421_), .A2(KEYINPUT99), .A3(new_n411_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n417_), .A2(new_n420_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n393_), .B1(new_n375_), .B2(new_n374_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n270_), .A2(KEYINPUT32), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n277_), .A2(new_n426_), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n265_), .A2(new_n426_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n423_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n412_), .A2(new_n405_), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT97), .B1(new_n430_), .B2(new_n411_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT98), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n399_), .A2(new_n404_), .A3(new_n400_), .A4(new_n402_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n431_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n430_), .A2(KEYINPUT97), .A3(new_n411_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n434_), .B(new_n435_), .C1(new_n432_), .C2(new_n433_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n265_), .B(new_n270_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT33), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n438_), .B1(new_n421_), .B2(new_n411_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n418_), .A2(KEYINPUT33), .A3(new_n419_), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n436_), .A2(new_n437_), .A3(new_n439_), .A4(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n425_), .B1(new_n429_), .B2(new_n441_), .ZN(new_n442_));
  AOI22_X1  g241(.A1(new_n395_), .A2(new_n424_), .B1(new_n442_), .B2(new_n317_), .ZN(new_n443_));
  XOR2_X1   g242(.A(G57gat), .B(G64gat), .Z(new_n444_));
  INV_X1    g243(.A(KEYINPUT11), .ZN(new_n445_));
  AOI22_X1  g244(.A1(new_n444_), .A2(new_n445_), .B1(G71gat), .B2(G78gat), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT70), .B1(new_n444_), .B2(new_n445_), .ZN(new_n447_));
  OR2_X1    g246(.A1(G71gat), .A2(G78gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G57gat), .B(G64gat), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT70), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n449_), .A2(new_n450_), .A3(KEYINPUT11), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n446_), .A2(new_n447_), .A3(new_n448_), .A4(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G71gat), .A2(G78gat), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n448_), .B(new_n453_), .C1(new_n449_), .C2(KEYINPUT11), .ZN(new_n454_));
  INV_X1    g253(.A(new_n451_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n450_), .B1(new_n449_), .B2(KEYINPUT11), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n454_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n452_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n459_), .A2(G231gat), .A3(G233gat), .ZN(new_n460_));
  INV_X1    g259(.A(G231gat), .ZN(new_n461_));
  INV_X1    g260(.A(G233gat), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n458_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n460_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G1gat), .B(G8gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT75), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n301_), .A2(new_n341_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G15gat), .A2(G22gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G1gat), .A2(G8gat), .ZN(new_n469_));
  AOI22_X1  g268(.A1(new_n467_), .A2(new_n468_), .B1(KEYINPUT14), .B2(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(new_n466_), .B(new_n470_), .Z(new_n471_));
  NAND2_X1  g270(.A1(new_n464_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G183gat), .B(G211gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G127gat), .B(G155gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n477_), .A2(KEYINPUT17), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n466_), .B(new_n470_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n460_), .A2(new_n463_), .A3(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n472_), .A2(new_n478_), .A3(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n477_), .A2(KEYINPUT17), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT77), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n481_), .B(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G232gat), .A2(G233gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT34), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT35), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G29gat), .B(G36gat), .ZN(new_n488_));
  INV_X1    g287(.A(G43gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(G50gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n488_), .B(G43gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(new_n318_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(G99gat), .ZN(new_n496_));
  INV_X1    g295(.A(G106gat), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT67), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n496_), .B(new_n497_), .C1(new_n498_), .C2(KEYINPUT7), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT7), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n500_), .B(KEYINPUT67), .C1(G99gat), .C2(G106gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n499_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT68), .ZN(new_n503_));
  AND3_X1   g302(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n504_));
  AOI21_X1  g303(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n503_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G99gat), .A2(G106gat), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT6), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n509_), .A2(KEYINPUT68), .A3(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n502_), .A2(new_n506_), .A3(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G85gat), .B(G92gat), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT66), .B1(new_n504_), .B2(new_n505_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT66), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n509_), .A2(new_n517_), .A3(new_n510_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n502_), .A2(new_n516_), .A3(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n513_), .A2(KEYINPUT8), .ZN(new_n520_));
  AOI22_X1  g319(.A1(new_n515_), .A2(KEYINPUT8), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  XOR2_X1   g320(.A(KEYINPUT10), .B(G99gat), .Z(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(new_n497_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n269_), .A2(KEYINPUT65), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT65), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(G92gat), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n525_), .A2(new_n527_), .A3(G85gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n529_));
  INV_X1    g328(.A(G85gat), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n530_), .A2(KEYINPUT9), .ZN(new_n531_));
  AOI22_X1  g330(.A1(new_n528_), .A2(new_n529_), .B1(new_n513_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n516_), .A2(new_n518_), .ZN(new_n533_));
  NOR3_X1   g332(.A1(new_n524_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT69), .B1(new_n521_), .B2(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n532_), .A2(new_n533_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(new_n523_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT69), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT8), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n539_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n519_), .A2(new_n520_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n537_), .B(new_n538_), .C1(new_n540_), .C2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n535_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT15), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n492_), .A2(new_n318_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n490_), .A2(G50gat), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n545_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n491_), .A2(new_n493_), .A3(KEYINPUT15), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n515_), .A2(KEYINPUT8), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(new_n541_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n548_), .A2(new_n549_), .B1(new_n551_), .B2(new_n537_), .ZN(new_n552_));
  AOI22_X1  g351(.A1(new_n495_), .A2(new_n544_), .B1(new_n552_), .B2(KEYINPUT73), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n552_), .A2(KEYINPUT73), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n487_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT36), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G190gat), .B(G218gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT74), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(G134gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(G162gat), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n544_), .A2(new_n495_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n552_), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n486_), .B(KEYINPUT35), .Z(new_n564_));
  NAND3_X1  g363(.A1(new_n562_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n556_), .A2(new_n557_), .A3(new_n561_), .A4(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n561_), .A2(new_n557_), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n561_), .A2(new_n557_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n565_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n567_), .B(new_n568_), .C1(new_n555_), .C2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n566_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT37), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n566_), .A2(KEYINPUT37), .A3(new_n570_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NOR3_X1   g374(.A1(new_n443_), .A2(new_n484_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT78), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n548_), .A2(new_n549_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(new_n479_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G229gat), .A2(G233gat), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n471_), .A2(new_n495_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n579_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n479_), .A2(new_n494_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n580_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n577_), .B1(new_n582_), .B2(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(KEYINPUT78), .B1(new_n584_), .B2(new_n585_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G113gat), .B(G141gat), .ZN(new_n590_));
  INV_X1    g389(.A(G169gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(G197gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT79), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n589_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n595_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n587_), .A2(new_n598_), .A3(new_n588_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n597_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n544_), .A2(new_n458_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n535_), .A2(new_n459_), .A3(new_n543_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G230gat), .A2(G233gat), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT12), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n603_), .A2(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n458_), .B1(new_n551_), .B2(new_n537_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT12), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n609_), .A2(new_n602_), .A3(new_n611_), .A4(new_n605_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n607_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G120gat), .B(G148gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G176gat), .B(G204gat), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n616_), .B(new_n617_), .Z(new_n618_));
  NAND2_X1  g417(.A1(new_n613_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n618_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n607_), .A2(new_n612_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT13), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n619_), .A2(KEYINPUT13), .A3(new_n621_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT72), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n576_), .A2(new_n601_), .A3(new_n628_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n629_), .A2(G1gat), .A3(new_n424_), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n630_), .A2(KEYINPUT38), .ZN(new_n631_));
  INV_X1    g430(.A(new_n571_), .ZN(new_n632_));
  OAI21_X1  g431(.A(KEYINPUT100), .B1(new_n443_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n484_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n274_), .A2(new_n279_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n425_), .A2(new_n317_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n392_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n424_), .B(new_n635_), .C1(new_n636_), .C2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n429_), .A2(new_n441_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n425_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n639_), .A2(new_n317_), .A3(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n638_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT100), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n642_), .A2(new_n643_), .A3(new_n571_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n601_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n645_), .A2(new_n626_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n633_), .A2(new_n634_), .A3(new_n644_), .A4(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G1gat), .B1(new_n647_), .B2(new_n424_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n630_), .A2(KEYINPUT38), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n631_), .A2(new_n648_), .A3(new_n649_), .ZN(G1324gat));
  INV_X1    g449(.A(KEYINPUT40), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT101), .ZN(new_n652_));
  OAI21_X1  g451(.A(G8gat), .B1(new_n647_), .B2(new_n635_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(KEYINPUT39), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT39), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n655_), .B(G8gat), .C1(new_n647_), .C2(new_n635_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n629_), .A2(G8gat), .A3(new_n635_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n652_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n660_));
  AOI211_X1 g459(.A(KEYINPUT101), .B(new_n658_), .C1(new_n654_), .C2(new_n656_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n651_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n643_), .B1(new_n642_), .B2(new_n571_), .ZN(new_n663_));
  AOI211_X1 g462(.A(KEYINPUT100), .B(new_n632_), .C1(new_n638_), .C2(new_n641_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n665_), .A2(new_n634_), .A3(new_n280_), .A4(new_n646_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n655_), .B1(new_n666_), .B2(G8gat), .ZN(new_n667_));
  INV_X1    g466(.A(new_n656_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n659_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT101), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n657_), .A2(new_n652_), .A3(new_n659_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n670_), .A2(KEYINPUT40), .A3(new_n671_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n662_), .A2(new_n672_), .ZN(G1325gat));
  OAI21_X1  g472(.A(G15gat), .B1(new_n647_), .B2(new_n317_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT41), .Z(new_n675_));
  INV_X1    g474(.A(new_n629_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n676_), .A2(new_n301_), .A3(new_n392_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(G1326gat));
  OAI21_X1  g477(.A(G22gat), .B1(new_n647_), .B2(new_n640_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT42), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n676_), .A2(new_n341_), .A3(new_n425_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1327gat));
  AND4_X1   g481(.A1(new_n484_), .A2(new_n642_), .A3(new_n632_), .A4(new_n646_), .ZN(new_n683_));
  AOI21_X1  g482(.A(G29gat), .B1(new_n683_), .B2(new_n423_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n685_));
  INV_X1    g484(.A(new_n575_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n685_), .B1(new_n443_), .B2(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n642_), .A2(KEYINPUT43), .A3(new_n575_), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n687_), .A2(new_n484_), .A3(new_n646_), .A4(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(KEYINPUT102), .A3(KEYINPUT44), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(KEYINPUT44), .B1(new_n689_), .B2(KEYINPUT102), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n693_), .A2(new_n424_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n684_), .B1(new_n694_), .B2(G29gat), .ZN(G1328gat));
  OAI21_X1  g494(.A(G36gat), .B1(new_n693_), .B2(new_n635_), .ZN(new_n696_));
  OR2_X1    g495(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n697_));
  INV_X1    g496(.A(G36gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n683_), .A2(new_n698_), .A3(new_n280_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(KEYINPUT103), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n683_), .A2(new_n701_), .A3(new_n698_), .A4(new_n280_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT45), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT45), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n700_), .A2(new_n705_), .A3(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n696_), .A2(new_n697_), .A3(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(KEYINPUT105), .B1(KEYINPUT104), .B2(KEYINPUT46), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT106), .Z(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n708_), .A2(new_n711_), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n696_), .A2(new_n710_), .A3(new_n697_), .A4(new_n707_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1329gat));
  OAI21_X1  g513(.A(new_n392_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n317_), .A2(G43gat), .ZN(new_n716_));
  AOI22_X1  g515(.A1(new_n715_), .A2(G43gat), .B1(new_n683_), .B2(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n717_), .B(new_n719_), .ZN(G1330gat));
  OAI21_X1  g519(.A(G50gat), .B1(new_n693_), .B2(new_n640_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n683_), .A2(new_n318_), .A3(new_n425_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1331gat));
  NOR3_X1   g522(.A1(new_n596_), .A2(new_n484_), .A3(new_n599_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n665_), .A2(new_n627_), .A3(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(G57gat), .B1(new_n725_), .B2(new_n424_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n626_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n727_), .A2(new_n601_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n576_), .A2(new_n728_), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n424_), .A2(G57gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n726_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT108), .ZN(G1332gat));
  OAI21_X1  g531(.A(G64gat), .B1(new_n725_), .B2(new_n635_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT48), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n635_), .A2(G64gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(new_n729_), .B2(new_n735_), .ZN(G1333gat));
  OAI21_X1  g535(.A(G71gat), .B1(new_n725_), .B2(new_n317_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT49), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n317_), .A2(G71gat), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n729_), .B2(new_n739_), .ZN(G1334gat));
  OAI21_X1  g539(.A(G78gat), .B1(new_n725_), .B2(new_n640_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT50), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n640_), .A2(G78gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n742_), .B1(new_n729_), .B2(new_n743_), .ZN(G1335gat));
  NOR3_X1   g543(.A1(new_n443_), .A2(new_n634_), .A3(new_n571_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n745_), .A2(new_n645_), .A3(new_n627_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n530_), .B1(new_n746_), .B2(new_n424_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n687_), .A2(new_n484_), .A3(new_n688_), .A4(new_n728_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n423_), .A2(G85gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n747_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(G1336gat));
  OAI21_X1  g550(.A(new_n269_), .B1(new_n746_), .B2(new_n635_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n280_), .A2(new_n525_), .A3(new_n527_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n752_), .B1(new_n748_), .B2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(G1337gat));
  NAND2_X1  g554(.A1(new_n392_), .A2(new_n522_), .ZN(new_n756_));
  OR2_X1    g555(.A1(new_n746_), .A2(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(G99gat), .B1(new_n748_), .B2(new_n317_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT109), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT51), .ZN(G1338gat));
  NOR3_X1   g560(.A1(new_n746_), .A2(G106gat), .A3(new_n640_), .ZN(new_n762_));
  XOR2_X1   g561(.A(new_n762_), .B(KEYINPUT110), .Z(new_n763_));
  OAI21_X1  g562(.A(G106gat), .B1(new_n748_), .B2(new_n640_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765_));
  OR2_X1    g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n765_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n763_), .A2(new_n766_), .A3(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(KEYINPUT53), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT53), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n763_), .A2(new_n770_), .A3(new_n766_), .A4(new_n767_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(G1339gat));
  NAND3_X1  g571(.A1(new_n724_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT111), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT111), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n724_), .A2(new_n624_), .A3(new_n775_), .A4(new_n625_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n686_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n777_), .A2(KEYINPUT113), .A3(new_n686_), .ZN(new_n781_));
  XOR2_X1   g580(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n782_));
  NAND3_X1  g581(.A1(new_n780_), .A2(new_n781_), .A3(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n782_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT113), .B1(new_n777_), .B2(new_n686_), .ZN(new_n785_));
  AOI211_X1 g584(.A(new_n779_), .B(new_n575_), .C1(new_n774_), .C2(new_n776_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n784_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n783_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n621_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n597_), .B2(new_n600_), .ZN(new_n790_));
  AOI22_X1  g589(.A1(new_n544_), .A2(new_n458_), .B1(KEYINPUT12), .B2(new_n610_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n605_), .B1(new_n791_), .B2(new_n609_), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n791_), .A2(new_n605_), .A3(new_n609_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n793_), .B2(KEYINPUT55), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT55), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n612_), .A2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT114), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n612_), .A2(new_n798_), .A3(new_n795_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n794_), .A2(new_n797_), .A3(new_n799_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n800_), .A2(KEYINPUT56), .A3(new_n618_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT56), .B1(new_n800_), .B2(new_n618_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n790_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT115), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n579_), .A2(new_n585_), .A3(new_n581_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n585_), .B1(new_n581_), .B2(new_n583_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n594_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n807_), .B1(new_n589_), .B2(new_n594_), .ZN(new_n808_));
  XOR2_X1   g607(.A(new_n808_), .B(KEYINPUT116), .Z(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n622_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n811_), .B(new_n790_), .C1(new_n801_), .C2(new_n802_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n804_), .A2(new_n810_), .A3(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n571_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT56), .ZN(new_n817_));
  INV_X1    g616(.A(new_n799_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n609_), .A2(new_n602_), .A3(new_n611_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n606_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n791_), .A2(KEYINPUT55), .A3(new_n605_), .A4(new_n609_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n798_), .B1(new_n612_), .B2(new_n795_), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n818_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n817_), .B1(new_n824_), .B2(new_n620_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n800_), .A2(KEYINPUT56), .A3(new_n618_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n825_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n789_), .B1(new_n802_), .B2(KEYINPUT117), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n829_), .A3(new_n809_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(KEYINPUT118), .A2(KEYINPUT58), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n831_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n828_), .A2(new_n829_), .A3(new_n809_), .A4(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n832_), .A2(new_n575_), .A3(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n813_), .A2(KEYINPUT57), .A3(new_n571_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n816_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n788_), .B1(new_n837_), .B2(new_n484_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n280_), .A2(new_n424_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n636_), .ZN(new_n840_));
  XOR2_X1   g639(.A(new_n840_), .B(KEYINPUT119), .Z(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n838_), .A2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(G113gat), .B1(new_n843_), .B2(new_n601_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n788_), .ZN(new_n845_));
  AND3_X1   g644(.A1(new_n813_), .A2(KEYINPUT57), .A3(new_n571_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n832_), .A2(new_n575_), .A3(new_n834_), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT57), .B1(new_n813_), .B2(new_n571_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n846_), .A2(new_n847_), .A3(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n845_), .B1(new_n849_), .B2(new_n634_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n851_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n850_), .A2(new_n841_), .A3(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(KEYINPUT120), .B1(new_n841_), .B2(KEYINPUT121), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n853_), .B1(new_n838_), .B2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n645_), .B1(new_n855_), .B2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n844_), .B1(new_n858_), .B2(G113gat), .ZN(G1340gat));
  NAND2_X1  g658(.A1(new_n855_), .A2(new_n857_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n727_), .A2(G120gat), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n843_), .B1(KEYINPUT60), .B2(new_n861_), .ZN(new_n862_));
  AND3_X1   g661(.A1(new_n860_), .A2(new_n862_), .A3(new_n627_), .ZN(new_n863_));
  OAI22_X1  g662(.A1(new_n863_), .A2(new_n287_), .B1(KEYINPUT60), .B2(new_n862_), .ZN(G1341gat));
  AOI21_X1  g663(.A(G127gat), .B1(new_n843_), .B2(new_n634_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n866_));
  OR2_X1    g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n866_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n860_), .A2(G127gat), .A3(new_n634_), .ZN(new_n869_));
  AND3_X1   g668(.A1(new_n867_), .A2(new_n868_), .A3(new_n869_), .ZN(G1342gat));
  INV_X1    g669(.A(G134gat), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n843_), .A2(new_n871_), .A3(new_n632_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n686_), .B1(new_n855_), .B2(new_n857_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(new_n871_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(KEYINPUT123), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT123), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n876_), .B(new_n872_), .C1(new_n873_), .C2(new_n871_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(G1343gat));
  NAND2_X1  g677(.A1(new_n839_), .A2(new_n637_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(KEYINPUT124), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n838_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n601_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n627_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(KEYINPUT125), .B(G148gat), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n884_), .B(new_n885_), .ZN(G1345gat));
  NAND2_X1  g685(.A1(new_n881_), .A2(new_n634_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(KEYINPUT61), .B(G155gat), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1346gat));
  AOI21_X1  g688(.A(G162gat), .B1(new_n881_), .B2(new_n632_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n575_), .A2(G162gat), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n890_), .B1(new_n881_), .B2(new_n891_), .ZN(G1347gat));
  NOR4_X1   g691(.A1(new_n838_), .A2(new_n423_), .A3(new_n394_), .A4(new_n635_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n219_), .ZN(new_n894_));
  AND3_X1   g693(.A1(new_n893_), .A2(new_n894_), .A3(new_n601_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n591_), .B1(new_n893_), .B2(new_n601_), .ZN(new_n896_));
  OAI21_X1  g695(.A(KEYINPUT62), .B1(new_n895_), .B2(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n897_), .B1(KEYINPUT62), .B2(new_n896_), .ZN(G1348gat));
  AOI21_X1  g697(.A(G176gat), .B1(new_n893_), .B2(new_n626_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n628_), .A2(new_n246_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n893_), .B2(new_n900_), .ZN(G1349gat));
  NAND2_X1  g700(.A1(new_n893_), .A2(new_n634_), .ZN(new_n902_));
  MUX2_X1   g701(.A(new_n202_), .B(G183gat), .S(new_n902_), .Z(G1350gat));
  NAND3_X1  g702(.A1(new_n893_), .A2(new_n632_), .A3(new_n203_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n893_), .A2(new_n575_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n905_), .B2(new_n241_), .ZN(G1351gat));
  NAND4_X1  g705(.A1(new_n850_), .A2(new_n424_), .A3(new_n637_), .A4(new_n280_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT126), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n838_), .A2(new_n423_), .ZN(new_n910_));
  NAND4_X1  g709(.A1(new_n910_), .A2(KEYINPUT126), .A3(new_n637_), .A4(new_n280_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(G197gat), .B1(new_n912_), .B2(new_n601_), .ZN(new_n913_));
  AOI211_X1 g712(.A(new_n593_), .B(new_n645_), .C1(new_n909_), .C2(new_n911_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1352gat));
  NOR3_X1   g714(.A1(new_n838_), .A2(new_n423_), .A3(new_n635_), .ZN(new_n916_));
  AOI21_X1  g715(.A(KEYINPUT126), .B1(new_n916_), .B2(new_n637_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n907_), .A2(new_n908_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n627_), .B1(new_n917_), .B2(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(G204gat), .ZN(new_n920_));
  INV_X1    g719(.A(G204gat), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n912_), .A2(new_n921_), .A3(new_n627_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n920_), .A2(new_n922_), .ZN(G1353gat));
  OR2_X1    g722(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n924_), .B1(new_n912_), .B2(new_n634_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(KEYINPUT63), .B(G211gat), .ZN(new_n926_));
  AOI211_X1 g725(.A(new_n484_), .B(new_n926_), .C1(new_n909_), .C2(new_n911_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n925_), .A2(new_n927_), .ZN(G1354gat));
  AOI21_X1  g727(.A(G218gat), .B1(new_n912_), .B2(new_n632_), .ZN(new_n929_));
  INV_X1    g728(.A(G218gat), .ZN(new_n930_));
  AOI211_X1 g729(.A(new_n930_), .B(new_n686_), .C1(new_n909_), .C2(new_n911_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n929_), .A2(new_n931_), .ZN(G1355gat));
endmodule


