//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 0 0 0 1 1 0 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n836_, new_n838_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n848_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n892_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_;
  XNOR2_X1  g000(.A(KEYINPUT26), .B(G190gat), .ZN(new_n202_));
  INV_X1    g001(.A(G183gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT25), .B1(new_n203_), .B2(KEYINPUT78), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n203_), .A2(KEYINPUT25), .ZN(new_n205_));
  OAI211_X1 g004(.A(new_n202_), .B(new_n204_), .C1(new_n205_), .C2(KEYINPUT78), .ZN(new_n206_));
  XOR2_X1   g005(.A(G169gat), .B(G176gat), .Z(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT24), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n209_));
  INV_X1    g008(.A(G190gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n209_), .B1(new_n203_), .B2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n212_));
  AND2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT24), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n206_), .A2(new_n208_), .A3(new_n213_), .A4(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G176gat), .ZN(new_n218_));
  INV_X1    g017(.A(G169gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT22), .B1(new_n219_), .B2(KEYINPUT79), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n219_), .A2(KEYINPUT22), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n218_), .B(new_n220_), .C1(new_n221_), .C2(KEYINPUT79), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n211_), .B(new_n212_), .C1(G183gat), .C2(G190gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n217_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT30), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G15gat), .B(G43gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(KEYINPUT80), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(G99gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G227gat), .A2(G233gat), .ZN(new_n231_));
  INV_X1    g030(.A(G71gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n230_), .B(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n227_), .B1(new_n234_), .B2(KEYINPUT81), .ZN(new_n235_));
  INV_X1    g034(.A(new_n233_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n230_), .B(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT81), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n235_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n237_), .A2(new_n238_), .A3(new_n227_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n240_), .A2(KEYINPUT83), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT31), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT31), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n240_), .A2(KEYINPUT83), .A3(new_n244_), .A4(new_n241_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G127gat), .B(G134gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT82), .ZN(new_n248_));
  XOR2_X1   g047(.A(G113gat), .B(G120gat), .Z(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n246_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n250_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n243_), .A2(new_n252_), .A3(new_n245_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G225gat), .A2(G233gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G155gat), .B(G162gat), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n257_), .A2(KEYINPUT1), .ZN(new_n258_));
  INV_X1    g057(.A(G141gat), .ZN(new_n259_));
  INV_X1    g058(.A(G148gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G141gat), .A2(G148gat), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n261_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n258_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n263_), .B(KEYINPUT2), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT84), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT3), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n261_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n259_), .B(new_n260_), .C1(new_n267_), .C2(new_n268_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n266_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  OR2_X1    g072(.A1(new_n273_), .A2(KEYINPUT85), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n257_), .B1(new_n273_), .B2(KEYINPUT85), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n265_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT92), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(new_n278_), .A3(new_n252_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n280_), .B1(new_n276_), .B2(new_n250_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n277_), .A2(new_n278_), .A3(new_n280_), .A4(new_n252_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n256_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  XOR2_X1   g084(.A(G1gat), .B(G29gat), .Z(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT93), .B(G85gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT0), .B(G57gat), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n288_), .B(new_n289_), .Z(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n276_), .B(new_n250_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(new_n256_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n285_), .A2(new_n291_), .A3(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n293_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n290_), .B1(new_n284_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT97), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n294_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n285_), .A2(KEYINPUT97), .A3(new_n291_), .A4(new_n293_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n298_), .A2(KEYINPUT98), .A3(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(KEYINPUT98), .B1(new_n298_), .B2(new_n299_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n224_), .B(KEYINPUT90), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT22), .B(G169gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT91), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n223_), .B(new_n303_), .C1(new_n305_), .C2(G176gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n214_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n213_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT89), .ZN(new_n310_));
  INV_X1    g109(.A(new_n307_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT25), .B(G183gat), .ZN(new_n312_));
  AOI22_X1  g111(.A1(new_n311_), .A2(new_n207_), .B1(new_n202_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n310_), .A2(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n309_), .A2(KEYINPUT89), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n306_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(G197gat), .A2(G204gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT86), .B(G204gat), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n317_), .B1(new_n318_), .B2(G197gat), .ZN(new_n319_));
  OR2_X1    g118(.A1(new_n319_), .A2(KEYINPUT21), .ZN(new_n320_));
  XOR2_X1   g119(.A(G211gat), .B(G218gat), .Z(new_n321_));
  OR2_X1    g120(.A1(new_n318_), .A2(G197gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT21), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n323_), .B1(G197gat), .B2(G204gat), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n321_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n320_), .A2(new_n325_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n321_), .A2(KEYINPUT21), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(new_n319_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n316_), .A2(new_n329_), .ZN(new_n330_));
  AOI22_X1  g129(.A1(new_n320_), .A2(new_n325_), .B1(new_n319_), .B2(new_n327_), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT20), .B1(new_n331_), .B2(new_n226_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G226gat), .A2(G233gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT19), .ZN(new_n334_));
  OR3_X1    g133(.A1(new_n330_), .A2(new_n332_), .A3(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n316_), .A2(new_n329_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n331_), .A2(new_n226_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(KEYINPUT20), .A3(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(new_n334_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n335_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G8gat), .B(G36gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT18), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G64gat), .B(G92gat), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n342_), .B(new_n343_), .Z(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n340_), .A2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n335_), .A2(new_n339_), .A3(new_n344_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n348_), .A2(KEYINPUT27), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT27), .ZN(new_n350_));
  INV_X1    g149(.A(new_n347_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n334_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n352_), .B(KEYINPUT96), .C1(new_n334_), .C2(new_n338_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT96), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n354_), .B(new_n334_), .C1(new_n330_), .C2(new_n332_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n353_), .A2(new_n345_), .A3(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n351_), .B1(new_n356_), .B2(KEYINPUT99), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT99), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n353_), .A2(new_n358_), .A3(new_n345_), .A4(new_n355_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n350_), .B1(new_n357_), .B2(new_n359_), .ZN(new_n360_));
  OAI22_X1  g159(.A1(new_n301_), .A2(new_n302_), .B1(new_n349_), .B2(new_n360_), .ZN(new_n361_));
  NOR3_X1   g160(.A1(new_n277_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT28), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT29), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n363_), .B1(new_n276_), .B2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G22gat), .B(G50gat), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  OR3_X1    g166(.A1(new_n362_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n367_), .B1(new_n362_), .B2(new_n365_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(KEYINPUT87), .A3(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n331_), .B1(new_n277_), .B2(KEYINPUT29), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G228gat), .A2(G233gat), .ZN(new_n372_));
  INV_X1    g171(.A(G78gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(G106gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n371_), .B(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n370_), .A2(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT87), .B1(new_n368_), .B2(new_n369_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n370_), .A2(new_n378_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n255_), .B1(new_n361_), .B2(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n291_), .B1(new_n292_), .B2(new_n256_), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n282_), .A2(new_n283_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n385_), .B1(new_n386_), .B2(new_n256_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n348_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT94), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n296_), .A2(new_n389_), .A3(KEYINPUT33), .ZN(new_n390_));
  AOI21_X1  g189(.A(KEYINPUT33), .B1(new_n296_), .B2(new_n389_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n388_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT95), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n383_), .ZN(new_n395_));
  OAI211_X1 g194(.A(KEYINPUT95), .B(new_n388_), .C1(new_n390_), .C2(new_n391_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n353_), .A2(new_n355_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n344_), .A2(KEYINPUT32), .ZN(new_n398_));
  MUX2_X1   g197(.A(new_n397_), .B(new_n340_), .S(new_n398_), .Z(new_n399_));
  NAND3_X1  g198(.A1(new_n399_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .A4(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n356_), .A2(KEYINPUT99), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(new_n347_), .A3(new_n359_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n349_), .B1(new_n403_), .B2(KEYINPUT27), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT100), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT100), .B1(new_n360_), .B2(new_n349_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n383_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n302_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n254_), .B1(new_n300_), .B2(new_n409_), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n384_), .A2(new_n401_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT70), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G230gat), .A2(G233gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT68), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n232_), .A2(KEYINPUT67), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT67), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(G71gat), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n416_), .A2(new_n418_), .A3(new_n373_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n373_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT11), .ZN(new_n422_));
  INV_X1    g221(.A(G64gat), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n423_), .A2(G57gat), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(G57gat), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n422_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n415_), .B1(new_n421_), .B2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n417_), .A2(G71gat), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n232_), .A2(KEYINPUT67), .ZN(new_n429_));
  OAI21_X1  g228(.A(G78gat), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n416_), .A2(new_n418_), .A3(new_n373_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n426_), .A2(new_n430_), .A3(new_n415_), .A4(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n424_), .A2(new_n425_), .ZN(new_n434_));
  OAI22_X1  g233(.A1(new_n427_), .A2(new_n433_), .B1(new_n422_), .B2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n426_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT68), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n434_), .A2(new_n422_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(new_n432_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n435_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT64), .ZN(new_n441_));
  OR2_X1    g240(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n441_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n442_), .A2(new_n441_), .A3(new_n443_), .ZN(new_n446_));
  AOI21_X1  g245(.A(G106gat), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G99gat), .A2(G106gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT6), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT6), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n450_), .A2(G99gat), .A3(G106gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n449_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G85gat), .A2(G92gat), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT9), .ZN(new_n454_));
  OR3_X1    g253(.A1(new_n453_), .A2(new_n454_), .A3(KEYINPUT65), .ZN(new_n455_));
  OR2_X1    g254(.A1(G85gat), .A2(G92gat), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n454_), .B1(new_n456_), .B2(new_n453_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n453_), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT65), .B1(new_n458_), .B2(KEYINPUT9), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n452_), .B(new_n455_), .C1(new_n457_), .C2(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n447_), .A2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n450_), .B1(G99gat), .B2(G106gat), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n448_), .A2(KEYINPUT6), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT66), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT66), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n449_), .A2(new_n451_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT7), .ZN(new_n467_));
  INV_X1    g266(.A(G99gat), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n467_), .A2(new_n468_), .A3(new_n375_), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n464_), .A2(new_n466_), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n456_), .A2(new_n453_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT8), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n471_), .A2(new_n452_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT8), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(new_n478_), .A3(new_n474_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n461_), .B1(new_n476_), .B2(new_n479_), .ZN(new_n480_));
  AOI211_X1 g279(.A(new_n412_), .B(new_n414_), .C1(new_n440_), .C2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n446_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n375_), .B1(new_n482_), .B2(new_n444_), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n457_), .A2(new_n459_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n483_), .A2(new_n484_), .A3(new_n452_), .A4(new_n455_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n469_), .A2(new_n470_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n486_), .B1(KEYINPUT66), .B2(new_n452_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n473_), .B1(new_n487_), .B2(new_n466_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n479_), .B1(new_n488_), .B2(new_n478_), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n437_), .A2(new_n438_), .A3(new_n432_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n438_), .B1(new_n437_), .B2(new_n432_), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n485_), .B(new_n489_), .C1(new_n490_), .C2(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT70), .B1(new_n492_), .B2(new_n413_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n478_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n494_));
  AOI211_X1 g293(.A(KEYINPUT8), .B(new_n473_), .C1(new_n471_), .C2(new_n452_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n485_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n496_), .A2(new_n439_), .A3(new_n435_), .ZN(new_n497_));
  AOI21_X1  g296(.A(KEYINPUT12), .B1(new_n497_), .B2(KEYINPUT69), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT69), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT12), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n490_), .A2(new_n491_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n502_), .B1(new_n503_), .B2(new_n496_), .ZN(new_n504_));
  OAI22_X1  g303(.A1(new_n481_), .A2(new_n493_), .B1(new_n498_), .B2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n413_), .B1(new_n492_), .B2(new_n497_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  XOR2_X1   g306(.A(G120gat), .B(G148gat), .Z(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G176gat), .B(G204gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n505_), .A2(new_n507_), .A3(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT72), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n496_), .B1(new_n439_), .B2(new_n435_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n412_), .B1(new_n516_), .B2(new_n414_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n492_), .A2(KEYINPUT70), .A3(new_n413_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n497_), .A2(new_n501_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n499_), .B1(new_n503_), .B2(new_n496_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n520_), .B1(new_n521_), .B2(KEYINPUT12), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n506_), .B1(new_n519_), .B2(new_n522_), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n523_), .A2(new_n513_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n515_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(KEYINPUT73), .B(KEYINPUT13), .Z(new_n528_));
  OAI21_X1  g327(.A(new_n527_), .B1(new_n525_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(KEYINPUT76), .B(G1gat), .Z(new_n531_));
  INV_X1    g330(.A(G8gat), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT14), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G15gat), .B(G22gat), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G1gat), .B(G8gat), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n535_), .A2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n533_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(G29gat), .B(G36gat), .Z(new_n541_));
  XOR2_X1   g340(.A(G43gat), .B(G50gat), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G229gat), .A2(G233gat), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT15), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n543_), .B(new_n546_), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n544_), .B(new_n545_), .C1(new_n547_), .C2(new_n540_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n543_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n540_), .B(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n548_), .B1(new_n550_), .B2(new_n545_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G113gat), .B(G141gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G169gat), .B(G197gat), .ZN(new_n553_));
  XOR2_X1   g352(.A(new_n552_), .B(new_n553_), .Z(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n551_), .A2(new_n555_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n548_), .B(new_n554_), .C1(new_n550_), .C2(new_n545_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT77), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NOR3_X1   g359(.A1(new_n411_), .A2(new_n530_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n480_), .A2(new_n543_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n543_), .B(KEYINPUT15), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(new_n496_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G232gat), .A2(G233gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT34), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n566_), .A2(KEYINPUT35), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n562_), .A2(new_n564_), .A3(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(KEYINPUT35), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n569_), .B(KEYINPUT74), .Z(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n568_), .A2(new_n571_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n562_), .A2(new_n564_), .A3(new_n567_), .A4(new_n570_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT75), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G190gat), .B(G218gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G134gat), .B(G162gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  OAI22_X1  g377(.A1(new_n574_), .A2(new_n575_), .B1(KEYINPUT36), .B2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(KEYINPUT36), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n572_), .A2(KEYINPUT75), .A3(new_n573_), .A4(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n574_), .A2(KEYINPUT36), .A3(new_n578_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT37), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT37), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n582_), .A2(new_n583_), .A3(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n440_), .B(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(new_n540_), .ZN(new_n591_));
  XOR2_X1   g390(.A(G127gat), .B(G155gat), .Z(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT16), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G183gat), .B(G211gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT17), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n595_), .A2(new_n596_), .ZN(new_n598_));
  OR3_X1    g397(.A1(new_n591_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n591_), .A2(new_n597_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n588_), .A2(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n561_), .A2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n301_), .A2(new_n302_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n603_), .A2(new_n604_), .A3(new_n531_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT38), .ZN(new_n606_));
  INV_X1    g405(.A(G1gat), .ZN(new_n607_));
  INV_X1    g406(.A(new_n584_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n529_), .A2(new_n558_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT101), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n408_), .A2(new_n410_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n404_), .B1(new_n409_), .B2(new_n300_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n254_), .B1(new_n613_), .B2(new_n395_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n401_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n612_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n601_), .ZN(new_n617_));
  AND4_X1   g416(.A1(new_n608_), .A2(new_n611_), .A3(new_n616_), .A4(new_n617_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n618_), .A2(new_n604_), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n606_), .B1(new_n607_), .B2(new_n619_), .ZN(G1324gat));
  NAND2_X1  g419(.A1(new_n406_), .A2(new_n407_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n603_), .A2(new_n532_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT39), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n618_), .A2(new_n622_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n624_), .B1(new_n625_), .B2(G8gat), .ZN(new_n626_));
  AOI211_X1 g425(.A(KEYINPUT39), .B(new_n532_), .C1(new_n618_), .C2(new_n622_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n623_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n628_), .B(new_n630_), .ZN(G1325gat));
  INV_X1    g430(.A(G15gat), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n632_), .B1(new_n618_), .B2(new_n255_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT41), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n603_), .A2(new_n632_), .A3(new_n255_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(G1326gat));
  INV_X1    g435(.A(G22gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n383_), .B(KEYINPUT103), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n618_), .B2(new_n638_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT42), .Z(new_n640_));
  NAND2_X1  g439(.A1(new_n638_), .A2(new_n637_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT104), .Z(new_n642_));
  NAND2_X1  g441(.A1(new_n603_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(new_n643_), .ZN(G1327gat));
  NOR2_X1   g443(.A1(new_n617_), .A2(new_n608_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n561_), .A2(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(G29gat), .B1(new_n646_), .B2(new_n604_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n611_), .A2(new_n601_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n588_), .ZN(new_n649_));
  OAI21_X1  g448(.A(KEYINPUT43), .B1(new_n411_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n616_), .A2(new_n651_), .A3(new_n588_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n648_), .A2(KEYINPUT44), .A3(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(KEYINPUT44), .B1(new_n648_), .B2(new_n653_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n604_), .A2(G29gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n647_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT105), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n658_), .B(new_n659_), .ZN(G1328gat));
  INV_X1    g459(.A(G36gat), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n646_), .A2(new_n661_), .A3(new_n622_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT45), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n654_), .A2(new_n655_), .A3(new_n621_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n663_), .B1(new_n661_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT46), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  OAI211_X1 g466(.A(new_n663_), .B(KEYINPUT46), .C1(new_n664_), .C2(new_n661_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1329gat));
  AOI21_X1  g468(.A(G43gat), .B1(new_n646_), .B2(new_n255_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n255_), .A2(G43gat), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n656_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT47), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n672_), .B(new_n673_), .ZN(G1330gat));
  AOI21_X1  g473(.A(G50gat), .B1(new_n646_), .B2(new_n638_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n383_), .A2(G50gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n656_), .B2(new_n676_), .ZN(G1331gat));
  INV_X1    g476(.A(new_n558_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n530_), .A2(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n411_), .A2(new_n679_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n680_), .A2(new_n602_), .ZN(new_n681_));
  AOI21_X1  g480(.A(G57gat), .B1(new_n681_), .B2(new_n604_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n617_), .A2(new_n560_), .ZN(new_n683_));
  NOR4_X1   g482(.A1(new_n411_), .A2(new_n584_), .A3(new_n529_), .A4(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n604_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n685_), .A2(KEYINPUT106), .ZN(new_n686_));
  MUX2_X1   g485(.A(KEYINPUT106), .B(new_n686_), .S(G57gat), .Z(new_n687_));
  AOI21_X1  g486(.A(new_n682_), .B1(new_n684_), .B2(new_n687_), .ZN(G1332gat));
  AOI21_X1  g487(.A(new_n423_), .B1(new_n684_), .B2(new_n622_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT48), .Z(new_n690_));
  NAND3_X1  g489(.A1(new_n681_), .A2(new_n423_), .A3(new_n622_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1333gat));
  AOI21_X1  g491(.A(new_n232_), .B1(new_n684_), .B2(new_n255_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT49), .Z(new_n694_));
  NAND3_X1  g493(.A1(new_n681_), .A2(new_n232_), .A3(new_n255_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1334gat));
  AOI21_X1  g495(.A(new_n373_), .B1(new_n684_), .B2(new_n638_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT50), .Z(new_n698_));
  NAND3_X1  g497(.A1(new_n681_), .A2(new_n373_), .A3(new_n638_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1335gat));
  AND2_X1   g499(.A1(new_n680_), .A2(new_n645_), .ZN(new_n701_));
  INV_X1    g500(.A(G85gat), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n701_), .A2(new_n702_), .A3(new_n604_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n650_), .A2(new_n652_), .A3(new_n705_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n679_), .A2(new_n617_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n705_), .B1(new_n650_), .B2(new_n652_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n704_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n653_), .A2(KEYINPUT107), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n711_), .A2(KEYINPUT108), .A3(new_n706_), .A4(new_n707_), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n710_), .A2(new_n604_), .A3(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n703_), .B1(new_n713_), .B2(new_n702_), .ZN(G1336gat));
  AOI21_X1  g513(.A(G92gat), .B1(new_n701_), .B2(new_n622_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT109), .ZN(new_n716_));
  NAND4_X1  g515(.A1(new_n710_), .A2(new_n712_), .A3(G92gat), .A4(new_n622_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1337gat));
  NAND3_X1  g517(.A1(new_n710_), .A2(new_n255_), .A3(new_n712_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(G99gat), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT110), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n254_), .B1(new_n446_), .B2(new_n445_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n701_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n720_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT51), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT51), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n720_), .A2(new_n726_), .A3(new_n723_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(G1338gat));
  NAND3_X1  g527(.A1(new_n701_), .A2(new_n375_), .A3(new_n383_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n653_), .A2(new_n383_), .A3(new_n707_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(G106gat), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n731_), .A2(KEYINPUT52), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n731_), .A2(KEYINPUT52), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n729_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g534(.A(KEYINPUT117), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT54), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n683_), .A2(new_n588_), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n529_), .A2(new_n737_), .A3(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n737_), .B1(new_n529_), .B2(new_n738_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT57), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT72), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n744_), .B1(new_n523_), .B2(new_n513_), .ZN(new_n745_));
  AND4_X1   g544(.A1(new_n744_), .A2(new_n505_), .A3(new_n507_), .A4(new_n513_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n558_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT55), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n505_), .A2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n519_), .A2(KEYINPUT55), .A3(new_n522_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n498_), .A2(new_n504_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n414_), .B1(new_n751_), .B2(new_n516_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n749_), .A2(new_n750_), .A3(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(new_n512_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT56), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n753_), .A2(KEYINPUT56), .A3(new_n512_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n747_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n545_), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n544_), .B(new_n759_), .C1(new_n547_), .C2(new_n540_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n760_), .B(new_n555_), .C1(new_n550_), .C2(new_n759_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT111), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n557_), .A2(new_n761_), .A3(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n557_), .A2(new_n761_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT111), .ZN(new_n765_));
  AOI22_X1  g564(.A1(new_n515_), .A2(new_n524_), .B1(new_n763_), .B2(new_n765_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n758_), .A2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n743_), .B1(new_n767_), .B2(new_n584_), .ZN(new_n768_));
  OAI211_X1 g567(.A(KEYINPUT57), .B(new_n608_), .C1(new_n758_), .C2(new_n766_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT113), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n765_), .A2(new_n763_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n771_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n772_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n770_), .B(new_n588_), .C1(new_n773_), .C2(KEYINPUT58), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(KEYINPUT58), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT58), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n753_), .A2(KEYINPUT56), .A3(new_n512_), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT56), .B1(new_n753_), .B2(new_n512_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n777_), .B1(new_n780_), .B2(new_n772_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n770_), .B1(new_n781_), .B2(new_n588_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n768_), .B(new_n769_), .C1(new_n776_), .C2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n601_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n742_), .A2(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n408_), .A2(new_n604_), .A3(new_n255_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n786_), .A2(KEYINPUT59), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(G113gat), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n560_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n793_));
  OAI21_X1  g592(.A(KEYINPUT114), .B1(new_n776_), .B2(new_n782_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n756_), .A2(new_n757_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n772_), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT58), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT113), .B1(new_n797_), .B2(new_n649_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n798_), .A2(new_n799_), .A3(new_n774_), .A4(new_n775_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT112), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n769_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n768_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n801_), .B(new_n743_), .C1(new_n767_), .C2(new_n584_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n794_), .A2(new_n800_), .A3(new_n803_), .A4(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n601_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n786_), .B1(new_n806_), .B2(new_n742_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT59), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n793_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n741_), .B1(new_n805_), .B2(new_n601_), .ZN(new_n810_));
  OAI211_X1 g609(.A(KEYINPUT116), .B(KEYINPUT59), .C1(new_n810_), .C2(new_n786_), .ZN(new_n811_));
  AOI211_X1 g610(.A(new_n789_), .B(new_n792_), .C1(new_n809_), .C2(new_n811_), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n810_), .A2(new_n678_), .A3(new_n786_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT115), .B1(new_n813_), .B2(G113gat), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n806_), .A2(new_n742_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n786_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n558_), .A3(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n790_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n814_), .A2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n736_), .B1(new_n812_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n809_), .A2(new_n811_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n822_), .A2(new_n788_), .A3(new_n791_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n814_), .A2(new_n819_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(KEYINPUT117), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n821_), .A2(new_n825_), .ZN(G1340gat));
  INV_X1    g625(.A(G120gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n529_), .B2(KEYINPUT60), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n807_), .B(new_n828_), .C1(KEYINPUT60), .C2(new_n827_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n789_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n830_), .A2(new_n530_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n829_), .B1(new_n831_), .B2(new_n827_), .ZN(G1341gat));
  AOI21_X1  g631(.A(G127gat), .B1(new_n807_), .B2(new_n617_), .ZN(new_n833_));
  INV_X1    g632(.A(G127gat), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n834_), .B1(new_n617_), .B2(KEYINPUT118), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n835_), .B1(KEYINPUT118), .B2(new_n834_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n833_), .B1(new_n830_), .B2(new_n836_), .ZN(G1342gat));
  AOI21_X1  g636(.A(G134gat), .B1(new_n807_), .B2(new_n584_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n588_), .A2(G134gat), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(KEYINPUT119), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n838_), .B1(new_n830_), .B2(new_n840_), .ZN(G1343gat));
  NOR2_X1   g640(.A1(new_n255_), .A2(new_n395_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n842_), .A2(new_n604_), .A3(new_n621_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(KEYINPUT120), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n815_), .A2(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n845_), .A2(new_n678_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(new_n259_), .ZN(G1344gat));
  NOR2_X1   g646(.A1(new_n845_), .A2(new_n529_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(new_n260_), .ZN(G1345gat));
  NOR2_X1   g648(.A1(new_n845_), .A2(new_n601_), .ZN(new_n850_));
  XOR2_X1   g649(.A(KEYINPUT61), .B(G155gat), .Z(new_n851_));
  XNOR2_X1  g650(.A(new_n850_), .B(new_n851_), .ZN(G1346gat));
  INV_X1    g651(.A(G162gat), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n845_), .A2(new_n853_), .A3(new_n649_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n845_), .B2(new_n608_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT121), .ZN(new_n856_));
  OR2_X1    g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n856_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n854_), .B1(new_n857_), .B2(new_n858_), .ZN(G1347gat));
  AOI21_X1  g658(.A(new_n638_), .B1(new_n742_), .B2(new_n784_), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n621_), .A2(new_n604_), .A3(new_n254_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n558_), .A3(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT62), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n862_), .A2(new_n863_), .A3(G169gat), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n862_), .A2(new_n305_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n863_), .B1(new_n862_), .B2(G169gat), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n865_), .B1(new_n866_), .B2(new_n867_), .ZN(G1348gat));
  NAND3_X1  g667(.A1(new_n860_), .A2(new_n530_), .A3(new_n861_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n810_), .A2(new_n383_), .ZN(new_n870_));
  AND3_X1   g669(.A1(new_n861_), .A2(new_n530_), .A3(G176gat), .ZN(new_n871_));
  AOI22_X1  g670(.A1(new_n869_), .A2(new_n218_), .B1(new_n870_), .B2(new_n871_), .ZN(G1349gat));
  NAND3_X1  g671(.A1(new_n870_), .A2(new_n617_), .A3(new_n861_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n861_), .A2(new_n617_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n874_), .A2(new_n312_), .ZN(new_n875_));
  AOI22_X1  g674(.A1(new_n873_), .A2(new_n203_), .B1(new_n860_), .B2(new_n875_), .ZN(G1350gat));
  NAND2_X1  g675(.A1(new_n584_), .A2(new_n202_), .ZN(new_n877_));
  XOR2_X1   g676(.A(new_n877_), .B(KEYINPUT123), .Z(new_n878_));
  NAND3_X1  g677(.A1(new_n860_), .A2(new_n861_), .A3(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n860_), .A2(new_n588_), .A3(new_n861_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n880_), .A2(KEYINPUT122), .A3(G190gat), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(KEYINPUT122), .B1(new_n880_), .B2(G190gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n879_), .B1(new_n882_), .B2(new_n883_), .ZN(G1351gat));
  NAND3_X1  g683(.A1(new_n622_), .A2(new_n685_), .A3(new_n842_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n810_), .A2(new_n885_), .ZN(new_n886_));
  AND3_X1   g685(.A1(new_n886_), .A2(G197gat), .A3(new_n558_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n887_), .A2(KEYINPUT124), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n887_), .A2(KEYINPUT124), .ZN(new_n889_));
  AOI21_X1  g688(.A(G197gat), .B1(new_n886_), .B2(new_n558_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n888_), .A2(new_n889_), .A3(new_n890_), .ZN(G1352gat));
  NOR3_X1   g690(.A1(new_n810_), .A2(new_n529_), .A3(new_n885_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n318_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n893_), .B1(G204gat), .B2(new_n892_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(KEYINPUT125), .ZN(G1353gat));
  INV_X1    g694(.A(KEYINPUT63), .ZN(new_n896_));
  INV_X1    g695(.A(G211gat), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n617_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(KEYINPUT126), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n886_), .A2(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n896_), .A2(new_n897_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n900_), .B(new_n901_), .ZN(G1354gat));
  AOI21_X1  g701(.A(G218gat), .B1(new_n886_), .B2(new_n584_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n588_), .A2(G218gat), .ZN(new_n904_));
  XOR2_X1   g703(.A(new_n904_), .B(KEYINPUT127), .Z(new_n905_));
  AOI21_X1  g704(.A(new_n903_), .B1(new_n886_), .B2(new_n905_), .ZN(G1355gat));
endmodule


