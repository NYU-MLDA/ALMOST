//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 1 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 0 1 1 1 0 1 0 0 1 1 1 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n651_, new_n652_, new_n653_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n826_, new_n827_, new_n828_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n843_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n861_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n868_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT23), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND3_X1  g003(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n205_));
  OAI211_X1 g004(.A(new_n204_), .B(new_n205_), .C1(G183gat), .C2(G190gat), .ZN(new_n206_));
  INV_X1    g005(.A(G169gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT22), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT22), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G169gat), .ZN(new_n210_));
  INV_X1    g009(.A(G176gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n208_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT82), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  AND3_X1   g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n213_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n206_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n207_), .A2(new_n211_), .ZN(new_n218_));
  AND3_X1   g017(.A1(new_n218_), .A2(KEYINPUT24), .A3(new_n214_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT24), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n220_), .A2(new_n207_), .A3(new_n211_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n219_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT26), .B(G190gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT81), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT25), .B(G183gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT26), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(G190gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(new_n225_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n227_), .A2(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n223_), .B1(new_n226_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n217_), .A2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(new_n233_), .B(KEYINPUT30), .Z(new_n234_));
  XOR2_X1   g033(.A(G71gat), .B(G99gat), .Z(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT31), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(new_n237_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(KEYINPUT84), .B(G15gat), .Z(new_n241_));
  NAND2_X1  g040(.A1(G227gat), .A2(G233gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT83), .B(G43gat), .ZN(new_n244_));
  XOR2_X1   g043(.A(new_n243_), .B(new_n244_), .Z(new_n245_));
  XOR2_X1   g044(.A(G127gat), .B(G134gat), .Z(new_n246_));
  XOR2_X1   g045(.A(G113gat), .B(G120gat), .Z(new_n247_));
  XOR2_X1   g046(.A(new_n246_), .B(new_n247_), .Z(new_n248_));
  XNOR2_X1  g047(.A(new_n245_), .B(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n240_), .A2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n238_), .A2(new_n239_), .A3(new_n249_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT86), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT85), .ZN(new_n255_));
  INV_X1    g054(.A(G155gat), .ZN(new_n256_));
  INV_X1    g055(.A(G162gat), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G155gat), .A2(G162gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT1), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(G155gat), .A3(G162gat), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT85), .B1(G155gat), .B2(G162gat), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n258_), .A2(new_n260_), .A3(new_n262_), .A4(new_n263_), .ZN(new_n264_));
  XOR2_X1   g063(.A(G141gat), .B(G148gat), .Z(new_n265_));
  AND2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n258_), .A2(new_n263_), .A3(new_n259_), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NOR3_X1   g068(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n267_), .B1(new_n271_), .B2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n254_), .B1(new_n266_), .B2(new_n276_), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n258_), .A2(new_n263_), .A3(new_n259_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT3), .ZN(new_n279_));
  INV_X1    g078(.A(G141gat), .ZN(new_n280_));
  INV_X1    g079(.A(G148gat), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G141gat), .A2(G148gat), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT2), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n282_), .A2(new_n285_), .A3(new_n272_), .A4(new_n268_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n278_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n264_), .A2(new_n265_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n287_), .A2(KEYINPUT86), .A3(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n277_), .A2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT28), .B(G22gat), .ZN(new_n291_));
  INV_X1    g090(.A(G50gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT87), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT29), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n290_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(new_n293_), .B(KEYINPUT87), .Z(new_n297_));
  AND3_X1   g096(.A1(new_n287_), .A2(KEYINPUT86), .A3(new_n288_), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT86), .B1(new_n287_), .B2(new_n288_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n295_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G228gat), .A2(G233gat), .ZN(new_n302_));
  OR2_X1    g101(.A1(G197gat), .A2(G204gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G197gat), .A2(G204gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT21), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT89), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT89), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n305_), .A2(new_n309_), .A3(new_n306_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n303_), .A2(KEYINPUT21), .A3(new_n304_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G211gat), .B(G218gat), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n308_), .A2(new_n310_), .A3(new_n311_), .A4(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n311_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n312_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  OAI211_X1 g116(.A(new_n302_), .B(new_n317_), .C1(new_n290_), .C2(new_n295_), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n287_), .A2(new_n288_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n319_), .A2(new_n295_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n311_), .A2(new_n312_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n321_), .B1(KEYINPUT89), .B2(new_n307_), .ZN(new_n322_));
  AOI22_X1  g121(.A1(new_n322_), .A2(new_n310_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n323_));
  OAI211_X1 g122(.A(G228gat), .B(G233gat), .C1(new_n320_), .C2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G78gat), .B(G106gat), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n318_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n325_), .B1(new_n318_), .B2(new_n324_), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n296_), .B(new_n301_), .C1(new_n327_), .C2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n318_), .A2(new_n324_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n325_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(KEYINPUT88), .B1(new_n301_), .B2(new_n296_), .ZN(new_n333_));
  AND3_X1   g132(.A1(new_n301_), .A2(new_n296_), .A3(KEYINPUT88), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n332_), .B(new_n326_), .C1(new_n333_), .C2(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n329_), .A2(new_n335_), .A3(KEYINPUT90), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n327_), .A2(new_n328_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT90), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n337_), .B(new_n338_), .C1(new_n333_), .C2(new_n334_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n336_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G1gat), .B(G29gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G57gat), .B(G85gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n277_), .A2(KEYINPUT94), .A3(new_n248_), .A4(new_n289_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n246_), .B(new_n247_), .ZN(new_n347_));
  NOR3_X1   g146(.A1(new_n298_), .A2(new_n299_), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT94), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n287_), .A2(new_n288_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n349_), .B1(new_n248_), .B2(new_n350_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n346_), .B1(new_n348_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT4), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT95), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n277_), .A2(new_n248_), .A3(new_n289_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n356_), .B1(new_n357_), .B2(KEYINPUT4), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n353_), .A2(new_n354_), .A3(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT4), .ZN(new_n361_));
  AOI21_X1  g160(.A(KEYINPUT94), .B1(new_n319_), .B2(new_n347_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n357_), .A2(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n361_), .B1(new_n363_), .B2(new_n346_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT95), .B1(new_n364_), .B2(new_n358_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n360_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n352_), .A2(new_n355_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n345_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n345_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n369_), .B1(new_n360_), .B2(new_n365_), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT99), .B1(new_n368_), .B2(new_n370_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n367_), .A2(new_n345_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n354_), .B1(new_n353_), .B2(new_n359_), .ZN(new_n373_));
  NOR3_X1   g172(.A1(new_n364_), .A2(KEYINPUT95), .A3(new_n358_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n372_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT99), .ZN(new_n376_));
  AOI22_X1  g175(.A1(new_n360_), .A2(new_n365_), .B1(new_n352_), .B2(new_n355_), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n375_), .B(new_n376_), .C1(new_n377_), .C2(new_n345_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G8gat), .B(G36gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT18), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G64gat), .B(G92gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n217_), .A2(new_n313_), .A3(new_n232_), .A4(new_n316_), .ZN(new_n383_));
  INV_X1    g182(.A(G190gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT26), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT91), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n229_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n386_), .B1(new_n229_), .B2(new_n385_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n219_), .B1(new_n389_), .B2(new_n227_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT92), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n222_), .A2(new_n391_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n221_), .A2(new_n204_), .A3(KEYINPUT92), .A4(new_n205_), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n212_), .A2(new_n214_), .ZN(new_n395_));
  AOI22_X1  g194(.A1(new_n390_), .A2(new_n394_), .B1(new_n206_), .B2(new_n395_), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n383_), .B(KEYINPUT20), .C1(new_n396_), .C2(new_n323_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT93), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G226gat), .A2(G233gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT19), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n397_), .A2(new_n398_), .A3(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n233_), .A2(new_n317_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n388_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n224_), .A2(new_n386_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(new_n404_), .A3(new_n227_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n219_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n405_), .A2(new_n406_), .A3(new_n392_), .A4(new_n393_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n395_), .A2(new_n206_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n407_), .A2(new_n313_), .A3(new_n316_), .A4(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n400_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n402_), .A2(new_n409_), .A3(KEYINPUT20), .A4(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n401_), .A2(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n398_), .B1(new_n397_), .B2(new_n400_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n382_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n397_), .A2(new_n400_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(KEYINPUT93), .ZN(new_n416_));
  INV_X1    g215(.A(new_n382_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n416_), .A2(new_n411_), .A3(new_n401_), .A4(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n414_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT27), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n407_), .A2(new_n408_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n317_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n422_), .A2(KEYINPUT20), .A3(new_n410_), .A4(new_n383_), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n402_), .A2(new_n409_), .A3(KEYINPUT20), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n423_), .B1(new_n424_), .B2(new_n410_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n420_), .B1(new_n425_), .B2(new_n382_), .ZN(new_n426_));
  AOI22_X1  g225(.A1(new_n419_), .A2(new_n420_), .B1(new_n418_), .B2(new_n426_), .ZN(new_n427_));
  AND4_X1   g226(.A1(new_n340_), .A2(new_n371_), .A3(new_n378_), .A4(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n419_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT97), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n430_), .A2(KEYINPUT33), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n375_), .A2(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n345_), .B1(new_n352_), .B2(new_n356_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n355_), .B1(new_n357_), .B2(KEYINPUT4), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n433_), .B1(new_n364_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n431_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n370_), .A2(new_n436_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n429_), .A2(new_n432_), .A3(new_n435_), .A4(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n412_), .A2(new_n413_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n417_), .A2(KEYINPUT32), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n440_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n425_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(KEYINPUT98), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT98), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n425_), .A2(new_n445_), .A3(new_n442_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n446_), .ZN(new_n447_));
  OAI211_X1 g246(.A(new_n441_), .B(new_n447_), .C1(new_n368_), .C2(new_n370_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n340_), .B1(new_n438_), .B2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n253_), .B1(new_n428_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT100), .ZN(new_n451_));
  INV_X1    g250(.A(new_n253_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n340_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n371_), .A2(new_n378_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n452_), .A2(new_n453_), .A3(new_n455_), .A4(new_n427_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT100), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n457_), .B(new_n253_), .C1(new_n428_), .C2(new_n449_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n451_), .A2(new_n456_), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(G1gat), .ZN(new_n460_));
  INV_X1    g259(.A(G8gat), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT14), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT75), .ZN(new_n463_));
  OR2_X1    g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n463_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G15gat), .B(G22gat), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n464_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT76), .ZN(new_n468_));
  XOR2_X1   g267(.A(G1gat), .B(G8gat), .Z(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G29gat), .B(G36gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT71), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G43gat), .B(G50gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n470_), .B(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT78), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G229gat), .A2(G233gat), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n470_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n474_), .B(KEYINPUT15), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n481_), .B(KEYINPUT79), .Z(new_n482_));
  AOI21_X1  g281(.A(new_n478_), .B1(new_n470_), .B2(new_n474_), .ZN(new_n483_));
  AOI22_X1  g282(.A1(new_n476_), .A2(new_n478_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G113gat), .B(G141gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT80), .ZN(new_n486_));
  XOR2_X1   g285(.A(G169gat), .B(G197gat), .Z(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n484_), .B(new_n488_), .Z(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n459_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT37), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT68), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G99gat), .A2(G106gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT6), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT6), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n496_), .A2(G99gat), .A3(G106gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT66), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT66), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n495_), .A2(new_n497_), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT7), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n502_), .A2(KEYINPUT65), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT65), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n504_), .A2(KEYINPUT7), .ZN(new_n505_));
  OAI22_X1  g304(.A1(new_n503_), .A2(new_n505_), .B1(G99gat), .B2(G106gat), .ZN(new_n506_));
  INV_X1    g305(.A(G99gat), .ZN(new_n507_));
  INV_X1    g306(.A(G106gat), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n507_), .B(new_n508_), .C1(new_n502_), .C2(KEYINPUT65), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n499_), .A2(new_n501_), .A3(new_n506_), .A4(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT67), .ZN(new_n511_));
  XOR2_X1   g310(.A(G85gat), .B(G92gat), .Z(new_n512_));
  NAND3_X1  g311(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT8), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n511_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n493_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n510_), .A2(new_n512_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT67), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n518_), .A2(KEYINPUT68), .A3(KEYINPUT8), .A4(new_n513_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n506_), .A2(new_n498_), .A3(new_n509_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT8), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n512_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n516_), .A2(new_n519_), .A3(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(KEYINPUT10), .B(G99gat), .Z(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(new_n508_), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n526_), .B(KEYINPUT64), .Z(new_n527_));
  NAND2_X1  g326(.A1(new_n512_), .A2(KEYINPUT9), .ZN(new_n528_));
  INV_X1    g327(.A(G85gat), .ZN(new_n529_));
  INV_X1    g328(.A(G92gat), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n528_), .B(new_n498_), .C1(KEYINPUT9), .C2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n527_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n524_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT35), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G232gat), .A2(G233gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT34), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n536_), .A2(new_n480_), .B1(new_n537_), .B2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n524_), .A2(new_n535_), .A3(new_n474_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT72), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n542_), .A2(new_n543_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n541_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n540_), .A2(new_n537_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  OAI221_X1 g347(.A(new_n541_), .B1(new_n537_), .B2(new_n540_), .C1(new_n544_), .C2(new_n545_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT74), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n548_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G190gat), .B(G218gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT73), .ZN(new_n553_));
  XOR2_X1   g352(.A(G134gat), .B(G162gat), .Z(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n555_), .A2(KEYINPUT36), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n551_), .A2(new_n557_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n548_), .A2(new_n549_), .A3(new_n550_), .A4(new_n556_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n555_), .A2(KEYINPUT36), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n561_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n492_), .B1(new_n560_), .B2(new_n563_), .ZN(new_n564_));
  AOI211_X1 g363(.A(KEYINPUT37), .B(new_n562_), .C1(new_n558_), .C2(new_n559_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G57gat), .B(G64gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT69), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT11), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(G71gat), .B(G78gat), .Z(new_n571_));
  OR2_X1    g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n568_), .A2(new_n569_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n570_), .A2(new_n573_), .A3(new_n571_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(new_n470_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT17), .ZN(new_n580_));
  XOR2_X1   g379(.A(G127gat), .B(G155gat), .Z(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT16), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G183gat), .B(G211gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  OR3_X1    g383(.A1(new_n579_), .A2(new_n580_), .A3(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(KEYINPUT17), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n579_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n566_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n575_), .ZN(new_n590_));
  AOI21_X1  g389(.A(KEYINPUT12), .B1(new_n536_), .B2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n536_), .A2(new_n590_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n524_), .A2(new_n575_), .A3(new_n535_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n591_), .B1(new_n594_), .B2(KEYINPUT12), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G230gat), .A2(G233gat), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n594_), .A2(G230gat), .A3(G233gat), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(G120gat), .B(G148gat), .Z(new_n600_));
  XNOR2_X1  g399(.A(G176gat), .B(G204gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n602_), .B(new_n603_), .Z(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n599_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n597_), .A2(new_n598_), .A3(new_n604_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT13), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n589_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT77), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n491_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n612_), .B1(new_n611_), .B2(new_n610_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT101), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n615_), .A2(new_n460_), .A3(new_n454_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT38), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n560_), .A2(new_n563_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n459_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n588_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n621_), .A2(new_n609_), .A3(new_n622_), .A4(new_n490_), .ZN(new_n623_));
  OAI21_X1  g422(.A(G1gat), .B1(new_n623_), .B2(new_n455_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n616_), .A2(new_n617_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n618_), .A2(new_n624_), .A3(new_n625_), .ZN(G1324gat));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT102), .ZN(new_n628_));
  OR3_X1    g427(.A1(new_n623_), .A2(new_n628_), .A3(new_n427_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n628_), .B1(new_n623_), .B2(new_n427_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(G8gat), .A3(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n631_), .A2(KEYINPUT103), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n631_), .A2(KEYINPUT103), .ZN(new_n633_));
  OAI211_X1 g432(.A(KEYINPUT104), .B(new_n627_), .C1(new_n632_), .C2(new_n633_), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n631_), .A2(KEYINPUT103), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n631_), .A2(KEYINPUT103), .ZN(new_n636_));
  XNOR2_X1  g435(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n635_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n427_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n615_), .A2(new_n461_), .A3(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n634_), .A2(new_n638_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT40), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n634_), .A2(new_n638_), .A3(new_n640_), .A4(KEYINPUT40), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(G1325gat));
  OAI21_X1  g444(.A(G15gat), .B1(new_n623_), .B2(new_n253_), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n646_), .B(KEYINPUT41), .Z(new_n647_));
  INV_X1    g446(.A(new_n615_), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n253_), .A2(G15gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n647_), .B1(new_n648_), .B2(new_n649_), .ZN(G1326gat));
  OAI21_X1  g449(.A(G22gat), .B1(new_n623_), .B2(new_n453_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT42), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n453_), .A2(G22gat), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n652_), .B1(new_n648_), .B2(new_n653_), .ZN(G1327gat));
  INV_X1    g453(.A(new_n609_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n655_), .A2(new_n622_), .A3(new_n620_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(new_n491_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(G29gat), .B1(new_n658_), .B2(new_n454_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n655_), .A2(new_n622_), .A3(new_n489_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT106), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT43), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n458_), .A2(new_n456_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n438_), .A2(new_n448_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(new_n453_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n340_), .A2(new_n371_), .A3(new_n427_), .A4(new_n378_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n457_), .B1(new_n667_), .B2(new_n253_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n662_), .B1(new_n663_), .B2(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n564_), .A2(new_n565_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n661_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n566_), .A2(new_n459_), .A3(KEYINPUT106), .A4(new_n662_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n670_), .B1(new_n459_), .B2(new_n674_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n451_), .A2(KEYINPUT105), .A3(new_n456_), .A4(new_n458_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n662_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n660_), .B1(new_n673_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  OAI211_X1 g479(.A(KEYINPUT44), .B(new_n660_), .C1(new_n673_), .C2(new_n677_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n454_), .A2(G29gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n659_), .B1(new_n682_), .B2(new_n683_), .ZN(G1328gat));
  INV_X1    g483(.A(KEYINPUT109), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n680_), .A2(new_n639_), .A3(new_n681_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT107), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n686_), .A2(new_n687_), .A3(G36gat), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n427_), .A2(G36gat), .ZN(new_n689_));
  OR3_X1    g488(.A1(new_n657_), .A2(KEYINPUT108), .A3(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(KEYINPUT108), .B1(new_n657_), .B2(new_n689_), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n690_), .A2(KEYINPUT45), .A3(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(KEYINPUT45), .B1(new_n690_), .B2(new_n691_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n688_), .A2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n687_), .B1(new_n686_), .B2(G36gat), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n685_), .B(KEYINPUT46), .C1(new_n695_), .C2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n686_), .A2(G36gat), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(KEYINPUT107), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n700_), .A2(new_n688_), .A3(new_n694_), .ZN(new_n701_));
  AOI21_X1  g500(.A(KEYINPUT46), .B1(new_n701_), .B2(new_n685_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n698_), .A2(new_n702_), .ZN(G1329gat));
  AOI21_X1  g502(.A(G43gat), .B1(new_n658_), .B2(new_n452_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n452_), .A2(G43gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n682_), .B2(new_n705_), .ZN(new_n706_));
  XOR2_X1   g505(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n707_));
  XNOR2_X1  g506(.A(new_n706_), .B(new_n707_), .ZN(G1330gat));
  NAND3_X1  g507(.A1(new_n658_), .A2(new_n292_), .A3(new_n340_), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT111), .B1(new_n682_), .B2(new_n340_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n680_), .A2(KEYINPUT111), .A3(new_n340_), .A4(new_n681_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(G50gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n709_), .B1(new_n710_), .B2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT112), .ZN(G1331gat));
  NOR2_X1   g513(.A1(new_n609_), .A2(new_n490_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n715_), .A2(new_n459_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n716_), .A2(new_n589_), .ZN(new_n717_));
  INV_X1    g516(.A(G57gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n717_), .A2(new_n718_), .A3(new_n454_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n621_), .A2(new_n622_), .A3(new_n715_), .ZN(new_n720_));
  OAI21_X1  g519(.A(G57gat), .B1(new_n720_), .B2(new_n455_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(G1332gat));
  OAI21_X1  g521(.A(G64gat), .B1(new_n720_), .B2(new_n427_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT48), .ZN(new_n724_));
  INV_X1    g523(.A(G64gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n717_), .A2(new_n725_), .A3(new_n639_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1333gat));
  OAI21_X1  g526(.A(G71gat), .B1(new_n720_), .B2(new_n253_), .ZN(new_n728_));
  XOR2_X1   g527(.A(KEYINPUT113), .B(KEYINPUT49), .Z(new_n729_));
  XNOR2_X1  g528(.A(new_n728_), .B(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(G71gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n717_), .A2(new_n731_), .A3(new_n452_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(G1334gat));
  OAI21_X1  g532(.A(G78gat), .B1(new_n720_), .B2(new_n453_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT50), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n453_), .A2(G78gat), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT114), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n717_), .A2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n735_), .A2(new_n738_), .ZN(G1335gat));
  NAND3_X1  g538(.A1(new_n716_), .A2(new_n588_), .A3(new_n619_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT115), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n741_), .A2(new_n529_), .A3(new_n454_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n673_), .A2(new_n677_), .ZN(new_n743_));
  NOR4_X1   g542(.A1(new_n743_), .A2(new_n609_), .A3(new_n622_), .A4(new_n490_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n454_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n742_), .B1(new_n746_), .B2(new_n529_), .ZN(G1336gat));
  NAND3_X1  g546(.A1(new_n741_), .A2(new_n530_), .A3(new_n639_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n744_), .A2(new_n639_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n748_), .B1(new_n750_), .B2(new_n530_), .ZN(G1337gat));
  AOI21_X1  g550(.A(new_n507_), .B1(new_n744_), .B2(new_n452_), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n741_), .A2(new_n525_), .A3(new_n452_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g554(.A1(new_n741_), .A2(new_n508_), .A3(new_n340_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n744_), .A2(new_n340_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n758_), .B2(G106gat), .ZN(new_n759_));
  AOI211_X1 g558(.A(KEYINPUT52), .B(new_n508_), .C1(new_n744_), .C2(new_n340_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n756_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT53), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT53), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n763_), .B(new_n756_), .C1(new_n759_), .C2(new_n760_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(G1339gat));
  NOR3_X1   g564(.A1(new_n455_), .A2(new_n253_), .A3(new_n639_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n477_), .B1(new_n470_), .B2(new_n474_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n488_), .B1(new_n482_), .B2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n476_), .A2(new_n477_), .ZN(new_n769_));
  AOI22_X1  g568(.A1(new_n484_), .A2(new_n488_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n608_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT55), .ZN(new_n772_));
  OAI21_X1  g571(.A(KEYINPUT116), .B1(new_n597_), .B2(new_n772_), .ZN(new_n773_));
  OR2_X1    g572(.A1(new_n595_), .A2(new_n596_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n597_), .A2(new_n772_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n595_), .A2(new_n776_), .A3(KEYINPUT55), .A4(new_n596_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n773_), .A2(new_n774_), .A3(new_n775_), .A4(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n605_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT117), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT56), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n778_), .A2(KEYINPUT117), .A3(new_n605_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n607_), .B(new_n490_), .C1(new_n783_), .C2(KEYINPUT118), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n778_), .A2(KEYINPUT56), .A3(new_n605_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT118), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n786_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n771_), .B1(new_n784_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n620_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT57), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n619_), .A2(new_n790_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n770_), .A2(new_n607_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT119), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n770_), .A2(KEYINPUT119), .A3(new_n607_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT56), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n779_), .A2(new_n797_), .ZN(new_n798_));
  AOI22_X1  g597(.A1(new_n795_), .A2(new_n796_), .B1(new_n798_), .B2(new_n785_), .ZN(new_n799_));
  OR2_X1    g598(.A1(new_n799_), .A2(KEYINPUT58), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n670_), .B1(new_n799_), .B2(KEYINPUT58), .ZN(new_n801_));
  AOI22_X1  g600(.A1(new_n788_), .A2(new_n792_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n622_), .B1(new_n791_), .B2(new_n802_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n610_), .A2(new_n490_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT54), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n453_), .B(new_n766_), .C1(new_n803_), .C2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT59), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n788_), .A2(new_n792_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n800_), .A2(new_n801_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT57), .B1(new_n788_), .B2(new_n620_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n588_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n805_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n815_), .A2(KEYINPUT59), .A3(new_n453_), .A4(new_n766_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n489_), .B1(new_n808_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(G113gat), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n490_), .A2(new_n818_), .ZN(new_n819_));
  OAI22_X1  g618(.A1(new_n817_), .A2(new_n818_), .B1(new_n806_), .B2(new_n819_), .ZN(G1340gat));
  AOI21_X1  g619(.A(new_n609_), .B1(new_n808_), .B2(new_n816_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(KEYINPUT120), .B(G120gat), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n822_), .B1(new_n609_), .B2(KEYINPUT60), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(KEYINPUT60), .B2(new_n822_), .ZN(new_n824_));
  OAI22_X1  g623(.A1(new_n821_), .A2(new_n822_), .B1(new_n806_), .B2(new_n824_), .ZN(G1341gat));
  AOI21_X1  g624(.A(new_n588_), .B1(new_n808_), .B2(new_n816_), .ZN(new_n826_));
  INV_X1    g625(.A(G127gat), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n622_), .A2(new_n827_), .ZN(new_n828_));
  OAI22_X1  g627(.A1(new_n826_), .A2(new_n827_), .B1(new_n806_), .B2(new_n828_), .ZN(G1342gat));
  INV_X1    g628(.A(G134gat), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(new_n806_), .B2(new_n620_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT121), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT121), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n833_), .B(new_n830_), .C1(new_n806_), .C2(new_n620_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n808_), .A2(new_n816_), .ZN(new_n835_));
  XOR2_X1   g634(.A(KEYINPUT122), .B(G134gat), .Z(new_n836_));
  NOR2_X1   g635(.A1(new_n670_), .A2(new_n836_), .ZN(new_n837_));
  AOI22_X1  g636(.A1(new_n832_), .A2(new_n834_), .B1(new_n835_), .B2(new_n837_), .ZN(G1343gat));
  NOR4_X1   g637(.A1(new_n452_), .A2(new_n455_), .A3(new_n453_), .A4(new_n639_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n815_), .A2(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n840_), .A2(new_n489_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(new_n280_), .ZN(G1344gat));
  NOR2_X1   g641(.A1(new_n840_), .A2(new_n609_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(new_n281_), .ZN(G1345gat));
  NOR2_X1   g643(.A1(new_n840_), .A2(new_n588_), .ZN(new_n845_));
  XOR2_X1   g644(.A(KEYINPUT61), .B(G155gat), .Z(new_n846_));
  XNOR2_X1  g645(.A(new_n845_), .B(new_n846_), .ZN(G1346gat));
  OAI21_X1  g646(.A(G162gat), .B1(new_n840_), .B2(new_n670_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n619_), .A2(new_n257_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n840_), .B2(new_n849_), .ZN(G1347gat));
  NOR3_X1   g649(.A1(new_n253_), .A2(new_n454_), .A3(new_n427_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n490_), .A2(new_n851_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(KEYINPUT123), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n815_), .A2(new_n453_), .A3(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT62), .ZN(new_n855_));
  AND3_X1   g654(.A1(new_n854_), .A2(new_n855_), .A3(G169gat), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n855_), .B1(new_n854_), .B2(G169gat), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n815_), .A2(new_n453_), .A3(new_n851_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n490_), .A2(new_n208_), .A3(new_n210_), .ZN(new_n859_));
  OAI22_X1  g658(.A1(new_n856_), .A2(new_n857_), .B1(new_n858_), .B2(new_n859_), .ZN(G1348gat));
  NOR2_X1   g659(.A1(new_n858_), .A2(new_n609_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(new_n211_), .ZN(G1349gat));
  NOR2_X1   g661(.A1(new_n858_), .A2(new_n588_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(G183gat), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n858_), .A2(new_n588_), .A3(new_n227_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n864_), .A2(new_n865_), .ZN(G1350gat));
  OAI21_X1  g665(.A(G190gat), .B1(new_n858_), .B2(new_n670_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n619_), .A2(new_n389_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n858_), .B2(new_n868_), .ZN(G1351gat));
  NOR2_X1   g668(.A1(new_n452_), .A2(new_n453_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n870_), .A2(new_n455_), .A3(new_n639_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n871_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n490_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g673(.A1(new_n872_), .A2(new_n655_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT124), .B(G204gat), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n875_), .B(new_n876_), .ZN(G1353gat));
  INV_X1    g676(.A(KEYINPUT126), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n588_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n879_));
  XOR2_X1   g678(.A(new_n879_), .B(KEYINPUT125), .Z(new_n880_));
  NAND3_X1  g679(.A1(new_n872_), .A2(new_n878_), .A3(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n871_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n882_), .B(new_n880_), .C1(new_n803_), .C2(new_n805_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(KEYINPUT126), .ZN(new_n884_));
  NOR2_X1   g683(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n881_), .A2(new_n884_), .A3(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n885_), .B1(new_n881_), .B2(new_n884_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1354gat));
  INV_X1    g687(.A(KEYINPUT127), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n620_), .A2(G218gat), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n872_), .A2(new_n890_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n872_), .A2(new_n566_), .ZN(new_n892_));
  INV_X1    g691(.A(G218gat), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n889_), .B(new_n891_), .C1(new_n892_), .C2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n891_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n872_), .B2(new_n566_), .ZN(new_n896_));
  OAI21_X1  g695(.A(KEYINPUT127), .B1(new_n895_), .B2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n894_), .A2(new_n897_), .ZN(G1355gat));
endmodule


