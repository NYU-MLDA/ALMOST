//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 1 1 0 1 1 0 0 0 1 0 1 1 0 1 0 1 0 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1 0 1 1 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n868_, new_n869_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(new_n202_), .A2(KEYINPUT23), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT85), .B(KEYINPUT23), .ZN(new_n204_));
  INV_X1    g003(.A(new_n202_), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n203_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G169gat), .ZN(new_n207_));
  INV_X1    g006(.A(G176gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n209_), .A2(KEYINPUT24), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n209_), .A2(KEYINPUT24), .A3(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT25), .B(G183gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT83), .ZN(new_n214_));
  INV_X1    g013(.A(G190gat), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n215_), .A2(KEYINPUT26), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n213_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT26), .B(G190gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n218_), .A2(KEYINPUT83), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n212_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n206_), .B(new_n210_), .C1(new_n220_), .C2(KEYINPUT84), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n220_), .A2(KEYINPUT84), .ZN(new_n222_));
  MUX2_X1   g021(.A(KEYINPUT23), .B(new_n204_), .S(new_n205_), .Z(new_n223_));
  NOR2_X1   g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(new_n207_), .ZN(new_n228_));
  OAI22_X1  g027(.A1(new_n221_), .A2(new_n222_), .B1(new_n226_), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G227gat), .A2(G233gat), .ZN(new_n230_));
  INV_X1    g029(.A(G71gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(G99gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n229_), .B(new_n233_), .ZN(new_n234_));
  XOR2_X1   g033(.A(G127gat), .B(G134gat), .Z(new_n235_));
  XOR2_X1   g034(.A(G113gat), .B(G120gat), .Z(new_n236_));
  XOR2_X1   g035(.A(new_n235_), .B(new_n236_), .Z(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n234_), .B(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G15gat), .B(G43gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT86), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT30), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT31), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n239_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT94), .B(G204gat), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT93), .B(G197gat), .ZN(new_n247_));
  OAI22_X1  g046(.A1(new_n246_), .A2(G197gat), .B1(new_n247_), .B2(G204gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT21), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(G204gat), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT21), .ZN(new_n251_));
  INV_X1    g050(.A(G197gat), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n250_), .B(new_n251_), .C1(new_n252_), .C2(new_n245_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G211gat), .B(G218gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n249_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n250_), .B1(new_n252_), .B2(new_n245_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n254_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(KEYINPUT21), .A3(new_n257_), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n255_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT2), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n260_), .A2(KEYINPUT88), .B1(G141gat), .B2(G148gat), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n261_), .B1(KEYINPUT88), .B2(new_n260_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT89), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  AND3_X1   g063(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT90), .ZN(new_n266_));
  NOR2_X1   g065(.A1(G141gat), .A2(G148gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT3), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n261_), .B(KEYINPUT89), .C1(KEYINPUT88), .C2(new_n260_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n264_), .A2(new_n266_), .A3(new_n268_), .A4(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(G155gat), .A2(G162gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT87), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G155gat), .A2(G162gat), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n270_), .A2(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(new_n273_), .B(KEYINPUT1), .Z(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(new_n272_), .ZN(new_n277_));
  XOR2_X1   g076(.A(G141gat), .B(G148gat), .Z(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n275_), .A2(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n259_), .B1(KEYINPUT29), .B2(new_n280_), .ZN(new_n281_));
  AND2_X1   g080(.A1(G228gat), .A2(G233gat), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n281_), .A2(new_n283_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G78gat), .B(G106gat), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n284_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n287_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n280_), .A2(KEYINPUT29), .ZN(new_n291_));
  XOR2_X1   g090(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  XOR2_X1   g094(.A(G22gat), .B(G50gat), .Z(new_n296_));
  NAND2_X1  g095(.A1(new_n291_), .A2(new_n293_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n295_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n296_), .B1(new_n295_), .B2(new_n297_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n290_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT92), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n303_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n284_), .A2(KEYINPUT95), .A3(new_n285_), .A4(new_n287_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n296_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n297_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n306_), .B1(new_n307_), .B2(new_n294_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n308_), .A2(new_n298_), .A3(KEYINPUT92), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n304_), .A2(new_n305_), .A3(new_n309_), .ZN(new_n310_));
  NOR3_X1   g109(.A1(new_n288_), .A2(new_n289_), .A3(KEYINPUT95), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n302_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n255_), .A2(new_n258_), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n229_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT20), .ZN(new_n316_));
  AND3_X1   g115(.A1(new_n223_), .A2(new_n212_), .A3(new_n210_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n213_), .B(KEYINPUT96), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(new_n218_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT22), .B(G169gat), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT98), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(new_n208_), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n211_), .B(KEYINPUT97), .Z(new_n324_));
  AOI21_X1  g123(.A(new_n324_), .B1(new_n206_), .B2(new_n225_), .ZN(new_n325_));
  AOI22_X1  g124(.A1(new_n317_), .A2(new_n319_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n316_), .B1(new_n327_), .B2(new_n314_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n315_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G226gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT19), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n316_), .B1(new_n259_), .B2(new_n326_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n229_), .A2(new_n314_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n331_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n333_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G8gat), .B(G36gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT18), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G64gat), .B(G92gat), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n338_), .B(new_n339_), .Z(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(KEYINPUT32), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n332_), .A2(new_n336_), .A3(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n333_), .A2(new_n334_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(new_n331_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n344_), .B1(new_n331_), .B2(new_n329_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n341_), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n342_), .A2(KEYINPUT102), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n280_), .A2(new_n237_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT99), .ZN(new_n349_));
  AOI22_X1  g148(.A1(new_n270_), .A2(new_n274_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n349_), .B1(new_n350_), .B2(new_n238_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n348_), .A2(new_n351_), .ZN(new_n352_));
  NOR3_X1   g151(.A1(new_n280_), .A2(new_n349_), .A3(new_n237_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT4), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT100), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n280_), .A2(new_n237_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n357_), .A2(KEYINPUT4), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n354_), .A2(new_n356_), .A3(new_n359_), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n352_), .A2(new_n353_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n355_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G1gat), .B(G29gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(G85gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT0), .B(G57gat), .ZN(new_n365_));
  XOR2_X1   g164(.A(new_n364_), .B(new_n365_), .Z(new_n366_));
  NAND3_X1  g165(.A1(new_n360_), .A2(new_n362_), .A3(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n366_), .B1(new_n360_), .B2(new_n362_), .ZN(new_n369_));
  OAI221_X1 g168(.A(new_n347_), .B1(KEYINPUT102), .B2(new_n342_), .C1(new_n368_), .C2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n340_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n335_), .B1(new_n315_), .B2(new_n328_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n336_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n371_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n332_), .A2(new_n340_), .A3(new_n336_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n354_), .A2(new_n355_), .A3(new_n359_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n356_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n366_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n374_), .B(new_n375_), .C1(new_n376_), .C2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n367_), .A2(KEYINPUT33), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT33), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n360_), .A2(new_n362_), .A3(new_n382_), .A4(new_n366_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n380_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n370_), .B1(new_n384_), .B2(KEYINPUT101), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT101), .ZN(new_n386_));
  AOI211_X1 g185(.A(new_n386_), .B(new_n380_), .C1(new_n381_), .C2(new_n383_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n313_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n368_), .A2(new_n369_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n312_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n374_), .A2(new_n375_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n391_), .A2(KEYINPUT27), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT103), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n375_), .A2(new_n393_), .B1(new_n345_), .B2(new_n371_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n394_), .B1(new_n393_), .B2(new_n375_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n392_), .B1(new_n395_), .B2(KEYINPUT27), .ZN(new_n396_));
  OR2_X1    g195(.A1(new_n390_), .A2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n244_), .B1(new_n388_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n396_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n313_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n389_), .A2(new_n244_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n398_), .A2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G113gat), .B(G141gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G169gat), .B(G197gat), .ZN(new_n405_));
  XOR2_X1   g204(.A(new_n404_), .B(new_n405_), .Z(new_n406_));
  NAND2_X1  g205(.A1(G229gat), .A2(G233gat), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT77), .B(G15gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(G22gat), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT14), .ZN(new_n411_));
  XOR2_X1   g210(.A(KEYINPUT78), .B(G1gat), .Z(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT79), .B(G8gat), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n411_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G1gat), .B(G8gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  OR3_X1    g215(.A1(new_n410_), .A2(new_n414_), .A3(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n416_), .B1(new_n410_), .B2(new_n414_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  XOR2_X1   g218(.A(G29gat), .B(G36gat), .Z(new_n420_));
  XOR2_X1   g219(.A(G43gat), .B(G50gat), .Z(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n419_), .A2(new_n422_), .ZN(new_n423_));
  XOR2_X1   g222(.A(new_n420_), .B(new_n421_), .Z(new_n424_));
  AOI21_X1  g223(.A(new_n424_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n408_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n422_), .B(KEYINPUT15), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n425_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(new_n429_), .A3(new_n407_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n406_), .B1(new_n426_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n426_), .A2(new_n430_), .A3(new_n406_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(KEYINPUT82), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n433_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT82), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n431_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n434_), .A2(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n403_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT37), .ZN(new_n440_));
  XOR2_X1   g239(.A(G85gat), .B(G92gat), .Z(new_n441_));
  XOR2_X1   g240(.A(KEYINPUT10), .B(G99gat), .Z(new_n442_));
  INV_X1    g241(.A(G106gat), .ZN(new_n443_));
  AOI22_X1  g242(.A1(KEYINPUT9), .A2(new_n441_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT64), .B(G92gat), .ZN(new_n445_));
  INV_X1    g244(.A(G85gat), .ZN(new_n446_));
  OR2_X1    g245(.A1(new_n446_), .A2(KEYINPUT9), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n444_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G99gat), .A2(G106gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT6), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT6), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n451_), .A2(G99gat), .A3(G106gat), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n450_), .A2(new_n452_), .A3(KEYINPUT65), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(KEYINPUT65), .B1(new_n450_), .B2(new_n452_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  OR2_X1    g256(.A1(new_n448_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT7), .ZN(new_n459_));
  INV_X1    g258(.A(G99gat), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(new_n460_), .A3(new_n443_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT67), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(G99gat), .A2(G106gat), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n464_), .A2(KEYINPUT67), .A3(new_n459_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n450_), .A2(new_n452_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT65), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT66), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT66), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n472_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n466_), .A2(new_n469_), .A3(new_n453_), .A4(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT8), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n475_), .A2(new_n476_), .A3(new_n441_), .ZN(new_n477_));
  AOI21_X1  g276(.A(KEYINPUT67), .B1(new_n464_), .B2(new_n459_), .ZN(new_n478_));
  NOR4_X1   g277(.A1(new_n462_), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n474_), .B(new_n467_), .C1(new_n478_), .C2(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n476_), .B1(new_n480_), .B2(new_n441_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n477_), .B1(new_n481_), .B2(KEYINPUT68), .ZN(new_n482_));
  INV_X1    g281(.A(new_n441_), .ZN(new_n483_));
  AOI22_X1  g282(.A1(new_n463_), .A2(new_n465_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n483_), .B1(new_n484_), .B2(new_n467_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT68), .ZN(new_n486_));
  NOR3_X1   g285(.A1(new_n485_), .A2(new_n486_), .A3(new_n476_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n458_), .B1(new_n482_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G232gat), .A2(G233gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT34), .ZN(new_n490_));
  OAI22_X1  g289(.A1(new_n488_), .A2(new_n424_), .B1(KEYINPUT35), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n490_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT35), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n488_), .A2(new_n427_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n492_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n497_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n495_), .B1(new_n499_), .B2(new_n491_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT36), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G190gat), .B(G218gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT75), .ZN(new_n503_));
  XOR2_X1   g302(.A(G134gat), .B(G162gat), .Z(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n498_), .A2(new_n500_), .A3(new_n501_), .A4(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n498_), .A2(new_n500_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n505_), .B(KEYINPUT36), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n506_), .B1(new_n509_), .B2(KEYINPUT76), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT76), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n511_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n440_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n509_), .A2(KEYINPUT37), .A3(new_n506_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G231gat), .A2(G233gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n419_), .B(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT70), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT11), .ZN(new_n519_));
  INV_X1    g318(.A(G64gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(G57gat), .ZN(new_n521_));
  INV_X1    g320(.A(G57gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(G64gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT69), .B(G71gat), .ZN(new_n525_));
  INV_X1    g324(.A(G78gat), .ZN(new_n526_));
  AOI22_X1  g325(.A1(new_n519_), .A2(new_n524_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT69), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n528_), .A2(G71gat), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n231_), .A2(KEYINPUT69), .ZN(new_n530_));
  OAI21_X1  g329(.A(G78gat), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n518_), .B1(new_n527_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n524_), .A2(new_n519_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n525_), .A2(new_n526_), .ZN(new_n534_));
  AND4_X1   g333(.A1(new_n518_), .A2(new_n533_), .A3(new_n534_), .A4(new_n531_), .ZN(new_n535_));
  OAI22_X1  g334(.A1(new_n532_), .A2(new_n535_), .B1(new_n519_), .B2(new_n524_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n533_), .A2(new_n534_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n531_), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT70), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n524_), .A2(new_n519_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n527_), .A2(new_n518_), .A3(new_n531_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n539_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n536_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n517_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n517_), .A2(new_n544_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT72), .ZN(new_n548_));
  XOR2_X1   g347(.A(G127gat), .B(G155gat), .Z(new_n549_));
  XNOR2_X1  g348(.A(G183gat), .B(G211gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n553_), .A2(KEYINPUT17), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT72), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n545_), .A2(new_n555_), .A3(new_n546_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n548_), .A2(new_n554_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT81), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT81), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n548_), .A2(new_n559_), .A3(new_n554_), .A4(new_n556_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n553_), .A2(KEYINPUT17), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n554_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n547_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n561_), .A2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n515_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT13), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G120gat), .B(G148gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT5), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G176gat), .B(G204gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT73), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G230gat), .A2(G233gat), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n481_), .A2(KEYINPUT68), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n486_), .B1(new_n485_), .B2(new_n476_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n574_), .A2(new_n575_), .A3(new_n477_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n543_), .B1(new_n576_), .B2(new_n458_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT71), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n573_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n488_), .A2(new_n544_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n576_), .A2(new_n543_), .A3(new_n458_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n580_), .A2(KEYINPUT71), .A3(new_n581_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n579_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n573_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT12), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n585_), .B(new_n458_), .C1(new_n482_), .C2(new_n487_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n448_), .A2(new_n457_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n441_), .A2(new_n476_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n588_), .B1(new_n456_), .B2(new_n484_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n480_), .A2(new_n441_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(KEYINPUT8), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n589_), .B1(new_n591_), .B2(new_n486_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n587_), .B1(new_n592_), .B2(new_n574_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(KEYINPUT72), .A2(KEYINPUT12), .ZN(new_n594_));
  OAI211_X1 g393(.A(new_n544_), .B(new_n586_), .C1(new_n593_), .C2(new_n594_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n488_), .A2(KEYINPUT72), .A3(KEYINPUT12), .A4(new_n543_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n584_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n572_), .B1(new_n583_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT74), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n586_), .A2(new_n544_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n594_), .B1(new_n576_), .B2(new_n458_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n596_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n573_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n579_), .A2(new_n582_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n604_), .A2(new_n605_), .A3(new_n571_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n598_), .A2(new_n599_), .A3(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n599_), .B1(new_n598_), .B2(new_n606_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n567_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n571_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n583_), .A2(new_n597_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n572_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n612_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n613_));
  OAI21_X1  g412(.A(KEYINPUT74), .B1(new_n611_), .B2(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n598_), .A2(new_n606_), .A3(new_n599_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n614_), .A2(KEYINPUT13), .A3(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n609_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n566_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n439_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n389_), .A2(new_n412_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(KEYINPUT38), .A3(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT104), .ZN(new_n625_));
  AOI21_X1  g424(.A(KEYINPUT38), .B1(new_n622_), .B2(new_n623_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n510_), .A2(new_n512_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n403_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n438_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n618_), .A2(KEYINPUT105), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT105), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n631_), .B1(new_n617_), .B2(new_n438_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n633_), .A2(new_n565_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n628_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n389_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n626_), .B1(G1gat), .B2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n625_), .A2(new_n639_), .ZN(G1324gat));
  OR3_X1    g439(.A1(new_n621_), .A2(new_n399_), .A3(new_n413_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n628_), .A2(new_n396_), .A3(new_n634_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT39), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n642_), .A2(new_n643_), .A3(G8gat), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n643_), .B1(new_n642_), .B2(G8gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n641_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n646_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g446(.A(new_n244_), .ZN(new_n648_));
  OR3_X1    g447(.A1(new_n621_), .A2(G15gat), .A3(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(G15gat), .B1(new_n635_), .B2(new_n648_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT41), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n650_), .A2(new_n651_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n649_), .B1(new_n652_), .B2(new_n653_), .ZN(G1326gat));
  OR3_X1    g453(.A1(new_n621_), .A2(G22gat), .A3(new_n313_), .ZN(new_n655_));
  OAI21_X1  g454(.A(G22gat), .B1(new_n635_), .B2(new_n313_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n656_), .A2(KEYINPUT42), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n656_), .A2(KEYINPUT42), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n655_), .B1(new_n657_), .B2(new_n658_), .ZN(G1327gat));
  INV_X1    g458(.A(new_n565_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n633_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n515_), .ZN(new_n663_));
  OAI21_X1  g462(.A(KEYINPUT43), .B1(new_n403_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT43), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n665_), .B(new_n515_), .C1(new_n398_), .C2(new_n402_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n662_), .B1(new_n664_), .B2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  OR2_X1    g468(.A1(new_n400_), .A2(new_n401_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n390_), .A2(new_n396_), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n384_), .A2(KEYINPUT101), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n384_), .A2(KEYINPUT101), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n672_), .A2(new_n673_), .A3(new_n370_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n671_), .B1(new_n674_), .B2(new_n313_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n670_), .B1(new_n675_), .B2(new_n244_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n665_), .B1(new_n676_), .B2(new_n515_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n666_), .ZN(new_n678_));
  OAI211_X1 g477(.A(KEYINPUT44), .B(new_n661_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n679_));
  AND4_X1   g478(.A1(G29gat), .A2(new_n669_), .A3(new_n637_), .A4(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n627_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n660_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n683_), .A2(new_n617_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n439_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(G29gat), .B1(new_n686_), .B2(new_n637_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n680_), .A2(new_n687_), .ZN(G1328gat));
  OAI211_X1 g487(.A(new_n679_), .B(new_n396_), .C1(new_n667_), .C2(new_n668_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(G36gat), .ZN(new_n690_));
  XNOR2_X1  g489(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n399_), .A2(G36gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n686_), .B2(new_n693_), .ZN(new_n694_));
  NOR4_X1   g493(.A1(new_n685_), .A2(G36gat), .A3(new_n399_), .A4(new_n691_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n690_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT46), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n690_), .A2(new_n696_), .A3(KEYINPUT46), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1329gat));
  INV_X1    g500(.A(G43gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n702_), .B1(new_n685_), .B2(new_n648_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT108), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n705_), .B(new_n702_), .C1(new_n685_), .C2(new_n648_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n648_), .A2(new_n702_), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n679_), .B(new_n708_), .C1(new_n667_), .C2(new_n668_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT47), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT47), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n707_), .A2(new_n712_), .A3(new_n709_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1330gat));
  AND4_X1   g513(.A1(G50gat), .A2(new_n669_), .A3(new_n312_), .A4(new_n679_), .ZN(new_n715_));
  AOI21_X1  g514(.A(G50gat), .B1(new_n686_), .B2(new_n312_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(G1331gat));
  INV_X1    g516(.A(KEYINPUT109), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n718_), .B1(new_n403_), .B2(new_n629_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n676_), .A2(KEYINPUT109), .A3(new_n438_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n721_), .A2(new_n566_), .A3(new_n617_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n722_), .A2(new_n522_), .A3(new_n637_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n628_), .A2(new_n438_), .A3(new_n660_), .A4(new_n617_), .ZN(new_n724_));
  OAI21_X1  g523(.A(G57gat), .B1(new_n724_), .B2(new_n389_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1332gat));
  OAI21_X1  g525(.A(G64gat), .B1(new_n724_), .B2(new_n399_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT48), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n722_), .A2(new_n520_), .A3(new_n396_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1333gat));
  OAI21_X1  g529(.A(G71gat), .B1(new_n724_), .B2(new_n648_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT49), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n722_), .A2(new_n231_), .A3(new_n244_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1334gat));
  OAI21_X1  g533(.A(G78gat), .B1(new_n724_), .B2(new_n313_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT110), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT50), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n735_), .A2(KEYINPUT110), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n735_), .A2(KEYINPUT110), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(KEYINPUT50), .A3(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n722_), .A2(new_n526_), .A3(new_n312_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n738_), .A2(new_n741_), .A3(new_n742_), .ZN(G1335gat));
  NOR2_X1   g542(.A1(new_n683_), .A2(new_n618_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n721_), .A2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n745_), .A2(new_n446_), .A3(new_n637_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n617_), .A2(new_n438_), .A3(new_n565_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT111), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n748_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  OAI211_X1 g550(.A(KEYINPUT112), .B(new_n748_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n389_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n746_), .B1(new_n753_), .B2(new_n446_), .ZN(G1336gat));
  AOI21_X1  g553(.A(G92gat), .B1(new_n745_), .B2(new_n396_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n751_), .A2(new_n752_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n399_), .A2(new_n445_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n755_), .B1(new_n756_), .B2(new_n757_), .ZN(G1337gat));
  NAND3_X1  g557(.A1(new_n745_), .A2(new_n244_), .A3(new_n442_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n648_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n759_), .B1(new_n760_), .B2(new_n460_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT51), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n763_), .B(new_n759_), .C1(new_n760_), .C2(new_n460_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(G1338gat));
  NOR2_X1   g564(.A1(new_n313_), .A2(G106gat), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n721_), .A2(new_n744_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT113), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n721_), .A2(new_n769_), .A3(new_n744_), .A4(new_n766_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n443_), .B1(KEYINPUT114), .B2(KEYINPUT52), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n772_), .B1(new_n749_), .B2(new_n313_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(KEYINPUT114), .A2(KEYINPUT52), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  OAI221_X1 g574(.A(new_n772_), .B1(KEYINPUT114), .B2(KEYINPUT52), .C1(new_n749_), .C2(new_n313_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n771_), .A2(new_n775_), .A3(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT53), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT53), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n771_), .A2(new_n775_), .A3(new_n779_), .A4(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(G1339gat));
  XNOR2_X1  g580(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(new_n619_), .B2(new_n629_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n566_), .A2(new_n438_), .A3(new_n618_), .A4(new_n782_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n438_), .A2(new_n611_), .ZN(new_n788_));
  OAI21_X1  g587(.A(KEYINPUT55), .B1(new_n573_), .B2(KEYINPUT116), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n790_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n595_), .A2(new_n596_), .A3(new_n789_), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n573_), .A2(KEYINPUT55), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n791_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(KEYINPUT56), .A3(new_n572_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT56), .B1(new_n794_), .B2(new_n572_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n788_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n428_), .A2(new_n429_), .A3(KEYINPUT117), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT117), .B1(new_n428_), .B2(new_n429_), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n799_), .A2(new_n800_), .A3(new_n407_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n407_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n406_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n433_), .B1(new_n801_), .B2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n805_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n798_), .B1(new_n806_), .B2(KEYINPUT118), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT118), .ZN(new_n808_));
  AOI211_X1 g607(.A(new_n808_), .B(new_n805_), .C1(new_n614_), .C2(new_n615_), .ZN(new_n809_));
  OAI211_X1 g608(.A(KEYINPUT57), .B(new_n681_), .C1(new_n807_), .C2(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n611_), .A2(new_n805_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n811_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT58), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n794_), .A2(new_n572_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT56), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n795_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n818_), .A2(KEYINPUT58), .A3(new_n811_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n814_), .A2(new_n515_), .A3(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n810_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n681_), .B1(new_n807_), .B2(new_n809_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n821_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n787_), .B1(new_n824_), .B2(new_n660_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT59), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n400_), .A2(new_n389_), .A3(new_n648_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n825_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n805_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n830_));
  AOI22_X1  g629(.A1(new_n830_), .A2(new_n808_), .B1(new_n818_), .B2(new_n788_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n806_), .A2(KEYINPUT118), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n627_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n833_), .A2(KEYINPUT119), .A3(KEYINPUT57), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT119), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n835_), .B1(new_n823_), .B2(new_n822_), .ZN(new_n836_));
  NOR3_X1   g635(.A1(new_n834_), .A2(new_n836_), .A3(new_n821_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n787_), .B1(new_n837_), .B2(new_n660_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n838_), .A2(new_n827_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n828_), .B1(new_n839_), .B2(new_n826_), .ZN(new_n840_));
  OAI21_X1  g639(.A(G113gat), .B1(new_n840_), .B2(new_n438_), .ZN(new_n841_));
  INV_X1    g640(.A(G113gat), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n839_), .A2(new_n842_), .A3(new_n629_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(G1340gat));
  OAI21_X1  g643(.A(G120gat), .B1(new_n840_), .B2(new_n618_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n618_), .A2(KEYINPUT60), .ZN(new_n846_));
  MUX2_X1   g645(.A(new_n846_), .B(KEYINPUT60), .S(G120gat), .Z(new_n847_));
  NAND2_X1  g646(.A1(new_n839_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n845_), .A2(new_n848_), .ZN(G1341gat));
  OAI21_X1  g648(.A(G127gat), .B1(new_n840_), .B2(new_n565_), .ZN(new_n850_));
  INV_X1    g649(.A(G127gat), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n839_), .A2(new_n851_), .A3(new_n660_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(G1342gat));
  OAI21_X1  g652(.A(G134gat), .B1(new_n840_), .B2(new_n663_), .ZN(new_n854_));
  INV_X1    g653(.A(G134gat), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n839_), .A2(new_n855_), .A3(new_n627_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n856_), .ZN(G1343gat));
  OAI21_X1  g656(.A(KEYINPUT119), .B1(new_n833_), .B2(KEYINPUT57), .ZN(new_n858_));
  AND3_X1   g657(.A1(new_n814_), .A2(new_n515_), .A3(new_n819_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n859_), .B1(new_n833_), .B2(KEYINPUT57), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n823_), .A2(new_n835_), .A3(new_n822_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n858_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n786_), .B1(new_n862_), .B2(new_n565_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n312_), .A2(new_n637_), .A3(new_n648_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n863_), .A2(new_n396_), .A3(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n629_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n617_), .ZN(new_n868_));
  XOR2_X1   g667(.A(KEYINPUT120), .B(G148gat), .Z(new_n869_));
  XNOR2_X1  g668(.A(new_n868_), .B(new_n869_), .ZN(G1345gat));
  NAND2_X1  g669(.A1(new_n865_), .A2(new_n660_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(KEYINPUT61), .B(G155gat), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n871_), .B(new_n872_), .ZN(G1346gat));
  AOI21_X1  g672(.A(G162gat), .B1(new_n865_), .B2(new_n627_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n515_), .A2(G162gat), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(KEYINPUT121), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n874_), .B1(new_n865_), .B2(new_n876_), .ZN(G1347gat));
  NOR2_X1   g676(.A1(new_n399_), .A2(new_n401_), .ZN(new_n878_));
  XOR2_X1   g677(.A(new_n878_), .B(KEYINPUT122), .Z(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(new_n312_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n825_), .A2(new_n880_), .ZN(new_n881_));
  AOI211_X1 g680(.A(KEYINPUT62), .B(new_n207_), .C1(new_n881_), .C2(new_n629_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT62), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n629_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n883_), .B1(new_n884_), .B2(G169gat), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n881_), .A2(new_n322_), .A3(new_n629_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n882_), .B1(new_n885_), .B2(new_n886_), .ZN(G1348gat));
  AOI21_X1  g686(.A(G176gat), .B1(new_n881_), .B2(new_n617_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n838_), .A2(new_n880_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n889_), .A2(new_n208_), .A3(new_n618_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n888_), .A2(new_n890_), .ZN(G1349gat));
  NOR2_X1   g690(.A1(new_n889_), .A2(new_n565_), .ZN(new_n892_));
  OR2_X1    g691(.A1(new_n892_), .A2(KEYINPUT123), .ZN(new_n893_));
  AOI21_X1  g692(.A(G183gat), .B1(new_n892_), .B2(KEYINPUT123), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n565_), .A2(new_n318_), .ZN(new_n895_));
  AOI22_X1  g694(.A1(new_n893_), .A2(new_n894_), .B1(new_n881_), .B2(new_n895_), .ZN(G1350gat));
  NAND3_X1  g695(.A1(new_n881_), .A2(new_n218_), .A3(new_n627_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n881_), .A2(new_n515_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n898_), .B2(new_n215_), .ZN(G1351gat));
  NOR3_X1   g698(.A1(new_n399_), .A2(new_n390_), .A3(new_n244_), .ZN(new_n900_));
  AOI21_X1  g699(.A(KEYINPUT124), .B1(new_n838_), .B2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n902_));
  INV_X1    g701(.A(new_n900_), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n863_), .A2(new_n902_), .A3(new_n903_), .ZN(new_n904_));
  OAI211_X1 g703(.A(G197gat), .B(new_n629_), .C1(new_n901_), .C2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(KEYINPUT125), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n629_), .B1(new_n901_), .B2(new_n904_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(new_n252_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n838_), .A2(KEYINPUT124), .A3(new_n900_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n902_), .B1(new_n863_), .B2(new_n903_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT125), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n911_), .A2(new_n912_), .A3(G197gat), .A4(new_n629_), .ZN(new_n913_));
  AND3_X1   g712(.A1(new_n906_), .A2(new_n908_), .A3(new_n913_), .ZN(G1352gat));
  AOI21_X1  g713(.A(new_n618_), .B1(new_n909_), .B2(new_n910_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(G204gat), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n916_), .B1(new_n245_), .B2(new_n915_), .ZN(G1353gat));
  AOI21_X1  g716(.A(new_n565_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n911_), .A2(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(KEYINPUT126), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n919_), .B(new_n921_), .ZN(G1354gat));
  NAND2_X1  g721(.A1(new_n911_), .A2(new_n627_), .ZN(new_n923_));
  XOR2_X1   g722(.A(KEYINPUT127), .B(G218gat), .Z(new_n924_));
  NOR2_X1   g723(.A1(new_n663_), .A2(new_n924_), .ZN(new_n925_));
  AOI22_X1  g724(.A1(new_n923_), .A2(new_n924_), .B1(new_n911_), .B2(new_n925_), .ZN(G1355gat));
endmodule


