//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 1 0 0 1 1 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n622_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n805_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n820_, new_n821_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n865_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_;
  XOR2_X1   g000(.A(G85gat), .B(G92gat), .Z(new_n202_));
  NOR3_X1   g001(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT66), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT6), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n202_), .B1(new_n204_), .B2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT8), .ZN(new_n210_));
  XOR2_X1   g009(.A(KEYINPUT10), .B(G99gat), .Z(new_n211_));
  INV_X1    g010(.A(G106gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n214_));
  XOR2_X1   g013(.A(new_n214_), .B(KEYINPUT64), .Z(new_n215_));
  NAND2_X1  g014(.A1(KEYINPUT9), .A2(G85gat), .ZN(new_n216_));
  INV_X1    g015(.A(G92gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n218_), .B1(KEYINPUT9), .B2(G85gat), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n206_), .B(new_n213_), .C1(new_n215_), .C2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n210_), .A2(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(G29gat), .B(G36gat), .Z(new_n224_));
  XOR2_X1   g023(.A(G43gat), .B(G50gat), .Z(new_n225_));
  OR2_X1    g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n225_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(KEYINPUT15), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n223_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n228_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G232gat), .A2(G233gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT34), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT69), .B(KEYINPUT35), .ZN(new_n234_));
  OAI221_X1 g033(.A(new_n230_), .B1(new_n231_), .B2(new_n223_), .C1(new_n233_), .C2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n234_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G190gat), .B(G218gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G134gat), .B(G162gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n240_), .A2(KEYINPUT36), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n237_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(new_n240_), .B(KEYINPUT36), .Z(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n237_), .A2(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT37), .B1(new_n243_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT37), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n242_), .B(new_n248_), .C1(new_n237_), .C2(new_n245_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(G1gat), .ZN(new_n251_));
  INV_X1    g050(.A(G8gat), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT14), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n254_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G15gat), .B(G22gat), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(G1gat), .B(G8gat), .Z(new_n259_));
  XOR2_X1   g058(.A(new_n258_), .B(new_n259_), .Z(new_n260_));
  AND2_X1   g059(.A1(G231gat), .A2(G233gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G57gat), .B(G64gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT11), .ZN(new_n265_));
  XOR2_X1   g064(.A(G71gat), .B(G78gat), .Z(new_n266_));
  OR2_X1    g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n264_), .A2(KEYINPUT11), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n266_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n267_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n263_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT17), .ZN(new_n272_));
  XOR2_X1   g071(.A(G127gat), .B(G155gat), .Z(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT16), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G183gat), .B(G211gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  NOR3_X1   g075(.A1(new_n271_), .A2(new_n272_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n270_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n277_), .B1(new_n278_), .B2(new_n262_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT67), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n270_), .B(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n263_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n281_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n262_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n276_), .B(KEYINPUT17), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n282_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n279_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n250_), .A2(new_n288_), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n289_), .B(KEYINPUT71), .Z(new_n290_));
  NAND3_X1  g089(.A1(KEYINPUT78), .A2(G183gat), .A3(G190gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(KEYINPUT78), .B1(G183gat), .B2(G190gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT23), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(G183gat), .ZN(new_n295_));
  INV_X1    g094(.A(G190gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G183gat), .A2(G190gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT23), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n294_), .A2(new_n297_), .A3(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(G169gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT24), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n305_), .B1(G169gat), .B2(G176gat), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT75), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n307_), .B1(G169gat), .B2(G176gat), .ZN(new_n308_));
  INV_X1    g107(.A(G169gat), .ZN(new_n309_));
  INV_X1    g108(.A(G176gat), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(new_n310_), .A3(KEYINPUT75), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n306_), .A2(new_n308_), .A3(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT76), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n311_), .A2(new_n308_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n305_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT74), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT26), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n317_), .B1(new_n318_), .B2(G190gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT25), .B(G183gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT26), .B(G190gat), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n319_), .B(new_n320_), .C1(new_n321_), .C2(new_n317_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n314_), .A2(new_n316_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n298_), .A2(KEYINPUT23), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT77), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n298_), .A2(KEYINPUT77), .A3(KEYINPUT23), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n293_), .ZN(new_n329_));
  AOI21_X1  g128(.A(KEYINPUT23), .B1(new_n329_), .B2(new_n291_), .ZN(new_n330_));
  OAI22_X1  g129(.A1(new_n328_), .A2(new_n330_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n304_), .B1(new_n323_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(G197gat), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT87), .B1(new_n334_), .B2(G204gat), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT87), .ZN(new_n336_));
  INV_X1    g135(.A(G204gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(new_n337_), .A3(G197gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n334_), .A2(G204gat), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n335_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT21), .ZN(new_n341_));
  INV_X1    g140(.A(G218gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(G211gat), .ZN(new_n343_));
  INV_X1    g142(.A(G211gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(G218gat), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n341_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n340_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT89), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n340_), .A2(new_n346_), .A3(KEYINPUT89), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n334_), .A2(G204gat), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n337_), .A2(G197gat), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT21), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n343_), .A2(new_n345_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT88), .B(KEYINPUT21), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n354_), .B(new_n355_), .C1(new_n340_), .C2(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(KEYINPUT90), .B1(new_n351_), .B2(new_n357_), .ZN(new_n358_));
  AND3_X1   g157(.A1(new_n340_), .A2(KEYINPUT89), .A3(new_n346_), .ZN(new_n359_));
  AOI21_X1  g158(.A(KEYINPUT89), .B1(new_n340_), .B2(new_n346_), .ZN(new_n360_));
  OAI211_X1 g159(.A(KEYINPUT90), .B(new_n357_), .C1(new_n359_), .C2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n333_), .B1(new_n358_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT93), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n363_), .A2(new_n364_), .A3(KEYINPUT20), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n357_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT90), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n332_), .B1(new_n368_), .B2(new_n361_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT20), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT93), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G226gat), .A2(G233gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT19), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n297_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(new_n303_), .ZN(new_n375_));
  NOR3_X1   g174(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n376_), .B1(new_n321_), .B2(new_n320_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n377_), .A2(new_n300_), .A3(new_n294_), .A4(new_n312_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n375_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(new_n366_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n365_), .A2(new_n371_), .A3(new_n373_), .A4(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n373_), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT94), .B1(new_n379_), .B2(new_n366_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n366_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT94), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n384_), .A2(new_n385_), .A3(new_n375_), .A4(new_n378_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n383_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n368_), .A2(new_n332_), .A3(new_n361_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT20), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n382_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n381_), .A2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G8gat), .B(G36gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(KEYINPUT18), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G64gat), .B(G92gat), .ZN(new_n394_));
  XOR2_X1   g193(.A(new_n393_), .B(new_n394_), .Z(new_n395_));
  NAND2_X1  g194(.A1(new_n391_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT95), .ZN(new_n397_));
  INV_X1    g196(.A(new_n395_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n381_), .A2(new_n390_), .A3(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n396_), .A2(new_n397_), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT27), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n381_), .A2(KEYINPUT95), .A3(new_n390_), .A4(new_n398_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n400_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n365_), .A2(new_n371_), .A3(new_n382_), .A4(new_n380_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT91), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n366_), .B(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n406_), .A2(new_n379_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n373_), .B1(new_n407_), .B2(new_n389_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n404_), .A2(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(KEYINPUT98), .B1(new_n409_), .B2(new_n398_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT98), .ZN(new_n411_));
  AOI211_X1 g210(.A(new_n411_), .B(new_n395_), .C1(new_n404_), .C2(new_n408_), .ZN(new_n412_));
  OAI211_X1 g211(.A(KEYINPUT27), .B(new_n396_), .C1(new_n410_), .C2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n403_), .A2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(G155gat), .A2(G162gat), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT81), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G155gat), .A2(G162gat), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G141gat), .A2(G148gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT2), .ZN(new_n422_));
  NOR2_X1   g221(.A1(G141gat), .A2(G148gat), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT3), .B1(new_n424_), .B2(KEYINPUT82), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT82), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT3), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n423_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n422_), .A2(new_n425_), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n420_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n421_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n431_), .A2(new_n423_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n418_), .B(KEYINPUT1), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n432_), .B1(new_n417_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n430_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT29), .ZN(new_n436_));
  INV_X1    g235(.A(G233gat), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT85), .ZN(new_n438_));
  OR2_X1    g237(.A1(new_n438_), .A2(G228gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(G228gat), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n437_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT86), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n436_), .A2(new_n442_), .A3(new_n368_), .A4(new_n361_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n384_), .A2(KEYINPUT91), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n366_), .A2(new_n405_), .ZN(new_n445_));
  AOI22_X1  g244(.A1(new_n444_), .A2(new_n445_), .B1(KEYINPUT29), .B2(new_n435_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n443_), .B1(new_n446_), .B2(new_n442_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G78gat), .B(G106gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n406_), .A2(new_n436_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n442_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n448_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n452_), .A2(new_n453_), .A3(new_n443_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n449_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT92), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n456_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n457_));
  XOR2_X1   g256(.A(KEYINPUT84), .B(KEYINPUT28), .Z(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT83), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n460_), .B1(new_n435_), .B2(KEYINPUT29), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT29), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n430_), .A2(KEYINPUT83), .A3(new_n462_), .A4(new_n434_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G22gat), .B(G50gat), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  AND3_X1   g264(.A1(new_n461_), .A2(new_n463_), .A3(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n465_), .B1(new_n461_), .B2(new_n463_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n459_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n461_), .A2(new_n463_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(new_n464_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n461_), .A2(new_n463_), .A3(new_n465_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(new_n458_), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n468_), .A2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n455_), .B1(new_n457_), .B2(new_n473_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n468_), .A2(new_n472_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n475_), .A2(new_n456_), .A3(new_n449_), .A4(new_n454_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n414_), .A2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G71gat), .B(G99gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(G43gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT31), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G127gat), .B(G134gat), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  XOR2_X1   g282(.A(G113gat), .B(G120gat), .Z(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G113gat), .B(G120gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n482_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT79), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n485_), .A2(KEYINPUT79), .A3(new_n487_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n481_), .B(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G227gat), .A2(G233gat), .ZN(new_n494_));
  INV_X1    g293(.A(G15gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT30), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n493_), .B(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n332_), .B(KEYINPUT80), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n499_), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  AOI22_X1  g301(.A1(new_n490_), .A2(new_n491_), .B1(new_n430_), .B2(new_n434_), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n430_), .A2(new_n488_), .A3(new_n434_), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT4), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G225gat), .A2(G233gat), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n492_), .A2(new_n435_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT4), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n505_), .A2(new_n507_), .A3(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G1gat), .B(G29gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT96), .B(G85gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT0), .B(G57gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n506_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n511_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n516_), .B1(new_n511_), .B2(new_n517_), .ZN(new_n519_));
  OR2_X1    g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n502_), .A2(new_n520_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n478_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n477_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n516_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n503_), .A2(new_n504_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n524_), .B1(new_n525_), .B2(new_n507_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n505_), .A2(new_n510_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n526_), .B1(new_n527_), .B2(new_n507_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT33), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n519_), .A2(new_n529_), .ZN(new_n530_));
  AOI211_X1 g329(.A(KEYINPUT33), .B(new_n516_), .C1(new_n511_), .C2(new_n517_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n528_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n532_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT32), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n391_), .B1(new_n534_), .B2(new_n398_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n409_), .A2(KEYINPUT32), .A3(new_n395_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n535_), .A2(new_n536_), .A3(new_n520_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n523_), .B1(new_n533_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT97), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n520_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n541_));
  AND3_X1   g340(.A1(new_n403_), .A2(new_n413_), .A3(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  OAI211_X1 g342(.A(KEYINPUT97), .B(new_n523_), .C1(new_n533_), .C2(new_n537_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n540_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n522_), .B1(new_n545_), .B2(new_n502_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n228_), .B(KEYINPUT72), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n547_), .A2(new_n260_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G229gat), .A2(G233gat), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n229_), .A2(new_n260_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n547_), .B(new_n260_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n549_), .ZN(new_n553_));
  AOI22_X1  g352(.A1(new_n550_), .A2(new_n551_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G113gat), .B(G141gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G169gat), .B(G197gat), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n555_), .B(new_n556_), .Z(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(KEYINPUT73), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n554_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n554_), .A2(new_n559_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n283_), .A2(new_n210_), .A3(new_n222_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n223_), .A2(new_n281_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n566_), .A2(G230gat), .A3(G233gat), .ZN(new_n567_));
  XOR2_X1   g366(.A(KEYINPUT68), .B(KEYINPUT12), .Z(new_n568_));
  NAND2_X1  g367(.A1(new_n565_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G230gat), .A2(G233gat), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n223_), .A2(KEYINPUT12), .A3(new_n278_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n569_), .A2(new_n564_), .A3(new_n570_), .A4(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n567_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G120gat), .B(G148gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT5), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G176gat), .B(G204gat), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n575_), .B(new_n576_), .Z(new_n577_));
  OR2_X1    g376(.A1(new_n573_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n573_), .A2(new_n577_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT13), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n578_), .A2(KEYINPUT13), .A3(new_n579_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NOR4_X1   g383(.A1(new_n290_), .A2(new_n546_), .A3(new_n563_), .A4(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n585_), .A2(new_n251_), .A3(new_n520_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT38), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n243_), .A2(new_n246_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n546_), .A2(new_n589_), .ZN(new_n590_));
  NOR3_X1   g389(.A1(new_n584_), .A2(new_n563_), .A3(new_n287_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n520_), .ZN(new_n593_));
  OAI21_X1  g392(.A(G1gat), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n586_), .A2(new_n587_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n588_), .A2(new_n594_), .A3(new_n595_), .ZN(G1324gat));
  AND3_X1   g395(.A1(new_n585_), .A2(new_n252_), .A3(new_n414_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n590_), .A2(new_n414_), .A3(new_n591_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(G8gat), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT99), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT99), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n598_), .A2(new_n601_), .A3(G8gat), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT39), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT39), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n600_), .A2(new_n605_), .A3(new_n602_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n597_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n607_), .B(new_n609_), .ZN(G1325gat));
  INV_X1    g409(.A(new_n502_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n585_), .A2(new_n495_), .A3(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n590_), .A2(new_n611_), .A3(new_n591_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n613_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n614_));
  AOI21_X1  g413(.A(KEYINPUT41), .B1(new_n613_), .B2(G15gat), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n612_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT101), .Z(G1326gat));
  OAI21_X1  g416(.A(G22gat), .B1(new_n592_), .B2(new_n523_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(G22gat), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n585_), .A2(new_n621_), .A3(new_n477_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(G1327gat));
  NAND2_X1  g422(.A1(new_n545_), .A2(new_n502_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n522_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n584_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n589_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n628_), .A2(new_n288_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n626_), .A2(new_n562_), .A3(new_n627_), .A4(new_n629_), .ZN(new_n630_));
  NOR3_X1   g429(.A1(new_n630_), .A2(G29gat), .A3(new_n593_), .ZN(new_n631_));
  AOI21_X1  g430(.A(KEYINPUT103), .B1(new_n247_), .B2(new_n249_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n247_), .A2(new_n249_), .A3(KEYINPUT103), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(KEYINPUT43), .B1(new_n546_), .B2(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n250_), .A2(KEYINPUT43), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n542_), .B1(new_n539_), .B2(new_n538_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n611_), .B1(new_n638_), .B2(new_n544_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n637_), .B1(new_n639_), .B2(new_n522_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n636_), .A2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n627_), .A2(new_n562_), .A3(new_n287_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(KEYINPUT44), .B1(new_n641_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT44), .ZN(new_n645_));
  AOI211_X1 g444(.A(new_n645_), .B(new_n642_), .C1(new_n636_), .C2(new_n640_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(new_n520_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n631_), .B1(new_n648_), .B2(G29gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT104), .ZN(G1328gat));
  NAND2_X1  g449(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n651_));
  NOR2_X1   g450(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n414_), .B(KEYINPUT106), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n653_), .A2(G36gat), .ZN(new_n654_));
  OR3_X1    g453(.A1(new_n630_), .A2(KEYINPUT45), .A3(new_n654_), .ZN(new_n655_));
  OAI21_X1  g454(.A(KEYINPUT45), .B1(new_n630_), .B2(new_n654_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n652_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT105), .B1(new_n647_), .B2(new_n414_), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n247_), .A2(new_n249_), .A3(KEYINPUT103), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n659_), .A2(new_n632_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n660_), .B1(new_n639_), .B2(new_n522_), .ZN(new_n661_));
  AOI22_X1  g460(.A1(new_n661_), .A2(KEYINPUT43), .B1(new_n626_), .B2(new_n637_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n645_), .B1(new_n662_), .B2(new_n642_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n641_), .A2(KEYINPUT44), .A3(new_n643_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n663_), .A2(KEYINPUT105), .A3(new_n414_), .A4(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(G36gat), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n651_), .B(new_n657_), .C1(new_n658_), .C2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n663_), .A2(new_n414_), .A3(new_n664_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT105), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n671_), .A2(G36gat), .A3(new_n665_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n651_), .B1(new_n672_), .B2(new_n657_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n668_), .A2(new_n673_), .ZN(G1329gat));
  NOR3_X1   g473(.A1(new_n630_), .A2(G43gat), .A3(new_n502_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n647_), .A2(new_n611_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n676_), .B2(G43gat), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g477(.A1(new_n647_), .A2(G50gat), .A3(new_n477_), .ZN(new_n679_));
  INV_X1    g478(.A(G50gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n680_), .B1(new_n630_), .B2(new_n523_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n679_), .A2(new_n681_), .ZN(G1331gat));
  NOR2_X1   g481(.A1(new_n290_), .A2(new_n627_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n546_), .A2(new_n562_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n686_), .A2(KEYINPUT108), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(KEYINPUT108), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(new_n520_), .A3(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(G57gat), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n287_), .A2(new_n562_), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n590_), .A2(new_n584_), .A3(new_n691_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n593_), .A2(new_n690_), .ZN(new_n693_));
  AOI22_X1  g492(.A1(new_n689_), .A2(new_n690_), .B1(new_n692_), .B2(new_n693_), .ZN(G1332gat));
  INV_X1    g493(.A(G64gat), .ZN(new_n695_));
  INV_X1    g494(.A(new_n653_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n692_), .B2(new_n696_), .ZN(new_n697_));
  XOR2_X1   g496(.A(new_n697_), .B(KEYINPUT48), .Z(new_n698_));
  NOR2_X1   g497(.A1(new_n653_), .A2(G64gat), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT109), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n698_), .B1(new_n685_), .B2(new_n700_), .ZN(G1333gat));
  INV_X1    g500(.A(G71gat), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n702_), .B1(new_n692_), .B2(new_n611_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT49), .Z(new_n704_));
  NAND3_X1  g503(.A1(new_n686_), .A2(new_n702_), .A3(new_n611_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1334gat));
  INV_X1    g505(.A(G78gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n707_), .B1(new_n692_), .B2(new_n477_), .ZN(new_n708_));
  XOR2_X1   g507(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n709_));
  XNOR2_X1  g508(.A(new_n708_), .B(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n477_), .A2(new_n707_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n710_), .B1(new_n685_), .B2(new_n711_), .ZN(G1335gat));
  NAND3_X1  g511(.A1(new_n684_), .A2(new_n584_), .A3(new_n629_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n713_), .A2(G85gat), .A3(new_n593_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n288_), .A2(new_n562_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n641_), .A2(new_n584_), .A3(new_n715_), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n716_), .A2(new_n593_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n714_), .B1(new_n717_), .B2(G85gat), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT111), .Z(G1336gat));
  INV_X1    g518(.A(new_n713_), .ZN(new_n720_));
  AOI21_X1  g519(.A(G92gat), .B1(new_n720_), .B2(new_n414_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT112), .Z(new_n722_));
  NOR3_X1   g521(.A1(new_n716_), .A2(new_n217_), .A3(new_n653_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1337gat));
  OAI21_X1  g523(.A(G99gat), .B1(new_n716_), .B2(new_n502_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n720_), .A2(new_n611_), .A3(new_n211_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g527(.A1(new_n720_), .A2(new_n212_), .A3(new_n477_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G106gat), .B1(new_n716_), .B2(new_n523_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n730_), .A2(KEYINPUT52), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n730_), .A2(KEYINPUT52), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n729_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT53), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT53), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n735_), .B(new_n729_), .C1(new_n731_), .C2(new_n732_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(G1339gat));
  NAND2_X1  g536(.A1(new_n572_), .A2(KEYINPUT113), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT55), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT55), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n572_), .A2(KEYINPUT113), .A3(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n569_), .A2(new_n564_), .A3(new_n571_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n742_), .A2(G230gat), .A3(G233gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n739_), .A2(new_n741_), .A3(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n577_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT56), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT115), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n744_), .A2(KEYINPUT56), .A3(new_n577_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n747_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n552_), .A2(new_n549_), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n548_), .A2(new_n553_), .A3(new_n551_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n558_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n753_), .B1(new_n558_), .B2(new_n554_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n578_), .A2(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT56), .B1(new_n744_), .B2(new_n577_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(KEYINPUT115), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n750_), .A2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT58), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n250_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n750_), .A2(new_n757_), .A3(KEYINPUT58), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT116), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT116), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n750_), .A2(new_n757_), .A3(new_n763_), .A4(KEYINPUT58), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n760_), .A2(new_n762_), .A3(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT117), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n562_), .A2(new_n578_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n767_), .B1(new_n747_), .B2(new_n749_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n580_), .A2(new_n754_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n628_), .B1(new_n768_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n766_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n765_), .B1(KEYINPUT57), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT57), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n744_), .A2(KEYINPUT56), .A3(new_n577_), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n562_), .B(new_n578_), .C1(new_n776_), .C2(new_n756_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n589_), .B1(new_n777_), .B2(new_n769_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT117), .B1(new_n778_), .B2(KEYINPUT114), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n771_), .A2(new_n766_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n775_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n287_), .B1(new_n774_), .B2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n627_), .A2(new_n250_), .A3(new_n691_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT54), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n414_), .A2(new_n502_), .A3(new_n477_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n785_), .A2(new_n520_), .A3(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(G113gat), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(new_n789_), .A3(new_n562_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT59), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n787_), .A2(new_n791_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n785_), .A2(KEYINPUT59), .A3(new_n520_), .A4(new_n786_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n563_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n790_), .B1(new_n794_), .B2(new_n789_), .ZN(G1340gat));
  INV_X1    g594(.A(KEYINPUT60), .ZN(new_n796_));
  AOI21_X1  g595(.A(G120gat), .B1(new_n584_), .B2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n797_), .B1(new_n796_), .B2(G120gat), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n785_), .A2(new_n520_), .A3(new_n786_), .A4(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT118), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n799_), .B(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n627_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n802_));
  INV_X1    g601(.A(G120gat), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n801_), .B1(new_n802_), .B2(new_n803_), .ZN(G1341gat));
  INV_X1    g603(.A(G127gat), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n788_), .A2(new_n805_), .A3(new_n288_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n287_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n807_), .B2(new_n805_), .ZN(G1342gat));
  AOI21_X1  g607(.A(G134gat), .B1(new_n788_), .B2(new_n589_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n792_), .A2(new_n793_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n250_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(G134gat), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(KEYINPUT119), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n809_), .B1(new_n810_), .B2(new_n813_), .ZN(G1343gat));
  NOR3_X1   g613(.A1(new_n696_), .A2(new_n611_), .A3(new_n523_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  AOI211_X1 g615(.A(new_n593_), .B(new_n816_), .C1(new_n782_), .C2(new_n784_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n562_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n584_), .ZN(new_n820_));
  XOR2_X1   g619(.A(KEYINPUT120), .B(G148gat), .Z(new_n821_));
  XNOR2_X1  g620(.A(new_n820_), .B(new_n821_), .ZN(G1345gat));
  XNOR2_X1  g621(.A(KEYINPUT61), .B(G155gat), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT121), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n825_), .B1(new_n817_), .B2(new_n288_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n785_), .A2(new_n520_), .A3(new_n288_), .A4(new_n815_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n827_), .A2(KEYINPUT121), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n824_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n817_), .A2(new_n825_), .A3(new_n288_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n827_), .A2(KEYINPUT121), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n830_), .A2(new_n831_), .A3(new_n823_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n829_), .A2(new_n832_), .ZN(G1346gat));
  AOI21_X1  g632(.A(G162gat), .B1(new_n817_), .B2(new_n589_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n660_), .A2(G162gat), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n817_), .B2(new_n835_), .ZN(G1347gat));
  AOI21_X1  g635(.A(new_n653_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT22), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n521_), .A2(new_n523_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n837_), .A2(new_n838_), .A3(new_n562_), .A4(new_n840_), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n841_), .A2(KEYINPUT62), .A3(new_n309_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(KEYINPUT62), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n837_), .A2(new_n562_), .A3(new_n840_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT62), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n309_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n842_), .B1(new_n843_), .B2(new_n846_), .ZN(G1348gat));
  AOI211_X1 g646(.A(new_n653_), .B(new_n839_), .C1(new_n782_), .C2(new_n784_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n584_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g649(.A1(new_n785_), .A2(new_n696_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n851_), .A2(new_n287_), .A3(new_n839_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n295_), .A2(KEYINPUT122), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(new_n320_), .A3(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(KEYINPUT122), .A2(G183gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n852_), .B2(new_n855_), .ZN(G1350gat));
  NAND2_X1  g655(.A1(new_n589_), .A2(new_n321_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(KEYINPUT123), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n848_), .A2(new_n858_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n851_), .A2(new_n250_), .A3(new_n839_), .ZN(new_n860_));
  OAI211_X1 g659(.A(KEYINPUT124), .B(new_n859_), .C1(new_n860_), .C2(new_n296_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT124), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n296_), .B1(new_n848_), .B2(new_n811_), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n837_), .A2(new_n840_), .A3(new_n858_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n862_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n861_), .A2(new_n865_), .ZN(G1351gat));
  AND2_X1   g665(.A1(new_n541_), .A2(new_n502_), .ZN(new_n867_));
  AND3_X1   g666(.A1(new_n785_), .A2(new_n696_), .A3(new_n867_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n868_), .A2(KEYINPUT125), .A3(G197gat), .A4(new_n562_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT125), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n837_), .A2(new_n562_), .A3(new_n867_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n871_), .B2(new_n334_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n334_), .ZN(new_n873_));
  AND3_X1   g672(.A1(new_n869_), .A2(new_n872_), .A3(new_n873_), .ZN(G1352gat));
  NAND2_X1  g673(.A1(new_n868_), .A2(new_n584_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT126), .B(G204gat), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n875_), .B(new_n876_), .ZN(G1353gat));
  AOI21_X1  g676(.A(new_n287_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n868_), .A2(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(KEYINPUT127), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n879_), .B(new_n882_), .ZN(G1354gat));
  NAND3_X1  g682(.A1(new_n868_), .A2(new_n342_), .A3(new_n589_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n868_), .A2(new_n811_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(new_n342_), .ZN(G1355gat));
endmodule


