//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 0 0 1 0 1 0 0 1 1 1 0 1 0 0 1 1 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_;
  INV_X1    g000(.A(KEYINPUT66), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT10), .B(G99gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT64), .B1(new_n203_), .B2(G106gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n205_));
  INV_X1    g004(.A(G106gat), .ZN(new_n206_));
  INV_X1    g005(.A(G99gat), .ZN(new_n207_));
  AND2_X1   g006(.A1(new_n207_), .A2(KEYINPUT10), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(KEYINPUT10), .ZN(new_n209_));
  OAI211_X1 g008(.A(new_n205_), .B(new_n206_), .C1(new_n208_), .C2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n204_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  AND2_X1   g015(.A1(G85gat), .A2(G92gat), .ZN(new_n217_));
  OR2_X1    g016(.A1(G85gat), .A2(G92gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT9), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n217_), .B1(new_n218_), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G85gat), .A2(G92gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n220_), .B1(new_n223_), .B2(new_n219_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n216_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n202_), .B1(new_n211_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT7), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(new_n207_), .A3(new_n206_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n228_), .A2(new_n214_), .A3(new_n215_), .A4(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(G85gat), .A2(G92gat), .ZN(new_n231_));
  NOR3_X1   g030(.A1(new_n217_), .A2(new_n231_), .A3(KEYINPUT67), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT8), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT8), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n230_), .A2(new_n235_), .A3(new_n232_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n214_), .A2(new_n215_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n224_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n223_), .B1(new_n231_), .B2(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n238_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n242_), .A2(KEYINPUT66), .A3(new_n204_), .A4(new_n210_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n226_), .A2(new_n237_), .A3(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT68), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n226_), .A2(new_n237_), .A3(new_n246_), .A4(new_n243_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT69), .B(G71gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(G78gat), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(G57gat), .B(G64gat), .Z(new_n252_));
  INV_X1    g051(.A(KEYINPUT11), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n252_), .A2(new_n253_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n251_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n250_), .A2(new_n254_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n226_), .A2(KEYINPUT70), .A3(new_n243_), .ZN(new_n260_));
  AOI21_X1  g059(.A(KEYINPUT70), .B1(new_n226_), .B2(new_n243_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n237_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT12), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n259_), .A2(new_n263_), .ZN(new_n264_));
  AOI22_X1  g063(.A1(new_n248_), .A2(new_n259_), .B1(new_n262_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G230gat), .A2(G233gat), .ZN(new_n266_));
  AND2_X1   g065(.A1(new_n257_), .A2(new_n258_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n245_), .A2(new_n247_), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(new_n263_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n265_), .A2(new_n266_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n248_), .A2(new_n259_), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n271_), .A2(new_n268_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n270_), .B1(new_n266_), .B2(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(G120gat), .B(G148gat), .Z(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(G204gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT5), .ZN(new_n276_));
  INV_X1    g075(.A(G176gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n273_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n273_), .A2(new_n279_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n273_), .A2(KEYINPUT71), .A3(new_n279_), .ZN(new_n284_));
  AND2_X1   g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n285_), .A2(KEYINPUT13), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(KEYINPUT13), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT72), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G229gat), .A2(G233gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G29gat), .B(G36gat), .ZN(new_n293_));
  INV_X1    g092(.A(G43gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G50gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n293_), .B(G43gat), .ZN(new_n297_));
  INV_X1    g096(.A(G50gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT78), .ZN(new_n302_));
  INV_X1    g101(.A(G1gat), .ZN(new_n303_));
  INV_X1    g102(.A(G8gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT14), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT75), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n306_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G15gat), .B(G22gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(G1gat), .B(G8gat), .Z(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT78), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n300_), .A2(new_n314_), .ZN(new_n315_));
  AND3_X1   g114(.A1(new_n302_), .A2(new_n313_), .A3(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n313_), .B1(new_n302_), .B2(new_n315_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n292_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n302_), .A2(new_n315_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n312_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT15), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n300_), .B(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(new_n313_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n320_), .A2(new_n323_), .A3(new_n291_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G113gat), .B(G141gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(G197gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT79), .ZN(new_n327_));
  INV_X1    g126(.A(G169gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n318_), .A2(new_n324_), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT80), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT80), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n318_), .A2(new_n324_), .A3(new_n332_), .A4(new_n329_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n318_), .A2(new_n324_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n329_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n334_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G155gat), .A2(G162gat), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT86), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(KEYINPUT86), .A2(G155gat), .A3(G162gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  OR2_X1    g142(.A1(G155gat), .A2(G162gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT87), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n343_), .A2(KEYINPUT87), .A3(new_n344_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(G141gat), .A2(G148gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT3), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G141gat), .A2(G148gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT2), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n347_), .A2(new_n348_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n343_), .A2(KEYINPUT1), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT1), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n341_), .A2(new_n355_), .A3(new_n342_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n354_), .A2(new_n344_), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n349_), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n353_), .B1(new_n359_), .B2(new_n351_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT29), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G22gat), .B(G50gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT28), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n360_), .A2(new_n361_), .A3(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n363_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n357_), .A2(new_n358_), .A3(new_n351_), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n347_), .A2(new_n348_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n350_), .A2(new_n352_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n366_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n365_), .B1(new_n369_), .B2(KEYINPUT29), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n364_), .A2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G197gat), .B(G204gat), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT21), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT88), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n373_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G211gat), .B(G218gat), .ZN(new_n377_));
  OR2_X1    g176(.A1(new_n377_), .A2(KEYINPUT89), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n372_), .A2(new_n373_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(KEYINPUT89), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n378_), .A2(KEYINPUT90), .A3(new_n379_), .A4(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n378_), .A2(new_n380_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(KEYINPUT90), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n376_), .A2(new_n381_), .A3(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n385_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n386_));
  INV_X1    g185(.A(G228gat), .ZN(new_n387_));
  INV_X1    g186(.A(G233gat), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n386_), .A2(new_n389_), .ZN(new_n390_));
  OAI221_X1 g189(.A(new_n385_), .B1(new_n387_), .B2(new_n388_), .C1(new_n360_), .C2(new_n361_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G78gat), .B(G106gat), .ZN(new_n393_));
  XOR2_X1   g192(.A(new_n393_), .B(KEYINPUT91), .Z(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  OAI211_X1 g194(.A(KEYINPUT92), .B(new_n371_), .C1(new_n392_), .C2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n371_), .A2(KEYINPUT92), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n397_), .A2(new_n394_), .A3(new_n390_), .A4(new_n391_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n392_), .A2(new_n395_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n396_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n392_), .A2(new_n395_), .A3(new_n371_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT93), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G71gat), .B(G99gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G227gat), .A2(G233gat), .ZN(new_n405_));
  XOR2_X1   g204(.A(new_n404_), .B(new_n405_), .Z(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT85), .ZN(new_n408_));
  XOR2_X1   g207(.A(G127gat), .B(G134gat), .Z(new_n409_));
  INV_X1    g208(.A(G113gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G127gat), .B(G134gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(G113gat), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n411_), .A2(G120gat), .A3(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(G120gat), .B1(new_n411_), .B2(new_n413_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n408_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n411_), .A2(new_n413_), .ZN(new_n417_));
  INV_X1    g216(.A(G120gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n411_), .A2(G120gat), .A3(new_n413_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(KEYINPUT85), .A3(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n416_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT30), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G183gat), .A2(G190gat), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT82), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT23), .ZN(new_n428_));
  NOR2_X1   g227(.A1(G183gat), .A2(G190gat), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT23), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n425_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n428_), .A2(new_n430_), .A3(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT84), .B(G176gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT22), .B(G169gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G169gat), .A2(G176gat), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n433_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n427_), .A2(new_n431_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT83), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n425_), .A2(KEYINPUT23), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT83), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n427_), .A2(new_n443_), .A3(new_n431_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n441_), .A2(new_n442_), .A3(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n328_), .A2(new_n277_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n446_), .A2(KEYINPUT24), .ZN(new_n447_));
  XNOR2_X1  g246(.A(KEYINPUT25), .B(G183gat), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(G190gat), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n450_), .A2(KEYINPUT81), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n449_), .B1(KEYINPUT26), .B2(new_n451_), .ZN(new_n452_));
  OR3_X1    g251(.A1(new_n450_), .A2(KEYINPUT81), .A3(KEYINPUT26), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n447_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n446_), .A2(KEYINPUT24), .A3(new_n437_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n445_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n424_), .A2(new_n439_), .A3(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n422_), .B(KEYINPUT30), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n439_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G15gat), .B(G43gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT31), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n457_), .A2(new_n460_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n463_), .B1(new_n457_), .B2(new_n460_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n407_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n466_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(new_n406_), .A3(new_n464_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G225gat), .A2(G233gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT97), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT4), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n414_), .A2(new_n415_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n360_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n369_), .A2(new_n421_), .A3(new_n416_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n474_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  AND2_X1   g277(.A1(new_n416_), .A2(new_n421_), .ZN(new_n479_));
  AOI21_X1  g278(.A(KEYINPUT4), .B1(new_n479_), .B2(new_n369_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n473_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n476_), .A2(new_n477_), .A3(new_n471_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT0), .B(G57gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(G85gat), .ZN(new_n484_));
  XOR2_X1   g283(.A(G1gat), .B(G29gat), .Z(new_n485_));
  XOR2_X1   g284(.A(new_n484_), .B(new_n485_), .Z(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n481_), .A2(new_n482_), .A3(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n487_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n470_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n376_), .A2(new_n381_), .A3(new_n384_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n456_), .A2(new_n493_), .A3(new_n439_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT26), .B(G190gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n448_), .A2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n428_), .A2(new_n432_), .A3(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n437_), .A2(KEYINPUT24), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n446_), .B1(new_n498_), .B2(KEYINPUT94), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n499_), .B1(KEYINPUT94), .B2(new_n498_), .ZN(new_n500_));
  NOR3_X1   g299(.A1(new_n497_), .A2(new_n500_), .A3(new_n447_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n445_), .A2(new_n430_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n501_), .B1(new_n502_), .B2(new_n438_), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n494_), .B(KEYINPUT20), .C1(new_n503_), .C2(new_n493_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G226gat), .A2(G233gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT19), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT20), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n508_), .B1(new_n459_), .B2(new_n385_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n503_), .A2(new_n493_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n506_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n509_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n507_), .A2(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(G8gat), .B(G36gat), .Z(new_n514_));
  XNOR2_X1  g313(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G64gat), .B(G92gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n513_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT96), .ZN(new_n520_));
  INV_X1    g319(.A(new_n518_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n507_), .A2(new_n512_), .A3(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n519_), .A2(new_n520_), .A3(new_n522_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n507_), .A2(new_n512_), .A3(KEYINPUT96), .A4(new_n521_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT27), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n502_), .A2(new_n438_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT99), .ZN(new_n528_));
  INV_X1    g327(.A(new_n501_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n527_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n438_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n531_), .B1(new_n445_), .B2(new_n430_), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT99), .B1(new_n532_), .B2(new_n501_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n530_), .A2(new_n493_), .A3(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n511_), .B1(new_n534_), .B2(new_n509_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n504_), .A2(new_n506_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n518_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT101), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n538_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n539_), .A2(KEYINPUT27), .A3(new_n522_), .A4(new_n540_), .ZN(new_n541_));
  AND4_X1   g340(.A1(new_n403_), .A2(new_n492_), .A3(new_n526_), .A4(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n521_), .A2(KEYINPUT32), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n544_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n507_), .A2(new_n512_), .A3(new_n543_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n545_), .B(new_n546_), .C1(new_n488_), .C2(new_n489_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n476_), .A2(new_n477_), .A3(new_n473_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(new_n486_), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n550_), .A2(KEYINPUT98), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n471_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(KEYINPUT98), .ZN(new_n553_));
  AND3_X1   g352(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n554_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n481_), .A2(new_n482_), .A3(new_n487_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT33), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n548_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n402_), .A2(KEYINPUT93), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT93), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n560_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(KEYINPUT100), .B1(new_n558_), .B2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n523_), .A2(new_n524_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n554_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n564_), .A2(new_n557_), .A3(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(new_n547_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT100), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(new_n403_), .A3(new_n568_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n562_), .A2(new_n490_), .A3(new_n526_), .A4(new_n541_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n563_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n542_), .B1(new_n571_), .B2(new_n470_), .ZN(new_n572_));
  XOR2_X1   g371(.A(G127gat), .B(G155gat), .Z(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT77), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G183gat), .B(G211gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n576_), .B(new_n577_), .Z(new_n578_));
  XOR2_X1   g377(.A(new_n578_), .B(KEYINPUT17), .Z(new_n579_));
  XNOR2_X1  g378(.A(new_n259_), .B(new_n312_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G231gat), .A2(G233gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n579_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n578_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n582_), .A2(KEYINPUT17), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT36), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(G134gat), .ZN(new_n589_));
  INV_X1    g388(.A(G162gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT34), .ZN(new_n594_));
  AOI22_X1  g393(.A1(new_n322_), .A2(new_n262_), .B1(new_n248_), .B2(new_n301_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT73), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n594_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n262_), .A2(new_n322_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n248_), .A2(new_n301_), .ZN(new_n599_));
  AND4_X1   g398(.A1(new_n596_), .A2(new_n598_), .A3(new_n599_), .A4(new_n594_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n593_), .B1(new_n597_), .B2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n598_), .A2(new_n599_), .ZN(new_n602_));
  OAI21_X1  g401(.A(KEYINPUT34), .B1(new_n602_), .B2(KEYINPUT73), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n595_), .A2(new_n596_), .A3(new_n594_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n603_), .A2(new_n604_), .A3(new_n592_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT35), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n601_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  AOI22_X1  g406(.A1(new_n601_), .A2(new_n605_), .B1(new_n606_), .B2(new_n595_), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n587_), .B(new_n591_), .C1(new_n607_), .C2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n601_), .A2(new_n605_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n595_), .A2(new_n606_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n591_), .A2(new_n587_), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n591_), .A2(new_n587_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n601_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n612_), .A2(new_n613_), .A3(new_n614_), .A4(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(KEYINPUT74), .B(KEYINPUT37), .ZN(new_n617_));
  AND3_X1   g416(.A1(new_n609_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(KEYINPUT74), .A2(KEYINPUT37), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n619_), .B1(new_n609_), .B2(new_n616_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n572_), .A2(new_n586_), .A3(new_n621_), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n290_), .A2(new_n338_), .A3(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n623_), .A2(new_n303_), .A3(new_n491_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT38), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n572_), .A2(new_n586_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n288_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n338_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n609_), .A2(new_n616_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n626_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G1gat), .B1(new_n631_), .B2(new_n490_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n625_), .A2(new_n632_), .ZN(G1324gat));
  AND2_X1   g432(.A1(new_n541_), .A2(new_n526_), .ZN(new_n634_));
  OAI21_X1  g433(.A(G8gat), .B1(new_n631_), .B2(new_n634_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n635_), .A2(KEYINPUT102), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(KEYINPUT102), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(KEYINPUT39), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n634_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n623_), .A2(new_n304_), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT39), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n635_), .A2(KEYINPUT102), .A3(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n638_), .A2(new_n640_), .A3(new_n642_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g443(.A(G15gat), .B1(new_n631_), .B2(new_n470_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT41), .Z(new_n646_));
  INV_X1    g445(.A(G15gat), .ZN(new_n647_));
  INV_X1    g446(.A(new_n470_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n623_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n649_), .ZN(G1326gat));
  OAI21_X1  g449(.A(G22gat), .B1(new_n631_), .B2(new_n403_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT42), .ZN(new_n652_));
  INV_X1    g451(.A(G22gat), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n623_), .A2(new_n653_), .A3(new_n562_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(G1327gat));
  NAND2_X1  g454(.A1(new_n629_), .A2(new_n586_), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n656_), .A2(new_n630_), .A3(new_n572_), .ZN(new_n657_));
  AOI21_X1  g456(.A(G29gat), .B1(new_n657_), .B2(new_n491_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT105), .ZN(new_n659_));
  INV_X1    g458(.A(new_n621_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n572_), .A2(new_n660_), .A3(KEYINPUT43), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT104), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT103), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n572_), .A2(new_n663_), .ZN(new_n664_));
  AOI211_X1 g463(.A(KEYINPUT103), .B(new_n542_), .C1(new_n571_), .C2(new_n470_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n664_), .A2(new_n665_), .A3(new_n660_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT43), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n662_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n571_), .A2(new_n470_), .ZN(new_n669_));
  OAI21_X1  g468(.A(KEYINPUT103), .B1(new_n669_), .B2(new_n542_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n572_), .A2(new_n663_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n670_), .A2(new_n621_), .A3(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n672_), .A2(KEYINPUT104), .A3(KEYINPUT43), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n661_), .B1(new_n668_), .B2(new_n673_), .ZN(new_n674_));
  OAI211_X1 g473(.A(new_n659_), .B(KEYINPUT44), .C1(new_n674_), .C2(new_n656_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n661_), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n666_), .A2(new_n662_), .A3(new_n667_), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT104), .B1(new_n672_), .B2(KEYINPUT43), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n676_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n656_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n659_), .A2(KEYINPUT44), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n659_), .A2(KEYINPUT44), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n679_), .A2(new_n680_), .A3(new_n681_), .A4(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n490_), .B1(new_n675_), .B2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n658_), .B1(new_n684_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g484(.A(G36gat), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n657_), .A2(new_n686_), .A3(new_n639_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT45), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n634_), .B1(new_n675_), .B2(new_n683_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(new_n686_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT107), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n690_), .B(new_n692_), .Z(G1329gat));
  NAND3_X1  g492(.A1(new_n657_), .A2(new_n294_), .A3(new_n648_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n470_), .B1(new_n675_), .B2(new_n683_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n694_), .B1(new_n695_), .B2(new_n294_), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g496(.A(G50gat), .B1(new_n657_), .B2(new_n562_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n298_), .B1(new_n675_), .B2(new_n683_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n699_), .B2(new_n562_), .ZN(G1331gat));
  AND4_X1   g499(.A1(new_n630_), .A2(new_n289_), .A3(new_n628_), .A4(new_n626_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n701_), .A2(G57gat), .A3(new_n491_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT108), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n288_), .A2(new_n338_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n622_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G57gat), .B1(new_n706_), .B2(new_n491_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n703_), .A2(new_n707_), .ZN(G1332gat));
  INV_X1    g507(.A(G64gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n701_), .B2(new_n639_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT48), .Z(new_n711_));
  NAND3_X1  g510(.A1(new_n706_), .A2(new_n709_), .A3(new_n639_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1333gat));
  INV_X1    g512(.A(G71gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n714_), .B1(new_n701_), .B2(new_n648_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT49), .Z(new_n716_));
  NAND3_X1  g515(.A1(new_n706_), .A2(new_n714_), .A3(new_n648_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1334gat));
  NAND2_X1  g517(.A1(new_n701_), .A2(new_n562_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(G78gat), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT50), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n705_), .A2(G78gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n403_), .B2(new_n722_), .ZN(G1335gat));
  INV_X1    g522(.A(new_n586_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n724_), .A2(new_n338_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  NOR4_X1   g525(.A1(new_n290_), .A2(new_n630_), .A3(new_n572_), .A4(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(G85gat), .B1(new_n727_), .B2(new_n491_), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n674_), .A2(new_n288_), .A3(new_n726_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n730_), .A2(new_n490_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n728_), .B1(new_n731_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g531(.A(G92gat), .B1(new_n727_), .B2(new_n639_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n730_), .A2(new_n634_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n734_), .B2(G92gat), .ZN(G1337gat));
  NAND4_X1  g534(.A1(new_n679_), .A2(new_n627_), .A3(new_n648_), .A4(new_n725_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(G99gat), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n727_), .B(new_n648_), .C1(new_n208_), .C2(new_n209_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT109), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT109), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n737_), .A2(new_n741_), .A3(new_n738_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g543(.A(KEYINPUT52), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n679_), .A2(new_n627_), .A3(new_n562_), .A4(new_n725_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT110), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n746_), .A2(new_n747_), .A3(G106gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n746_), .B2(G106gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n745_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n746_), .A2(G106gat), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT110), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n746_), .A2(new_n747_), .A3(G106gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(KEYINPUT52), .A3(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n727_), .A2(new_n206_), .A3(new_n562_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n750_), .A2(new_n754_), .A3(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT53), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT53), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n750_), .A2(new_n754_), .A3(new_n758_), .A4(new_n755_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(G1339gat));
  INV_X1    g559(.A(KEYINPUT119), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n266_), .B1(new_n265_), .B2(new_n269_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT55), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n270_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n265_), .A2(KEYINPUT55), .A3(new_n266_), .A4(new_n269_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n766_), .A2(KEYINPUT56), .A3(new_n279_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT113), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n262_), .A2(new_n264_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n269_), .A2(new_n271_), .A3(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n266_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n763_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n771_), .A2(new_n772_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n765_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n279_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT112), .ZN(new_n778_));
  XOR2_X1   g577(.A(KEYINPUT111), .B(KEYINPUT56), .Z(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n777_), .A2(new_n778_), .A3(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n278_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n782_));
  OAI21_X1  g581(.A(KEYINPUT112), .B1(new_n782_), .B2(new_n779_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n782_), .A2(KEYINPUT113), .A3(KEYINPUT56), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n769_), .A2(new_n781_), .A3(new_n783_), .A4(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n785_), .A2(new_n338_), .A3(new_n280_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n291_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n320_), .A2(new_n323_), .A3(new_n292_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n788_), .A3(new_n336_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n334_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n285_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n786_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(new_n630_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT57), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(KEYINPUT114), .A3(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT114), .ZN(new_n796_));
  INV_X1    g595(.A(new_n630_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n797_), .B1(new_n786_), .B2(new_n791_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n796_), .B1(new_n798_), .B2(KEYINPUT57), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n795_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT115), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n801_), .B1(new_n782_), .B2(KEYINPUT56), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT56), .ZN(new_n803_));
  AOI211_X1 g602(.A(new_n803_), .B(new_n278_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n802_), .A2(new_n804_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n766_), .A2(KEYINPUT115), .A3(KEYINPUT56), .A4(new_n279_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(new_n790_), .A3(new_n280_), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT116), .B1(new_n805_), .B2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n777_), .A2(new_n803_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n809_), .A2(new_n801_), .A3(new_n767_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n334_), .A2(new_n789_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n804_), .B2(KEYINPUT115), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n810_), .A2(new_n812_), .A3(new_n813_), .A4(new_n280_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT58), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n808_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n621_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT117), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n810_), .A2(new_n812_), .A3(KEYINPUT58), .A4(new_n280_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n816_), .A2(new_n621_), .A3(KEYINPUT117), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n819_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n798_), .A2(KEYINPUT57), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n800_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n800_), .A2(new_n822_), .A3(KEYINPUT118), .A4(new_n823_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n586_), .A3(new_n827_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n660_), .A2(new_n628_), .A3(new_n288_), .A4(new_n724_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n829_), .B(KEYINPUT54), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  NOR4_X1   g630(.A1(new_n639_), .A2(new_n490_), .A3(new_n562_), .A4(new_n470_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n761_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n831_), .A2(new_n761_), .A3(new_n832_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(G113gat), .B1(new_n836_), .B2(new_n338_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n831_), .A2(new_n832_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT59), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n793_), .A2(new_n794_), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n822_), .A2(new_n823_), .A3(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n830_), .B1(new_n841_), .B2(new_n724_), .ZN(new_n842_));
  XOR2_X1   g641(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n832_), .A3(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n839_), .A2(new_n844_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n845_), .A2(new_n410_), .A3(new_n628_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n837_), .A2(new_n846_), .ZN(G1340gat));
  OAI21_X1  g646(.A(new_n418_), .B1(new_n288_), .B2(KEYINPUT60), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n836_), .B(new_n848_), .C1(KEYINPUT60), .C2(new_n418_), .ZN(new_n849_));
  OAI21_X1  g648(.A(G120gat), .B1(new_n845_), .B2(new_n290_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1341gat));
  INV_X1    g650(.A(new_n835_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n724_), .B1(new_n852_), .B2(new_n833_), .ZN(new_n853_));
  INV_X1    g652(.A(G127gat), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(KEYINPUT121), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT121), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n853_), .A2(new_n857_), .A3(new_n854_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n845_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n586_), .A2(new_n854_), .ZN(new_n860_));
  AOI22_X1  g659(.A1(new_n856_), .A2(new_n858_), .B1(new_n859_), .B2(new_n860_), .ZN(G1342gat));
  AND3_X1   g660(.A1(new_n859_), .A2(G134gat), .A3(new_n621_), .ZN(new_n862_));
  AOI21_X1  g661(.A(G134gat), .B1(new_n836_), .B2(new_n797_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(G1343gat));
  AOI21_X1  g663(.A(new_n648_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n865_), .A2(new_n491_), .A3(new_n562_), .A4(new_n634_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n628_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT122), .B(G141gat), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(G1344gat));
  NOR2_X1   g668(.A1(new_n866_), .A2(new_n290_), .ZN(new_n870_));
  XOR2_X1   g669(.A(new_n870_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g670(.A1(new_n866_), .A2(new_n586_), .ZN(new_n872_));
  XOR2_X1   g671(.A(KEYINPUT61), .B(G155gat), .Z(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1346gat));
  NOR3_X1   g673(.A1(new_n866_), .A2(new_n590_), .A3(new_n660_), .ZN(new_n875_));
  OR2_X1    g674(.A1(new_n866_), .A2(new_n630_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n590_), .B2(new_n876_), .ZN(G1347gat));
  NAND2_X1  g676(.A1(new_n639_), .A2(new_n492_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n842_), .A2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n403_), .ZN(new_n881_));
  OAI21_X1  g680(.A(G169gat), .B1(new_n881_), .B2(new_n628_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT62), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n881_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n885_), .A2(new_n338_), .A3(new_n435_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n882_), .A2(new_n883_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n884_), .A2(new_n886_), .A3(new_n887_), .ZN(G1348gat));
  OAI21_X1  g687(.A(new_n434_), .B1(new_n881_), .B2(new_n288_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n562_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n890_), .A2(G176gat), .A3(new_n289_), .A4(new_n879_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n889_), .A2(new_n891_), .ZN(G1349gat));
  NOR3_X1   g691(.A1(new_n881_), .A2(new_n448_), .A3(new_n586_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(KEYINPUT123), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n878_), .A2(new_n586_), .ZN(new_n895_));
  AOI21_X1  g694(.A(G183gat), .B1(new_n890_), .B2(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n894_), .A2(new_n896_), .ZN(G1350gat));
  OAI21_X1  g696(.A(G190gat), .B1(new_n881_), .B2(new_n660_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n797_), .A2(new_n495_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n881_), .B2(new_n899_), .ZN(G1351gat));
  NOR2_X1   g699(.A1(new_n403_), .A2(new_n491_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n634_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n865_), .A2(G197gat), .A3(new_n338_), .A4(new_n903_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n904_), .A2(KEYINPUT124), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n904_), .A2(KEYINPUT124), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n831_), .A2(new_n338_), .A3(new_n470_), .A4(new_n903_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT125), .ZN(new_n908_));
  INV_X1    g707(.A(G197gat), .ZN(new_n909_));
  AND3_X1   g708(.A1(new_n907_), .A2(new_n908_), .A3(new_n909_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n908_), .B1(new_n907_), .B2(new_n909_), .ZN(new_n911_));
  OAI22_X1  g710(.A1(new_n905_), .A2(new_n906_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT126), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n904_), .A2(KEYINPUT124), .ZN(new_n915_));
  INV_X1    g714(.A(new_n903_), .ZN(new_n916_));
  AOI211_X1 g715(.A(new_n648_), .B(new_n916_), .C1(new_n828_), .C2(new_n830_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n917_), .A2(new_n918_), .A3(G197gat), .A4(new_n338_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n915_), .A2(new_n919_), .ZN(new_n920_));
  OAI211_X1 g719(.A(new_n920_), .B(KEYINPUT126), .C1(new_n911_), .C2(new_n910_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n914_), .A2(new_n921_), .ZN(G1352gat));
  NAND2_X1  g721(.A1(new_n917_), .A2(new_n289_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g723(.A1(new_n865_), .A2(new_n903_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n925_), .A2(new_n586_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT63), .ZN(new_n927_));
  INV_X1    g726(.A(G211gat), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n927_), .A2(new_n928_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n930_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n926_), .A2(new_n929_), .A3(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(KEYINPUT127), .ZN(new_n933_));
  OR2_X1    g732(.A1(new_n926_), .A2(new_n929_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT127), .ZN(new_n935_));
  NAND4_X1  g734(.A1(new_n926_), .A2(new_n935_), .A3(new_n929_), .A4(new_n931_), .ZN(new_n936_));
  AND3_X1   g735(.A1(new_n933_), .A2(new_n934_), .A3(new_n936_), .ZN(G1354gat));
  AND3_X1   g736(.A1(new_n917_), .A2(G218gat), .A3(new_n621_), .ZN(new_n938_));
  AOI21_X1  g737(.A(G218gat), .B1(new_n917_), .B2(new_n797_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1355gat));
endmodule


