//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 1 0 0 0 0 0 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 0 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n819_,
    new_n820_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n835_, new_n836_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G113gat), .B(G120gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n204_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(new_n202_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  XOR2_X1   g007(.A(new_n208_), .B(KEYINPUT31), .Z(new_n209_));
  INV_X1    g008(.A(KEYINPUT83), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(G183gat), .A3(G190gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  AND3_X1   g012(.A1(new_n213_), .A2(KEYINPUT80), .A3(KEYINPUT23), .ZN(new_n214_));
  AOI21_X1  g013(.A(KEYINPUT80), .B1(new_n213_), .B2(KEYINPUT23), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n212_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  OR2_X1    g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT22), .B(G169gat), .ZN(new_n221_));
  INV_X1    g020(.A(G176gat), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n220_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n218_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT25), .B(G183gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT26), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT78), .B1(new_n226_), .B2(G190gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT26), .B(G190gat), .ZN(new_n228_));
  OAI211_X1 g027(.A(new_n225_), .B(new_n227_), .C1(new_n228_), .C2(KEYINPUT78), .ZN(new_n229_));
  NOR3_X1   g028(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n213_), .A2(KEYINPUT23), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n230_), .B1(new_n212_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(G169gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(new_n222_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n234_), .A2(KEYINPUT24), .A3(new_n219_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT79), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT24), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n238_), .B1(G169gat), .B2(G176gat), .ZN(new_n239_));
  AOI21_X1  g038(.A(KEYINPUT79), .B1(new_n239_), .B2(new_n234_), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n229_), .B(new_n232_), .C1(new_n237_), .C2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n224_), .A2(new_n241_), .ZN(new_n242_));
  XOR2_X1   g041(.A(new_n242_), .B(KEYINPUT30), .Z(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT82), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n242_), .B(KEYINPUT30), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT82), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G227gat), .A2(G233gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT81), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(G71gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G15gat), .B(G43gat), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n251_), .B(G99gat), .Z(new_n252_));
  XNOR2_X1  g051(.A(new_n250_), .B(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n244_), .A2(new_n247_), .A3(new_n253_), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n247_), .A2(new_n253_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n210_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n209_), .B1(new_n256_), .B2(KEYINPUT84), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT83), .B1(new_n209_), .B2(KEYINPUT84), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n254_), .A2(new_n255_), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(G141gat), .A2(G148gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT3), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n261_), .A2(KEYINPUT85), .A3(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT85), .ZN(new_n264_));
  OAI22_X1  g063(.A1(new_n264_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G141gat), .A2(G148gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT2), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n263_), .A2(new_n265_), .A3(new_n268_), .A4(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(G155gat), .B(G162gat), .Z(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(G155gat), .ZN(new_n273_));
  INV_X1    g072(.A(G162gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT1), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT1), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n276_), .A2(G155gat), .A3(G162gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n273_), .A2(new_n274_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n275_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(G141gat), .B(G148gat), .Z(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n272_), .A2(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n282_), .A2(KEYINPUT29), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT88), .ZN(new_n284_));
  INV_X1    g083(.A(G211gat), .ZN(new_n285_));
  INV_X1    g084(.A(G218gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(G204gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(G197gat), .ZN(new_n289_));
  INV_X1    g088(.A(G197gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(G204gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G211gat), .A2(G218gat), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n287_), .A2(new_n289_), .A3(new_n291_), .A4(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT87), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n289_), .A2(new_n291_), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n287_), .A2(new_n292_), .ZN(new_n296_));
  AOI22_X1  g095(.A1(new_n293_), .A2(KEYINPUT21), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  AND3_X1   g096(.A1(new_n295_), .A2(KEYINPUT21), .A3(new_n296_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n284_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n295_), .A2(KEYINPUT21), .A3(new_n296_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT21), .ZN(new_n301_));
  XOR2_X1   g100(.A(G211gat), .B(G218gat), .Z(new_n302_));
  XNOR2_X1  g101(.A(G197gat), .B(G204gat), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n301_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  AOI22_X1  g103(.A1(new_n303_), .A2(new_n294_), .B1(new_n287_), .B2(new_n292_), .ZN(new_n305_));
  OAI211_X1 g104(.A(KEYINPUT88), .B(new_n300_), .C1(new_n304_), .C2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n299_), .A2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n282_), .A2(KEYINPUT86), .A3(KEYINPUT29), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G228gat), .A2(G233gat), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT86), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n270_), .A2(new_n271_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT29), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n310_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .A4(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n297_), .A2(new_n298_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n315_), .B1(new_n312_), .B2(new_n311_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n316_), .A2(G228gat), .A3(G233gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G78gat), .B(G106gat), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n314_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n318_), .B1(new_n314_), .B2(new_n317_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n283_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n314_), .A2(new_n317_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n318_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n283_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n314_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n324_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G22gat), .B(G50gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT28), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT89), .B(KEYINPUT90), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  AND3_X1   g130(.A1(new_n321_), .A2(new_n327_), .A3(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n331_), .B1(new_n321_), .B2(new_n327_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT20), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n231_), .A2(new_n212_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n217_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n223_), .A2(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n230_), .B1(new_n239_), .B2(new_n234_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n216_), .A2(new_n340_), .ZN(new_n341_));
  XOR2_X1   g140(.A(KEYINPUT26), .B(G190gat), .Z(new_n342_));
  NOR2_X1   g141(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n344_), .A2(KEYINPUT92), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT92), .ZN(new_n347_));
  INV_X1    g146(.A(new_n345_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n347_), .B1(new_n348_), .B2(new_n343_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n342_), .B1(new_n346_), .B2(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n339_), .B1(new_n341_), .B2(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n336_), .B1(new_n351_), .B2(new_n315_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n352_), .B1(new_n307_), .B2(new_n242_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G226gat), .A2(G233gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT19), .ZN(new_n355_));
  XOR2_X1   g154(.A(new_n355_), .B(KEYINPUT91), .Z(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n353_), .A2(new_n357_), .ZN(new_n358_));
  XOR2_X1   g157(.A(G8gat), .B(G36gat), .Z(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(G92gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT18), .B(G64gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT32), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n307_), .A2(new_n242_), .A3(KEYINPUT93), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(KEYINPUT93), .B1(new_n307_), .B2(new_n242_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT94), .B1(new_n351_), .B2(new_n315_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n225_), .A2(new_n347_), .ZN(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT92), .B1(new_n344_), .B2(new_n345_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n228_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n371_), .A2(new_n216_), .A3(new_n340_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT94), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n300_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n372_), .A2(new_n373_), .A3(new_n374_), .A4(new_n339_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n355_), .A2(new_n336_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n368_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n358_), .B(new_n363_), .C1(new_n367_), .C2(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n353_), .A2(new_n357_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n372_), .A2(new_n374_), .A3(new_n339_), .ZN(new_n380_));
  OAI211_X1 g179(.A(KEYINPUT20), .B(new_n380_), .C1(new_n365_), .C2(new_n366_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n379_), .B1(new_n381_), .B2(new_n355_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n378_), .B1(new_n382_), .B2(new_n363_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G225gat), .A2(G233gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n282_), .A2(new_n208_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n311_), .A2(new_n205_), .A3(new_n207_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n386_), .A3(KEYINPUT4), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT4), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n282_), .A2(new_n388_), .A3(new_n208_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n384_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n390_));
  AOI22_X1  g189(.A1(new_n385_), .A2(new_n386_), .B1(G225gat), .B2(G233gat), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G1gat), .B(G29gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(G85gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT0), .B(G57gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(KEYINPUT99), .B1(new_n392_), .B2(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n392_), .A2(new_n396_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT99), .ZN(new_n399_));
  INV_X1    g198(.A(new_n396_), .ZN(new_n400_));
  NOR4_X1   g199(.A1(new_n390_), .A2(new_n399_), .A3(new_n400_), .A4(new_n391_), .ZN(new_n401_));
  NOR3_X1   g200(.A1(new_n397_), .A2(new_n398_), .A3(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n383_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n362_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n366_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n377_), .B1(new_n405_), .B2(new_n364_), .ZN(new_n406_));
  OR2_X1    g205(.A1(new_n307_), .A2(new_n242_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n356_), .B1(new_n407_), .B2(new_n352_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n404_), .B1(new_n406_), .B2(new_n408_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n362_), .B(new_n358_), .C1(new_n367_), .C2(new_n377_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(KEYINPUT95), .A3(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n406_), .A2(new_n408_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT95), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n412_), .A2(new_n413_), .A3(new_n362_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n411_), .A2(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(KEYINPUT96), .A2(KEYINPUT33), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n416_), .B1(new_n392_), .B2(new_n396_), .ZN(new_n417_));
  OAI221_X1 g216(.A(new_n400_), .B1(KEYINPUT96), .B2(KEYINPUT33), .C1(new_n390_), .C2(new_n391_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n385_), .A2(new_n386_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n384_), .B1(new_n419_), .B2(KEYINPUT97), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n420_), .B1(KEYINPUT97), .B2(new_n419_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n387_), .A2(new_n384_), .A3(new_n389_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(new_n422_), .A3(new_n396_), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n417_), .A2(new_n418_), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n415_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT98), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n403_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n415_), .A2(KEYINPUT98), .A3(new_n424_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n335_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  XOR2_X1   g228(.A(KEYINPUT100), .B(KEYINPUT27), .Z(new_n430_));
  NAND3_X1  g229(.A1(new_n411_), .A2(new_n414_), .A3(new_n430_), .ZN(new_n431_));
  OAI211_X1 g230(.A(KEYINPUT27), .B(new_n410_), .C1(new_n382_), .C2(new_n362_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n433_), .A2(new_n402_), .A3(new_n335_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n260_), .B1(new_n429_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT102), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n334_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT101), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT101), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n334_), .A2(new_n431_), .A3(new_n439_), .A4(new_n432_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n438_), .A2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n257_), .A2(new_n402_), .A3(new_n259_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n436_), .B1(new_n441_), .B2(new_n443_), .ZN(new_n444_));
  AOI211_X1 g243(.A(KEYINPUT102), .B(new_n442_), .C1(new_n438_), .C2(new_n440_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n435_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G99gat), .A2(G106gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT6), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n449_));
  OR3_X1    g248(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT8), .ZN(new_n452_));
  XOR2_X1   g251(.A(G85gat), .B(G92gat), .Z(new_n453_));
  AND3_X1   g252(.A1(new_n451_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n452_), .B1(new_n451_), .B2(new_n453_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n456_), .B1(G85gat), .B2(G92gat), .ZN(new_n457_));
  XOR2_X1   g256(.A(KEYINPUT66), .B(G92gat), .Z(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(G85gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(KEYINPUT65), .B(KEYINPUT9), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n457_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  XOR2_X1   g260(.A(KEYINPUT10), .B(G99gat), .Z(new_n462_));
  XOR2_X1   g261(.A(KEYINPUT64), .B(G106gat), .Z(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(new_n448_), .ZN(new_n465_));
  OAI22_X1  g264(.A1(new_n454_), .A2(new_n455_), .B1(new_n461_), .B2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G57gat), .B(G64gat), .ZN(new_n467_));
  OR2_X1    g266(.A1(new_n467_), .A2(KEYINPUT11), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(KEYINPUT11), .ZN(new_n469_));
  XOR2_X1   g268(.A(G71gat), .B(G78gat), .Z(new_n470_));
  NAND3_X1  g269(.A1(new_n468_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  OR2_X1    g270(.A1(new_n469_), .A2(new_n470_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n466_), .A2(KEYINPUT12), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n466_), .A2(KEYINPUT67), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT67), .ZN(new_n477_));
  OAI221_X1 g276(.A(new_n477_), .B1(new_n461_), .B2(new_n465_), .C1(new_n454_), .C2(new_n455_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n475_), .B1(new_n479_), .B2(new_n473_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G230gat), .A2(G233gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n476_), .A2(new_n478_), .A3(new_n474_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT12), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n480_), .A2(new_n481_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n482_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n479_), .A2(new_n473_), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n487_), .A2(KEYINPUT68), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(KEYINPUT68), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n486_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n485_), .B1(new_n490_), .B2(new_n481_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G120gat), .B(G148gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(new_n288_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT5), .B(G176gat), .ZN(new_n494_));
  XOR2_X1   g293(.A(new_n493_), .B(new_n494_), .Z(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n491_), .A2(new_n496_), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n485_), .B(new_n495_), .C1(new_n490_), .C2(new_n481_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT13), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n497_), .A2(KEYINPUT13), .A3(new_n498_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G15gat), .B(G22gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G1gat), .A2(G8gat), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT73), .ZN(new_n506_));
  AND3_X1   g305(.A1(new_n505_), .A2(new_n506_), .A3(KEYINPUT14), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n506_), .B1(new_n505_), .B2(KEYINPUT14), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n504_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT74), .ZN(new_n510_));
  XOR2_X1   g309(.A(G1gat), .B(G8gat), .Z(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(G43gat), .B(G50gat), .Z(new_n513_));
  XNOR2_X1  g312(.A(G29gat), .B(G36gat), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n514_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT76), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n512_), .B(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G229gat), .A2(G233gat), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n512_), .ZN(new_n523_));
  XOR2_X1   g322(.A(new_n517_), .B(KEYINPUT15), .Z(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n512_), .A2(new_n518_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n525_), .A2(new_n520_), .A3(new_n526_), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n522_), .A2(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(G169gat), .B(G197gat), .Z(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT77), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G113gat), .B(G141gat), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n530_), .B(new_n531_), .Z(new_n532_));
  NOR2_X1   g331(.A1(new_n528_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n522_), .A2(new_n527_), .A3(new_n532_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n503_), .A2(new_n536_), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n446_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n517_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n479_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n524_), .A2(new_n466_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT69), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT69), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n524_), .A2(new_n543_), .A3(new_n466_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n540_), .A2(new_n542_), .A3(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G232gat), .A2(G233gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT34), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n547_), .A2(KEYINPUT35), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n545_), .A2(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n547_), .A2(KEYINPUT35), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n540_), .A2(new_n541_), .A3(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(G190gat), .B(G218gat), .Z(new_n553_));
  XNOR2_X1  g352(.A(G134gat), .B(G162gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT36), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n557_), .B(KEYINPUT70), .Z(new_n558_));
  NAND3_X1  g357(.A1(new_n549_), .A2(new_n552_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT71), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n549_), .A2(KEYINPUT71), .A3(new_n552_), .A4(new_n558_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT37), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n549_), .A2(new_n552_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n555_), .B(KEYINPUT36), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n564_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n563_), .A2(new_n567_), .ZN(new_n568_));
  AND2_X1   g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n512_), .B(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(new_n473_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT75), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G127gat), .B(G155gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(new_n285_), .ZN(new_n574_));
  XOR2_X1   g373(.A(KEYINPUT16), .B(G183gat), .Z(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT17), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  OR3_X1    g377(.A1(new_n571_), .A2(new_n572_), .A3(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n578_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n576_), .A2(KEYINPUT17), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n571_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n579_), .A2(new_n580_), .A3(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n565_), .A2(new_n566_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT72), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT72), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n565_), .A2(new_n586_), .A3(new_n566_), .ZN(new_n587_));
  AOI22_X1  g386(.A1(new_n585_), .A2(new_n587_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n568_), .B(new_n583_), .C1(new_n588_), .C2(KEYINPUT37), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n538_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(G1gat), .ZN(new_n592_));
  INV_X1    g391(.A(new_n402_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n591_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT38), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n537_), .A2(new_n583_), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n597_), .B(KEYINPUT103), .Z(new_n598_));
  INV_X1    g397(.A(new_n587_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n586_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n563_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT104), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n446_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n598_), .A2(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(G1gat), .B1(new_n604_), .B2(new_n402_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n594_), .A2(new_n595_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n596_), .A2(new_n605_), .A3(new_n606_), .ZN(G1324gat));
  INV_X1    g406(.A(G8gat), .ZN(new_n608_));
  INV_X1    g407(.A(new_n433_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n591_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n598_), .A2(new_n609_), .A3(new_n603_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT39), .ZN(new_n612_));
  AND3_X1   g411(.A1(new_n611_), .A2(new_n612_), .A3(G8gat), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n612_), .B1(new_n611_), .B2(G8gat), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n610_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT40), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(G1325gat));
  OAI21_X1  g416(.A(G15gat), .B1(new_n604_), .B2(new_n260_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(KEYINPUT41), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT41), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n620_), .B(G15gat), .C1(new_n604_), .C2(new_n260_), .ZN(new_n621_));
  INV_X1    g420(.A(G15gat), .ZN(new_n622_));
  INV_X1    g421(.A(new_n260_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n591_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n619_), .A2(new_n621_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT105), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(G1326gat));
  OAI21_X1  g426(.A(G22gat), .B1(new_n604_), .B2(new_n334_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT42), .ZN(new_n629_));
  INV_X1    g428(.A(G22gat), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n591_), .A2(new_n630_), .A3(new_n335_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n629_), .A2(new_n631_), .ZN(G1327gat));
  NOR3_X1   g431(.A1(new_n503_), .A2(new_n583_), .A3(new_n536_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT43), .ZN(new_n634_));
  AOI22_X1  g433(.A1(new_n601_), .A2(new_n564_), .B1(new_n563_), .B2(new_n567_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n446_), .A2(new_n634_), .A3(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n634_), .B1(new_n446_), .B2(new_n636_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n633_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT44), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  OAI211_X1 g440(.A(KEYINPUT44), .B(new_n633_), .C1(new_n637_), .C2(new_n638_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G29gat), .B1(new_n643_), .B2(new_n402_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n601_), .A2(new_n583_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n538_), .A2(new_n645_), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n402_), .A2(G29gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n644_), .B1(new_n646_), .B2(new_n647_), .ZN(G1328gat));
  NOR3_X1   g447(.A1(new_n646_), .A2(G36gat), .A3(new_n433_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT45), .Z(new_n650_));
  NAND3_X1  g449(.A1(new_n641_), .A2(new_n609_), .A3(new_n642_), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n651_), .A2(KEYINPUT106), .A3(G36gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(KEYINPUT106), .B1(new_n651_), .B2(G36gat), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n650_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT46), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  OAI211_X1 g455(.A(KEYINPUT46), .B(new_n650_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1329gat));
  NOR3_X1   g457(.A1(new_n646_), .A2(G43gat), .A3(new_n260_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n641_), .A2(new_n623_), .A3(new_n642_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n660_), .B2(G43gat), .ZN(new_n661_));
  XNOR2_X1  g460(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n661_), .B(new_n662_), .Z(G1330gat));
  OAI21_X1  g462(.A(G50gat), .B1(new_n643_), .B2(new_n334_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n334_), .A2(G50gat), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n664_), .B1(new_n646_), .B2(new_n665_), .ZN(G1331gat));
  INV_X1    g465(.A(new_n503_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n536_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n603_), .A2(new_n583_), .A3(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n670_), .A2(G57gat), .A3(new_n593_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT109), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n671_), .A2(new_n672_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n590_), .A2(new_n503_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT108), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n446_), .A2(new_n536_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(G57gat), .B1(new_n678_), .B2(new_n593_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n673_), .A2(new_n674_), .A3(new_n679_), .ZN(G1332gat));
  INV_X1    g479(.A(G64gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n681_), .B1(new_n670_), .B2(new_n609_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT48), .Z(new_n683_));
  NAND3_X1  g482(.A1(new_n678_), .A2(new_n681_), .A3(new_n609_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1333gat));
  INV_X1    g484(.A(G71gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n686_), .B1(new_n670_), .B2(new_n623_), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT49), .Z(new_n688_));
  NAND3_X1  g487(.A1(new_n678_), .A2(new_n686_), .A3(new_n623_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1334gat));
  INV_X1    g489(.A(G78gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n691_), .B1(new_n670_), .B2(new_n335_), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT50), .Z(new_n693_));
  NAND3_X1  g492(.A1(new_n678_), .A2(new_n691_), .A3(new_n335_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1335gat));
  OR2_X1    g494(.A1(new_n637_), .A2(new_n638_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n583_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n696_), .A2(new_n697_), .A3(new_n669_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n699_), .A2(G85gat), .A3(new_n593_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n677_), .A2(new_n503_), .A3(new_n645_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT110), .ZN(new_n702_));
  AOI21_X1  g501(.A(G85gat), .B1(new_n702_), .B2(new_n593_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n700_), .A2(new_n703_), .ZN(G1336gat));
  AOI21_X1  g503(.A(G92gat), .B1(new_n702_), .B2(new_n609_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n609_), .A2(new_n458_), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT111), .Z(new_n707_));
  AOI21_X1  g506(.A(new_n705_), .B1(new_n699_), .B2(new_n707_), .ZN(G1337gat));
  OAI21_X1  g507(.A(G99gat), .B1(new_n698_), .B2(new_n260_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n623_), .A2(new_n462_), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n702_), .A2(KEYINPUT112), .A3(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(KEYINPUT112), .B1(new_n702_), .B2(new_n710_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n709_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT51), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT51), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n715_), .B(new_n709_), .C1(new_n711_), .C2(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1338gat));
  NAND3_X1  g516(.A1(new_n702_), .A2(new_n463_), .A3(new_n335_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n696_), .A2(new_n697_), .A3(new_n335_), .A4(new_n669_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT52), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n719_), .A2(new_n720_), .A3(G106gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n719_), .B2(G106gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n718_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT53), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT53), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n725_), .B(new_n718_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1339gat));
  NAND3_X1  g526(.A1(new_n441_), .A2(new_n593_), .A3(new_n623_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n480_), .A2(KEYINPUT55), .A3(new_n484_), .A4(new_n481_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT114), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT55), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n485_), .A2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n480_), .A2(new_n484_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(G230gat), .A3(G233gat), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n731_), .A2(new_n733_), .A3(new_n735_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n730_), .A2(KEYINPUT114), .ZN(new_n737_));
  OAI211_X1 g536(.A(KEYINPUT56), .B(new_n496_), .C1(new_n736_), .C2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(KEYINPUT115), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n496_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT56), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n730_), .A2(KEYINPUT114), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n743_), .A2(new_n731_), .A3(new_n733_), .A4(new_n735_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT115), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n744_), .A2(new_n745_), .A3(KEYINPUT56), .A4(new_n496_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n739_), .A2(new_n742_), .A3(new_n746_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n668_), .A2(new_n498_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n519_), .A2(new_n520_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n532_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n525_), .A2(new_n521_), .A3(new_n526_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n750_), .A2(new_n751_), .A3(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n534_), .A2(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n754_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n749_), .A2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(KEYINPUT57), .B1(new_n757_), .B2(new_n601_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n755_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT57), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n759_), .A2(new_n760_), .A3(new_n588_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n758_), .A2(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n740_), .A2(KEYINPUT116), .A3(new_n741_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n754_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n498_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT116), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n738_), .A2(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(KEYINPUT56), .B1(new_n744_), .B2(new_n496_), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n763_), .B(new_n766_), .C1(new_n768_), .C2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT58), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n635_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT117), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n765_), .B1(new_n769_), .B2(KEYINPUT116), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n742_), .A2(new_n767_), .A3(new_n738_), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT58), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(KEYINPUT117), .B1(new_n777_), .B2(new_n635_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n775_), .A2(new_n776_), .A3(KEYINPUT58), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n774_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n583_), .B1(new_n762_), .B2(new_n780_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n501_), .A2(new_n536_), .A3(new_n502_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT54), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n782_), .A2(new_n590_), .A3(KEYINPUT113), .A4(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n501_), .A2(new_n536_), .A3(new_n502_), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT54), .B1(new_n785_), .B2(new_n589_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n785_), .A2(new_n589_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT113), .B1(new_n788_), .B2(new_n783_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n729_), .B1(new_n781_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(G113gat), .B1(new_n792_), .B2(new_n668_), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT118), .B1(new_n791_), .B2(KEYINPUT59), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n757_), .A2(KEYINPUT57), .A3(new_n601_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n760_), .B1(new_n759_), .B2(new_n588_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n779_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n777_), .A2(KEYINPUT117), .A3(new_n635_), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n796_), .B(new_n797_), .C1(new_n798_), .C2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n790_), .B1(new_n800_), .B2(new_n697_), .ZN(new_n801_));
  OAI211_X1 g600(.A(KEYINPUT118), .B(KEYINPUT59), .C1(new_n801_), .C2(new_n728_), .ZN(new_n802_));
  OAI22_X1  g601(.A1(new_n781_), .A2(KEYINPUT119), .B1(new_n789_), .B2(new_n787_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n800_), .A2(KEYINPUT119), .A3(new_n697_), .ZN(new_n804_));
  OR2_X1    g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n728_), .A2(KEYINPUT59), .ZN(new_n806_));
  AOI22_X1  g605(.A1(new_n795_), .A2(new_n802_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n668_), .A2(G113gat), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT120), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n793_), .B1(new_n807_), .B2(new_n809_), .ZN(G1340gat));
  OAI21_X1  g609(.A(new_n806_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n802_), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n503_), .B(new_n811_), .C1(new_n812_), .C2(new_n794_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(G120gat), .ZN(new_n814_));
  INV_X1    g613(.A(G120gat), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(new_n667_), .B2(KEYINPUT60), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n792_), .B(new_n816_), .C1(KEYINPUT60), .C2(new_n815_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n814_), .A2(new_n817_), .ZN(G1341gat));
  AOI21_X1  g617(.A(G127gat), .B1(new_n792_), .B2(new_n583_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n583_), .A2(G127gat), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n807_), .B2(new_n820_), .ZN(G1342gat));
  INV_X1    g620(.A(G134gat), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n822_), .B1(new_n791_), .B2(new_n602_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT121), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  OAI211_X1 g624(.A(KEYINPUT121), .B(new_n822_), .C1(new_n791_), .C2(new_n602_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n635_), .A2(new_n822_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n827_), .B1(new_n807_), .B2(new_n828_), .ZN(G1343gat));
  NOR3_X1   g628(.A1(new_n609_), .A2(new_n623_), .A3(new_n402_), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n335_), .B(new_n830_), .C1(new_n781_), .C2(new_n790_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n831_), .A2(new_n536_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(KEYINPUT122), .B(G141gat), .ZN(new_n833_));
  XOR2_X1   g632(.A(new_n832_), .B(new_n833_), .Z(G1344gat));
  NOR2_X1   g633(.A1(new_n831_), .A2(new_n667_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT123), .B(G148gat), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n835_), .B(new_n836_), .ZN(G1345gat));
  OR3_X1    g636(.A1(new_n831_), .A2(KEYINPUT124), .A3(new_n697_), .ZN(new_n838_));
  OAI21_X1  g637(.A(KEYINPUT124), .B1(new_n831_), .B2(new_n697_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(KEYINPUT61), .B(G155gat), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n838_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n840_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(G1346gat));
  INV_X1    g642(.A(KEYINPUT126), .ZN(new_n844_));
  OAI211_X1 g643(.A(KEYINPUT125), .B(new_n274_), .C1(new_n831_), .C2(new_n602_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n801_), .A2(new_n334_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n846_), .A2(G162gat), .A3(new_n636_), .A4(new_n830_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n801_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n602_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n849_), .A2(new_n335_), .A3(new_n850_), .A4(new_n830_), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT125), .B1(new_n851_), .B2(new_n274_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n844_), .B1(new_n848_), .B2(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n274_), .B1(new_n831_), .B2(new_n602_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT125), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n856_), .A2(KEYINPUT126), .A3(new_n845_), .A4(new_n847_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n853_), .A2(new_n857_), .ZN(G1347gat));
  NOR3_X1   g657(.A1(new_n442_), .A2(new_n433_), .A3(new_n335_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n668_), .B(new_n859_), .C1(new_n803_), .C2(new_n804_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(G169gat), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT62), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n860_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n805_), .A2(new_n221_), .A3(new_n668_), .A4(new_n859_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n863_), .A2(new_n864_), .A3(new_n865_), .ZN(G1348gat));
  AND4_X1   g665(.A1(G176gat), .A2(new_n849_), .A3(new_n503_), .A4(new_n859_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n503_), .B(new_n859_), .C1(new_n803_), .C2(new_n804_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n222_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT127), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n868_), .A2(KEYINPUT127), .A3(new_n222_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n867_), .B1(new_n871_), .B2(new_n872_), .ZN(G1349gat));
  AND2_X1   g672(.A1(new_n859_), .A2(new_n583_), .ZN(new_n874_));
  AOI21_X1  g673(.A(G183gat), .B1(new_n790_), .B2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n805_), .A2(new_n859_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n697_), .A2(new_n370_), .A3(new_n369_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n875_), .B1(new_n877_), .B2(new_n878_), .ZN(G1350gat));
  OAI21_X1  g678(.A(G190gat), .B1(new_n876_), .B2(new_n635_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n805_), .A2(new_n228_), .A3(new_n850_), .A4(new_n859_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1351gat));
  NOR3_X1   g681(.A1(new_n623_), .A2(new_n433_), .A3(new_n593_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n846_), .A2(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n536_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(new_n290_), .ZN(G1352gat));
  NOR2_X1   g685(.A1(new_n884_), .A2(new_n667_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(new_n288_), .ZN(G1353gat));
  AOI21_X1  g687(.A(new_n697_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n846_), .A2(new_n883_), .A3(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1354gat));
  NOR3_X1   g691(.A1(new_n884_), .A2(new_n286_), .A3(new_n635_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n884_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n850_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n286_), .B2(new_n895_), .ZN(G1355gat));
endmodule


