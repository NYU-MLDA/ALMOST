//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 0 0 0 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n897_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n937_, new_n938_, new_n940_, new_n941_, new_n943_, new_n944_,
    new_n945_, new_n947_, new_n948_, new_n949_, new_n951_, new_n952_,
    new_n953_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT19), .ZN(new_n204_));
  OR2_X1    g003(.A1(G197gat), .A2(G204gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G197gat), .A2(G204gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT21), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n205_), .A2(KEYINPUT21), .A3(new_n206_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G211gat), .B(G218gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n210_), .A2(new_n211_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n216_), .B1(G183gat), .B2(G190gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(G183gat), .A3(G190gat), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n219_), .A2(KEYINPUT83), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(KEYINPUT83), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n218_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT25), .B(G183gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT26), .B(G190gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT82), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT82), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n223_), .A2(new_n224_), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(G169gat), .ZN(new_n229_));
  INV_X1    g028(.A(G176gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G169gat), .A2(G176gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(KEYINPUT24), .A3(new_n232_), .ZN(new_n233_));
  OR3_X1    g032(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n222_), .A2(new_n226_), .A3(new_n228_), .A4(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT22), .B1(new_n229_), .B2(KEYINPUT84), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n229_), .A2(KEYINPUT22), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n230_), .B(new_n237_), .C1(new_n238_), .C2(KEYINPUT84), .ZN(new_n239_));
  INV_X1    g038(.A(new_n219_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n240_), .A2(new_n217_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(G183gat), .A2(G190gat), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n239_), .B(new_n232_), .C1(new_n241_), .C2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n236_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT85), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT85), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n236_), .A2(new_n246_), .A3(new_n243_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n215_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n222_), .B1(G183gat), .B2(G190gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n232_), .A2(KEYINPUT94), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n232_), .A2(KEYINPUT94), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT22), .B(G169gat), .ZN(new_n252_));
  AOI22_X1  g051(.A1(new_n250_), .A2(new_n251_), .B1(new_n252_), .B2(new_n230_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n249_), .A2(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n231_), .A2(KEYINPUT24), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n241_), .A2(new_n255_), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n225_), .A2(KEYINPUT93), .A3(new_n233_), .ZN(new_n257_));
  AOI21_X1  g056(.A(KEYINPUT93), .B1(new_n225_), .B2(new_n233_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n256_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n254_), .A2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT20), .B1(new_n260_), .B2(new_n214_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n204_), .B1(new_n248_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT20), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n263_), .B1(new_n260_), .B2(new_n214_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n245_), .A2(new_n247_), .A3(new_n215_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n204_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n264_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n262_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G64gat), .B(G92gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT96), .ZN(new_n270_));
  XOR2_X1   g069(.A(KEYINPUT95), .B(KEYINPUT18), .Z(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G8gat), .B(G36gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n202_), .B1(new_n268_), .B2(new_n274_), .ZN(new_n275_));
  AND3_X1   g074(.A1(new_n236_), .A2(new_n246_), .A3(new_n243_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n246_), .B1(new_n236_), .B2(new_n243_), .ZN(new_n277_));
  NOR3_X1   g076(.A1(new_n276_), .A2(new_n277_), .A3(new_n214_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n225_), .A2(new_n233_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT93), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n225_), .A2(KEYINPUT93), .A3(new_n233_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  AOI22_X1  g082(.A1(new_n283_), .A2(new_n256_), .B1(new_n249_), .B2(new_n253_), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT20), .B1(new_n284_), .B2(new_n215_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n204_), .B1(new_n278_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n274_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n263_), .B1(new_n284_), .B2(new_n215_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n214_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(new_n289_), .A3(new_n266_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n286_), .A2(new_n287_), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT100), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT100), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n286_), .A2(new_n293_), .A3(new_n287_), .A4(new_n290_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n275_), .A2(new_n292_), .A3(new_n294_), .ZN(new_n295_));
  AND3_X1   g094(.A1(new_n288_), .A2(new_n289_), .A3(new_n266_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n266_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n274_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(new_n291_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(new_n202_), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n295_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G78gat), .B(G106gat), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT3), .ZN(new_n305_));
  INV_X1    g104(.A(G141gat), .ZN(new_n306_));
  INV_X1    g105(.A(G148gat), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G141gat), .A2(G148gat), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT2), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n308_), .A2(new_n311_), .A3(new_n312_), .A4(new_n313_), .ZN(new_n314_));
  OR2_X1    g113(.A1(G155gat), .A2(G162gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n314_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(KEYINPUT1), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT1), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n320_), .A2(G155gat), .A3(G162gat), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n319_), .A2(new_n321_), .A3(new_n315_), .ZN(new_n322_));
  XOR2_X1   g121(.A(G141gat), .B(G148gat), .Z(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n318_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT29), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT90), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n326_), .A2(new_n327_), .A3(new_n214_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n327_), .B1(new_n326_), .B2(new_n214_), .ZN(new_n330_));
  INV_X1    g129(.A(G233gat), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT89), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n332_), .A2(G228gat), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(G228gat), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n331_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NOR3_X1   g136(.A1(new_n329_), .A2(new_n330_), .A3(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n326_), .A2(new_n214_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT90), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n336_), .B1(new_n340_), .B2(new_n328_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n304_), .B1(new_n338_), .B2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT92), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  OR3_X1    g143(.A1(new_n325_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT28), .B1(new_n325_), .B2(KEYINPUT29), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G22gat), .B(G50gat), .ZN(new_n347_));
  AND3_X1   g146(.A1(new_n345_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n347_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n337_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n340_), .A2(new_n336_), .A3(new_n328_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n353_), .A2(KEYINPUT92), .A3(new_n304_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n351_), .A2(new_n303_), .A3(new_n352_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n344_), .A2(new_n350_), .A3(new_n354_), .A4(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n355_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n342_), .A2(KEYINPUT91), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT91), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n353_), .A2(new_n359_), .A3(new_n304_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n357_), .B1(new_n358_), .B2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n356_), .B1(new_n361_), .B2(new_n350_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n276_), .A2(new_n277_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G71gat), .B(G99gat), .ZN(new_n364_));
  INV_X1    g163(.A(G43gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n363_), .B(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G113gat), .B(G120gat), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G127gat), .B(G134gat), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n371_), .A2(KEYINPUT87), .ZN(new_n372_));
  INV_X1    g171(.A(G134gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(G127gat), .ZN(new_n374_));
  INV_X1    g173(.A(G127gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(G134gat), .ZN(new_n376_));
  AND3_X1   g175(.A1(new_n374_), .A2(new_n376_), .A3(KEYINPUT87), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n370_), .B1(new_n372_), .B2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n374_), .A2(new_n376_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT87), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n371_), .A2(KEYINPUT87), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n381_), .A2(new_n382_), .A3(new_n369_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n378_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT31), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(KEYINPUT86), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G227gat), .A2(G233gat), .ZN(new_n388_));
  INV_X1    g187(.A(G15gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT30), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n387_), .B(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n368_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n391_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n387_), .B(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n367_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n393_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G225gat), .A2(G233gat), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n384_), .A2(new_n325_), .ZN(new_n401_));
  AOI22_X1  g200(.A1(new_n314_), .A2(new_n317_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n378_), .A2(new_n402_), .A3(new_n383_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n401_), .A2(KEYINPUT4), .A3(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n402_), .B1(new_n383_), .B2(new_n378_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT4), .ZN(new_n406_));
  AOI21_X1  g205(.A(KEYINPUT97), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  AND4_X1   g206(.A1(KEYINPUT97), .A2(new_n384_), .A3(new_n406_), .A4(new_n325_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n400_), .B(new_n404_), .C1(new_n407_), .C2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n401_), .A2(new_n403_), .A3(new_n399_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G1gat), .B(G29gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT98), .B(G85gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT0), .B(G57gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n411_), .A2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n409_), .A2(new_n410_), .A3(new_n416_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NOR4_X1   g219(.A1(new_n302_), .A2(new_n362_), .A3(new_n398_), .A4(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n359_), .B1(new_n353_), .B2(new_n304_), .ZN(new_n422_));
  AOI211_X1 g221(.A(KEYINPUT91), .B(new_n303_), .C1(new_n351_), .C2(new_n352_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n355_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n350_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n420_), .B1(new_n426_), .B2(new_n356_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n268_), .A2(KEYINPUT32), .A3(new_n287_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n287_), .A2(KEYINPUT32), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n429_), .A2(new_n286_), .A3(new_n290_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n420_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT33), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n419_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT99), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT99), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n419_), .A2(new_n435_), .A3(new_n432_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n409_), .A2(KEYINPUT33), .A3(new_n410_), .A4(new_n416_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n399_), .B(new_n404_), .C1(new_n407_), .C2(new_n408_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n401_), .A2(new_n403_), .A3(new_n400_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n417_), .A3(new_n440_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n298_), .A2(new_n291_), .A3(new_n438_), .A4(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n431_), .B1(new_n437_), .B2(new_n442_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n354_), .A2(new_n350_), .A3(new_n355_), .ZN(new_n444_));
  AOI22_X1  g243(.A1(new_n425_), .A2(new_n424_), .B1(new_n444_), .B2(new_n344_), .ZN(new_n445_));
  AOI22_X1  g244(.A1(new_n301_), .A2(new_n427_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n393_), .A2(new_n396_), .A3(KEYINPUT88), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT88), .B1(new_n393_), .B2(new_n396_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT101), .B1(new_n446_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n443_), .A2(new_n445_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n420_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n362_), .A2(new_n300_), .A3(new_n295_), .A4(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT101), .ZN(new_n455_));
  INV_X1    g254(.A(new_n449_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n454_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n421_), .B1(new_n450_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT81), .ZN(new_n459_));
  AND2_X1   g258(.A1(G15gat), .A2(G22gat), .ZN(new_n460_));
  NOR2_X1   g259(.A1(G15gat), .A2(G22gat), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G1gat), .A2(G8gat), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n463_), .A2(KEYINPUT14), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT78), .B1(new_n462_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(KEYINPUT14), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT78), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n466_), .B(new_n467_), .C1(new_n461_), .C2(new_n460_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n465_), .A2(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(G1gat), .B(G8gat), .Z(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(G29gat), .B(G36gat), .Z(new_n473_));
  XOR2_X1   g272(.A(G43gat), .B(G50gat), .Z(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n465_), .A2(new_n470_), .A3(new_n468_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n472_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n475_), .B1(new_n472_), .B2(new_n476_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n459_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n475_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n476_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n470_), .B1(new_n465_), .B2(new_n468_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n481_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n484_), .A2(KEYINPUT81), .A3(new_n477_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n480_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G229gat), .A2(G233gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n475_), .B(KEYINPUT15), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n489_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n478_), .A2(new_n488_), .ZN(new_n491_));
  AOI22_X1  g290(.A1(new_n486_), .A2(new_n488_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G113gat), .B(G141gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G169gat), .B(G197gat), .ZN(new_n494_));
  XOR2_X1   g293(.A(new_n493_), .B(new_n494_), .Z(new_n495_));
  XNOR2_X1  g294(.A(new_n492_), .B(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G232gat), .A2(G233gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT34), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n499_), .A2(KEYINPUT35), .ZN(new_n500_));
  OR2_X1    g299(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT64), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT64), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n501_), .A2(new_n505_), .A3(new_n502_), .ZN(new_n506_));
  AOI21_X1  g305(.A(G106gat), .B1(new_n504_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G99gat), .A2(G106gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT6), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT6), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n510_), .A2(G99gat), .A3(G106gat), .ZN(new_n511_));
  AND3_X1   g310(.A1(new_n509_), .A2(new_n511_), .A3(KEYINPUT66), .ZN(new_n512_));
  AOI21_X1  g311(.A(KEYINPUT66), .B1(new_n509_), .B2(new_n511_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(G85gat), .ZN(new_n515_));
  INV_X1    g314(.A(G92gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G85gat), .A2(G92gat), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(KEYINPUT65), .A3(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(KEYINPUT9), .B1(new_n515_), .B2(new_n516_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n517_), .A2(KEYINPUT65), .A3(KEYINPUT9), .A4(new_n518_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NOR3_X1   g322(.A1(new_n507_), .A2(new_n514_), .A3(new_n523_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(G99gat), .A2(G106gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT7), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n526_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT67), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n526_), .B(KEYINPUT67), .C1(new_n512_), .C2(new_n513_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n517_), .A2(new_n518_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(KEYINPUT68), .B(KEYINPUT8), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n529_), .A2(new_n530_), .A3(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n509_), .A2(new_n511_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT69), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT69), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n509_), .A2(new_n511_), .A3(new_n537_), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n536_), .A2(new_n526_), .A3(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT8), .B1(new_n539_), .B2(new_n531_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n524_), .B1(new_n534_), .B2(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n500_), .B1(new_n541_), .B2(new_n475_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n499_), .A2(KEYINPUT35), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT15), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n475_), .B(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n541_), .A2(new_n546_), .ZN(new_n547_));
  NOR3_X1   g346(.A1(new_n543_), .A2(new_n544_), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  XOR2_X1   g348(.A(G190gat), .B(G218gat), .Z(new_n550_));
  XNOR2_X1  g349(.A(G134gat), .B(G162gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT36), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n554_), .B(KEYINPUT76), .Z(new_n555_));
  INV_X1    g354(.A(KEYINPUT74), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n556_), .B1(new_n541_), .B2(new_n546_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n533_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n558_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n536_), .A2(new_n526_), .A3(new_n538_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n560_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n561_));
  AOI22_X1  g360(.A1(new_n559_), .A2(new_n530_), .B1(new_n561_), .B2(KEYINPUT8), .ZN(new_n562_));
  OAI211_X1 g361(.A(KEYINPUT74), .B(new_n489_), .C1(new_n562_), .C2(new_n524_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n557_), .A2(new_n542_), .A3(new_n563_), .ZN(new_n564_));
  AND3_X1   g363(.A1(new_n564_), .A2(KEYINPUT75), .A3(new_n544_), .ZN(new_n565_));
  AOI21_X1  g364(.A(KEYINPUT75), .B1(new_n564_), .B2(new_n544_), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n549_), .B(new_n555_), .C1(new_n565_), .C2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n564_), .A2(new_n544_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT75), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n564_), .A2(KEYINPUT75), .A3(new_n544_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n548_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n552_), .B(new_n553_), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n573_), .B(KEYINPUT77), .Z(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n567_), .B1(new_n572_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT37), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT37), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n567_), .B(new_n578_), .C1(new_n572_), .C2(new_n573_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT70), .B(KEYINPUT12), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G57gat), .B(G64gat), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n582_), .A2(KEYINPUT11), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(KEYINPUT11), .ZN(new_n584_));
  XOR2_X1   g383(.A(G71gat), .B(G78gat), .Z(new_n585_));
  NAND3_X1  g384(.A1(new_n583_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n584_), .A2(new_n585_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n581_), .B1(new_n541_), .B2(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(G230gat), .A2(G233gat), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n590_), .B1(new_n541_), .B2(new_n588_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n588_), .ZN(new_n592_));
  OAI211_X1 g391(.A(KEYINPUT12), .B(new_n592_), .C1(new_n562_), .C2(new_n524_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n589_), .A2(new_n591_), .A3(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT71), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n541_), .A2(new_n588_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n541_), .A2(new_n588_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n590_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT71), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n589_), .A2(new_n591_), .A3(new_n600_), .A4(new_n593_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n595_), .A2(new_n599_), .A3(new_n601_), .ZN(new_n602_));
  XOR2_X1   g401(.A(G120gat), .B(G148gat), .Z(new_n603_));
  XNOR2_X1  g402(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G176gat), .B(G204gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n607_), .B(KEYINPUT73), .Z(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n602_), .A2(new_n609_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n595_), .A2(new_n599_), .A3(new_n601_), .A4(new_n607_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT13), .ZN(new_n613_));
  NAND2_X1  g412(.A1(G231gat), .A2(G233gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n588_), .B(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n482_), .A2(new_n483_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n615_), .B(new_n616_), .Z(new_n617_));
  XOR2_X1   g416(.A(G127gat), .B(G155gat), .Z(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(G183gat), .B(G211gat), .Z(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  OAI21_X1  g421(.A(KEYINPUT17), .B1(new_n617_), .B2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT80), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n622_), .B1(new_n617_), .B2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  OAI211_X1 g425(.A(KEYINPUT17), .B(new_n622_), .C1(new_n617_), .C2(new_n624_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n580_), .A2(new_n613_), .A3(new_n628_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n458_), .A2(new_n497_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(G1gat), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n630_), .A2(new_n631_), .A3(new_n420_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT38), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT102), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n567_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n458_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n613_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n628_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n639_), .A2(new_n497_), .A3(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n638_), .A2(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G1gat), .B1(new_n642_), .B2(new_n452_), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n635_), .B(new_n643_), .C1(new_n633_), .C2(new_n632_), .ZN(G1324gat));
  INV_X1    g443(.A(G8gat), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n630_), .A2(new_n645_), .A3(new_n302_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n642_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(new_n302_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT39), .ZN(new_n649_));
  AND4_X1   g448(.A1(KEYINPUT103), .A2(new_n648_), .A3(new_n649_), .A4(G8gat), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n645_), .B1(new_n651_), .B2(KEYINPUT39), .ZN(new_n652_));
  AOI22_X1  g451(.A1(new_n648_), .A2(new_n652_), .B1(KEYINPUT103), .B2(new_n649_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n646_), .B1(new_n650_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT40), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(new_n655_), .ZN(G1325gat));
  OAI21_X1  g455(.A(G15gat), .B1(new_n642_), .B2(new_n456_), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n657_), .B(KEYINPUT41), .Z(new_n658_));
  NAND3_X1  g457(.A1(new_n630_), .A2(new_n389_), .A3(new_n449_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1326gat));
  OAI21_X1  g459(.A(G22gat), .B1(new_n642_), .B2(new_n445_), .ZN(new_n661_));
  XOR2_X1   g460(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(G22gat), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n630_), .A2(new_n664_), .A3(new_n362_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n665_), .ZN(G1327gat));
  NAND2_X1  g465(.A1(new_n637_), .A2(new_n640_), .ZN(new_n667_));
  NOR4_X1   g466(.A1(new_n458_), .A2(new_n497_), .A3(new_n639_), .A4(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(G29gat), .B1(new_n668_), .B2(new_n420_), .ZN(new_n669_));
  OAI21_X1  g468(.A(KEYINPUT43), .B1(new_n458_), .B2(new_n580_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n302_), .A2(new_n362_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n671_), .A2(new_n397_), .A3(new_n452_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n455_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n673_));
  AOI211_X1 g472(.A(KEYINPUT101), .B(new_n449_), .C1(new_n451_), .C2(new_n453_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n672_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n577_), .A2(new_n579_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n675_), .A2(new_n676_), .A3(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n670_), .A2(new_n678_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n639_), .A2(new_n497_), .A3(new_n628_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n681_), .B1(KEYINPUT105), .B2(KEYINPUT44), .ZN(new_n682_));
  NOR2_X1   g481(.A1(KEYINPUT105), .A2(KEYINPUT44), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n679_), .A2(new_n683_), .A3(new_n680_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n420_), .A2(G29gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n669_), .B1(new_n685_), .B2(new_n686_), .ZN(G1328gat));
  INV_X1    g486(.A(G36gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n668_), .A2(new_n688_), .A3(new_n302_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT45), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n301_), .B1(new_n682_), .B2(new_n684_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n690_), .B1(new_n691_), .B2(new_n688_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT46), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  OAI211_X1 g493(.A(new_n690_), .B(KEYINPUT46), .C1(new_n691_), .C2(new_n688_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1329gat));
  NAND3_X1  g495(.A1(new_n668_), .A2(new_n365_), .A3(new_n449_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n398_), .B1(new_n682_), .B2(new_n684_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n697_), .B1(new_n698_), .B2(new_n365_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT47), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  OAI211_X1 g500(.A(KEYINPUT47), .B(new_n697_), .C1(new_n698_), .C2(new_n365_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1330gat));
  AOI21_X1  g502(.A(G50gat), .B1(new_n668_), .B2(new_n362_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n362_), .A2(G50gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n685_), .B2(new_n705_), .ZN(G1331gat));
  NAND4_X1  g505(.A1(new_n638_), .A2(new_n497_), .A3(new_n628_), .A4(new_n639_), .ZN(new_n707_));
  INV_X1    g506(.A(G57gat), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n707_), .A2(new_n708_), .A3(new_n452_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n677_), .A2(new_n640_), .A3(new_n613_), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n710_), .A2(KEYINPUT106), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n458_), .A2(new_n496_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(KEYINPUT106), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n711_), .A2(new_n712_), .A3(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n715_), .A2(KEYINPUT107), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(KEYINPUT107), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n716_), .A2(new_n420_), .A3(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n709_), .B1(new_n718_), .B2(new_n708_), .ZN(G1332gat));
  OAI21_X1  g518(.A(G64gat), .B1(new_n707_), .B2(new_n301_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT48), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n301_), .A2(G64gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n714_), .B2(new_n722_), .ZN(G1333gat));
  OAI21_X1  g522(.A(G71gat), .B1(new_n707_), .B2(new_n456_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT49), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n456_), .A2(G71gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n714_), .B2(new_n726_), .ZN(G1334gat));
  OAI21_X1  g526(.A(G78gat), .B1(new_n707_), .B2(new_n445_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT50), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n445_), .A2(G78gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(new_n714_), .B2(new_n730_), .ZN(G1335gat));
  NOR2_X1   g530(.A1(new_n613_), .A2(new_n667_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n712_), .A2(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(G85gat), .B1(new_n733_), .B2(new_n420_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT108), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n639_), .A2(new_n497_), .A3(new_n640_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n736_), .B1(new_n670_), .B2(new_n678_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n738_), .A2(new_n515_), .A3(new_n452_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n735_), .A2(new_n739_), .ZN(G1336gat));
  OAI21_X1  g539(.A(G92gat), .B1(new_n738_), .B2(new_n301_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n733_), .A2(new_n516_), .A3(new_n302_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1337gat));
  OAI21_X1  g542(.A(G99gat), .B1(new_n738_), .B2(new_n456_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n733_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n504_), .A2(new_n506_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n397_), .A2(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n744_), .B1(new_n745_), .B2(new_n747_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g548(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n751_));
  INV_X1    g550(.A(new_n736_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n679_), .A2(new_n751_), .A3(new_n362_), .A4(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(G106gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n751_), .B1(new_n737_), .B2(new_n362_), .ZN(new_n755_));
  OAI21_X1  g554(.A(KEYINPUT52), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n679_), .A2(new_n362_), .A3(new_n752_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT109), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n758_), .A2(new_n759_), .A3(G106gat), .A4(new_n753_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n756_), .A2(new_n760_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n745_), .A2(G106gat), .A3(new_n445_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n750_), .B1(new_n761_), .B2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n750_), .ZN(new_n765_));
  AOI211_X1 g564(.A(new_n762_), .B(new_n765_), .C1(new_n756_), .C2(new_n760_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1339gat));
  INV_X1    g566(.A(new_n629_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT54), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n769_), .A2(KEYINPUT111), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n768_), .A2(new_n497_), .A3(new_n771_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n769_), .A2(KEYINPUT111), .ZN(new_n773_));
  OAI22_X1  g572(.A1(new_n629_), .A2(new_n496_), .B1(new_n773_), .B2(new_n770_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n772_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n595_), .A2(new_n776_), .A3(new_n601_), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n589_), .A2(new_n591_), .A3(new_n593_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n589_), .A2(new_n596_), .A3(new_n593_), .ZN(new_n779_));
  AOI22_X1  g578(.A1(new_n778_), .A2(KEYINPUT55), .B1(new_n590_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n777_), .A2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n609_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT56), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n781_), .A2(KEYINPUT56), .A3(new_n609_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n485_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT81), .B1(new_n484_), .B2(new_n477_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n487_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n495_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(KEYINPUT112), .A3(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n488_), .B1(new_n480_), .B2(new_n485_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n792_), .B1(new_n793_), .B2(new_n495_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n490_), .A2(new_n477_), .A3(new_n488_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n791_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n492_), .A2(new_n495_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n798_), .A2(new_n611_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT58), .B1(new_n786_), .B2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT115), .B1(new_n800_), .B2(new_n580_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n786_), .A2(KEYINPUT58), .A3(new_n799_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT56), .B1(new_n781_), .B2(new_n609_), .ZN(new_n803_));
  AOI211_X1 g602(.A(new_n783_), .B(new_n608_), .C1(new_n777_), .C2(new_n780_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n799_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT58), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n677_), .A3(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n801_), .A2(new_n802_), .A3(new_n809_), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n612_), .A2(KEYINPUT113), .A3(new_n798_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT113), .B1(new_n612_), .B2(new_n798_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n496_), .A2(new_n611_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n637_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(KEYINPUT114), .B1(new_n816_), .B2(KEYINPUT57), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(KEYINPUT57), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n612_), .A2(KEYINPUT113), .A3(new_n798_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n612_), .A2(new_n798_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n815_), .A2(new_n819_), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n636_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT114), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n824_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n810_), .A2(new_n817_), .A3(new_n818_), .A4(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n775_), .B1(new_n828_), .B2(new_n640_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n671_), .A2(new_n397_), .A3(new_n420_), .ZN(new_n830_));
  OAI21_X1  g629(.A(KEYINPUT59), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n775_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n824_), .A2(new_n826_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n810_), .A2(new_n818_), .A3(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n832_), .B1(new_n835_), .B2(new_n628_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n830_), .A2(KEYINPUT59), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n831_), .A2(new_n838_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(KEYINPUT118), .B(G113gat), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n497_), .A2(new_n840_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(KEYINPUT119), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n839_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT116), .B1(new_n829_), .B2(new_n830_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT116), .ZN(new_n845_));
  INV_X1    g644(.A(new_n830_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n824_), .A2(new_n826_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n802_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n580_), .B1(new_n806_), .B2(new_n805_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(new_n808_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n847_), .B1(new_n850_), .B2(new_n801_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n825_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n852_));
  AOI211_X1 g651(.A(KEYINPUT114), .B(KEYINPUT57), .C1(new_n823_), .C2(new_n636_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n628_), .B1(new_n851_), .B2(new_n854_), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n845_), .B(new_n846_), .C1(new_n855_), .C2(new_n775_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n844_), .A2(new_n856_), .A3(new_n496_), .ZN(new_n857_));
  INV_X1    g656(.A(G113gat), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(KEYINPUT117), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT117), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n857_), .A2(new_n861_), .A3(new_n858_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n843_), .B1(new_n860_), .B2(new_n862_), .ZN(G1340gat));
  OAI21_X1  g662(.A(G120gat), .B1(new_n839_), .B2(new_n613_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT60), .ZN(new_n865_));
  AOI21_X1  g664(.A(G120gat), .B1(new_n639_), .B2(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n866_), .B1(new_n865_), .B2(G120gat), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n844_), .A2(new_n856_), .A3(new_n867_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n868_), .A2(KEYINPUT120), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n868_), .A2(KEYINPUT120), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n864_), .B1(new_n869_), .B2(new_n870_), .ZN(G1341gat));
  OAI21_X1  g670(.A(G127gat), .B1(new_n839_), .B2(new_n640_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n844_), .A2(new_n856_), .A3(new_n375_), .A4(new_n628_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(G1342gat));
  NOR3_X1   g673(.A1(new_n839_), .A2(new_n373_), .A3(new_n580_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n844_), .A2(new_n856_), .A3(new_n637_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n373_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n876_), .A2(KEYINPUT121), .A3(new_n373_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n875_), .B1(new_n879_), .B2(new_n880_), .ZN(G1343gat));
  NAND2_X1  g680(.A1(new_n828_), .A2(new_n640_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n832_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n449_), .A2(new_n445_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n302_), .A2(new_n452_), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n883_), .A2(new_n496_), .A3(new_n884_), .A4(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(KEYINPUT123), .ZN(new_n887_));
  INV_X1    g686(.A(new_n884_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n829_), .A2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT123), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n889_), .A2(new_n890_), .A3(new_n496_), .A4(new_n885_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT122), .B(G141gat), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n887_), .A2(new_n891_), .A3(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n892_), .B1(new_n887_), .B2(new_n891_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1344gat));
  NAND2_X1  g694(.A1(new_n889_), .A2(new_n885_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(new_n613_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(new_n307_), .ZN(G1345gat));
  NOR2_X1   g697(.A1(new_n896_), .A2(new_n640_), .ZN(new_n899_));
  XOR2_X1   g698(.A(KEYINPUT61), .B(G155gat), .Z(new_n900_));
  XNOR2_X1  g699(.A(new_n899_), .B(new_n900_), .ZN(G1346gat));
  INV_X1    g700(.A(G162gat), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n889_), .A2(new_n902_), .A3(new_n637_), .A4(new_n885_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n885_), .ZN(new_n904_));
  NOR4_X1   g703(.A1(new_n829_), .A2(new_n580_), .A3(new_n888_), .A4(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n903_), .B1(new_n902_), .B2(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n903_), .B(KEYINPUT124), .C1(new_n902_), .C2(new_n905_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(G1347gat));
  AOI21_X1  g709(.A(new_n775_), .B1(new_n834_), .B2(new_n640_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n301_), .A2(new_n420_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n913_), .A2(new_n456_), .A3(new_n362_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n911_), .A2(new_n497_), .A3(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n252_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT125), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n918_), .B(new_n919_), .C1(new_n916_), .C2(new_n229_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n918_), .B1(new_n916_), .B2(new_n229_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(KEYINPUT62), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n916_), .A2(new_n918_), .A3(new_n229_), .ZN(new_n923_));
  OAI211_X1 g722(.A(new_n917_), .B(new_n920_), .C1(new_n922_), .C2(new_n923_), .ZN(G1348gat));
  NOR2_X1   g723(.A1(new_n911_), .A2(new_n915_), .ZN(new_n925_));
  AOI21_X1  g724(.A(G176gat), .B1(new_n925_), .B2(new_n639_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n927_));
  NOR4_X1   g726(.A1(new_n829_), .A2(new_n230_), .A3(new_n613_), .A4(new_n915_), .ZN(new_n928_));
  OR3_X1    g727(.A1(new_n926_), .A2(new_n927_), .A3(new_n928_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n927_), .B1(new_n926_), .B2(new_n928_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(new_n930_), .ZN(G1349gat));
  INV_X1    g730(.A(new_n925_), .ZN(new_n932_));
  NOR3_X1   g731(.A1(new_n932_), .A2(new_n223_), .A3(new_n640_), .ZN(new_n933_));
  INV_X1    g732(.A(G183gat), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n883_), .A2(new_n628_), .A3(new_n914_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n933_), .B1(new_n934_), .B2(new_n935_), .ZN(G1350gat));
  OAI21_X1  g735(.A(G190gat), .B1(new_n932_), .B2(new_n580_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n925_), .A2(new_n224_), .A3(new_n637_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n937_), .A2(new_n938_), .ZN(G1351gat));
  NOR3_X1   g738(.A1(new_n829_), .A2(new_n888_), .A3(new_n913_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(new_n496_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g741(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n943_));
  XNOR2_X1  g742(.A(KEYINPUT127), .B(G204gat), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n940_), .A2(new_n639_), .ZN(new_n945_));
  MUX2_X1   g744(.A(new_n943_), .B(new_n944_), .S(new_n945_), .Z(G1353gat));
  AOI21_X1  g745(.A(new_n640_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n940_), .A2(new_n947_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n949_));
  XOR2_X1   g748(.A(new_n948_), .B(new_n949_), .Z(G1354gat));
  INV_X1    g749(.A(G218gat), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n940_), .A2(new_n951_), .A3(new_n637_), .ZN(new_n952_));
  AND2_X1   g751(.A1(new_n940_), .A2(new_n677_), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n952_), .B1(new_n953_), .B2(new_n951_), .ZN(G1355gat));
endmodule


