//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1 1 0 0 0 0 0 0 0 1 1 0 0 0 1 0 0 1 0 0 0 1 1 0 0 1 0 0 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n783_,
    new_n784_, new_n785_, new_n787_, new_n788_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n848_, new_n849_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_, new_n952_,
    new_n954_, new_n955_, new_n956_, new_n958_, new_n959_, new_n961_,
    new_n962_, new_n964_, new_n965_, new_n966_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n985_, new_n986_, new_n988_, new_n989_, new_n990_,
    new_n991_, new_n993_, new_n995_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1003_, new_n1004_;
  XOR2_X1   g000(.A(G1gat), .B(G29gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT103), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT0), .B(G57gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G225gat), .A2(G233gat), .ZN(new_n208_));
  INV_X1    g007(.A(G120gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G113gat), .ZN(new_n210_));
  INV_X1    g009(.A(G113gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G120gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT88), .ZN(new_n213_));
  AND3_X1   g012(.A1(new_n210_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n213_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G127gat), .B(G134gat), .ZN(new_n216_));
  NOR3_X1   g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  XOR2_X1   g016(.A(G127gat), .B(G134gat), .Z(new_n218_));
  NOR2_X1   g017(.A1(new_n211_), .A2(G120gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n209_), .A2(G113gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT88), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n210_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n218_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT89), .B1(new_n217_), .B2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n221_), .A2(new_n222_), .A3(new_n218_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT89), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G141gat), .A2(G148gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT92), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT2), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT2), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n228_), .A2(new_n229_), .A3(new_n232_), .ZN(new_n233_));
  OAI22_X1  g032(.A1(KEYINPUT91), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(KEYINPUT91), .A2(KEYINPUT3), .ZN(new_n235_));
  INV_X1    g034(.A(G141gat), .ZN(new_n236_));
  INV_X1    g035(.A(G148gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n231_), .A2(new_n233_), .A3(new_n234_), .A4(new_n238_), .ZN(new_n239_));
  XOR2_X1   g038(.A(G155gat), .B(G162gat), .Z(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n236_), .A2(new_n237_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT1), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n243_), .A2(G155gat), .A3(G162gat), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n244_), .B1(G155gat), .B2(G162gat), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n243_), .B1(G155gat), .B2(G162gat), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n228_), .B(new_n242_), .C1(new_n245_), .C2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n241_), .A2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n224_), .A2(new_n227_), .A3(new_n248_), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n241_), .B(new_n247_), .C1(new_n217_), .C2(new_n223_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(KEYINPUT4), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT101), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT101), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n249_), .A2(new_n253_), .A3(KEYINPUT4), .A4(new_n250_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT4), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n224_), .A2(new_n256_), .A3(new_n248_), .A4(new_n227_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT102), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n216_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n226_), .B1(new_n260_), .B2(new_n225_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n214_), .A2(new_n215_), .ZN(new_n262_));
  AOI21_X1  g061(.A(KEYINPUT89), .B1(new_n262_), .B2(new_n218_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n264_), .A2(KEYINPUT102), .A3(new_n256_), .A4(new_n248_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n259_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n208_), .B1(new_n255_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n249_), .A2(new_n250_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(new_n208_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n207_), .B1(new_n268_), .B2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n266_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n206_), .B(new_n270_), .C1(new_n273_), .C2(new_n208_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G226gat), .A2(G233gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT19), .ZN(new_n277_));
  NOR2_X1   g076(.A1(G197gat), .A2(G204gat), .ZN(new_n278_));
  INV_X1    g077(.A(G197gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT93), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT93), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(G197gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n278_), .B1(new_n283_), .B2(G204gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G211gat), .B(G218gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT21), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n284_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(G204gat), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n280_), .A2(new_n282_), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT94), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n286_), .B1(G197gat), .B2(G204gat), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n291_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n285_), .B1(new_n284_), .B2(KEYINPUT21), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n288_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT96), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n290_), .A2(new_n292_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT94), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n285_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n278_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT93), .B(G197gat), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n305_), .B1(new_n306_), .B2(new_n289_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n304_), .B1(new_n307_), .B2(new_n286_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n303_), .A2(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(KEYINPUT96), .B1(new_n309_), .B2(new_n288_), .ZN(new_n310_));
  INV_X1    g109(.A(G183gat), .ZN(new_n311_));
  INV_X1    g110(.A(G190gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT23), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT23), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(G183gat), .A3(G190gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n312_), .A2(KEYINPUT26), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT26), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(G190gat), .ZN(new_n319_));
  AND2_X1   g118(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n320_));
  NOR2_X1   g119(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n317_), .B(new_n319_), .C1(new_n320_), .C2(new_n321_), .ZN(new_n322_));
  OR3_X1    g121(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n323_));
  OR2_X1    g122(.A1(G169gat), .A2(G176gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G169gat), .A2(G176gat), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n324_), .A2(KEYINPUT24), .A3(new_n325_), .ZN(new_n326_));
  AND4_X1   g125(.A1(new_n316_), .A2(new_n322_), .A3(new_n323_), .A4(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT86), .B(G176gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT22), .B(G169gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT98), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n325_), .B(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n314_), .B1(G183gat), .B2(G190gat), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT85), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n315_), .A2(new_n335_), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n314_), .A2(KEYINPUT85), .A3(G183gat), .A4(G190gat), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n334_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(G183gat), .A2(G190gat), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n331_), .B(new_n333_), .C1(new_n338_), .C2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n328_), .A2(new_n340_), .ZN(new_n341_));
  NOR3_X1   g140(.A1(new_n299_), .A2(new_n310_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n339_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n316_), .A2(new_n343_), .ZN(new_n344_));
  AND3_X1   g143(.A1(new_n329_), .A2(new_n330_), .A3(KEYINPUT87), .ZN(new_n345_));
  AOI21_X1  g144(.A(KEYINPUT87), .B1(new_n329_), .B2(new_n330_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n325_), .B(new_n344_), .C1(new_n345_), .C2(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n311_), .A2(KEYINPUT23), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT85), .B1(new_n348_), .B2(G190gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n337_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n313_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT83), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n352_), .B1(new_n311_), .B2(KEYINPUT84), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT25), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n352_), .B(KEYINPUT25), .C1(new_n311_), .C2(KEYINPUT84), .ZN(new_n356_));
  NAND2_X1  g155(.A1(KEYINPUT83), .A2(G183gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT26), .B(G190gat), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n355_), .A2(new_n356_), .A3(new_n357_), .A4(new_n358_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n326_), .A2(new_n323_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n351_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n347_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  AND2_X1   g162(.A1(new_n284_), .A2(new_n287_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n364_), .B1(new_n303_), .B2(new_n308_), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT20), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n277_), .B1(new_n342_), .B2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT20), .B1(new_n297_), .B2(new_n362_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT97), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT99), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n351_), .A2(new_n343_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n331_), .A2(new_n333_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n327_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n370_), .B1(new_n365_), .B2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n297_), .A2(KEYINPUT99), .A3(new_n341_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT97), .ZN(new_n377_));
  OAI211_X1 g176(.A(new_n377_), .B(KEYINPUT20), .C1(new_n297_), .C2(new_n362_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n369_), .A2(new_n376_), .A3(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n367_), .B1(new_n277_), .B2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G8gat), .B(G36gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT18), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G64gat), .B(G92gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n385_), .A2(KEYINPUT32), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n380_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n379_), .A2(new_n277_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n277_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n389_), .B1(new_n297_), .B2(new_n341_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n366_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n388_), .A2(new_n392_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n275_), .B(new_n387_), .C1(new_n386_), .C2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT100), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n385_), .B1(new_n388_), .B2(new_n392_), .ZN(new_n396_));
  AOI211_X1 g195(.A(new_n384_), .B(new_n391_), .C1(new_n379_), .C2(new_n277_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n395_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  OAI211_X1 g197(.A(KEYINPUT33), .B(new_n207_), .C1(new_n268_), .C2(new_n271_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT33), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n272_), .A2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n398_), .A2(new_n399_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n393_), .A2(new_n384_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n388_), .A2(new_n385_), .A3(new_n392_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(KEYINPUT100), .A3(new_n404_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n273_), .A2(new_n208_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n206_), .B1(new_n269_), .B2(new_n208_), .ZN(new_n407_));
  OR2_X1    g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n405_), .A2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n394_), .B1(new_n402_), .B2(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n248_), .A2(KEYINPUT29), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT28), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G22gat), .B(G50gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  XOR2_X1   g214(.A(G78gat), .B(G106gat), .Z(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n241_), .A2(new_n247_), .ZN(new_n418_));
  XOR2_X1   g217(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  OAI22_X1  g219(.A1(new_n299_), .A2(new_n310_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(G228gat), .ZN(new_n422_));
  INV_X1    g221(.A(G233gat), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n421_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n248_), .A2(KEYINPUT29), .ZN(new_n426_));
  INV_X1    g225(.A(new_n424_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n297_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n417_), .B1(new_n425_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n428_), .ZN(new_n430_));
  AOI211_X1 g229(.A(new_n416_), .B(new_n430_), .C1(new_n421_), .C2(new_n424_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n415_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n414_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n413_), .B(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n297_), .A2(new_n298_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n365_), .A2(KEYINPUT96), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n435_), .A2(new_n436_), .B1(new_n248_), .B2(new_n419_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n428_), .B1(new_n437_), .B2(new_n427_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n416_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n425_), .A2(new_n417_), .A3(new_n428_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n434_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n432_), .A2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G71gat), .B(G99gat), .ZN(new_n443_));
  INV_X1    g242(.A(G43gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT30), .ZN(new_n446_));
  OR2_X1    g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n446_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G227gat), .A2(G233gat), .ZN(new_n449_));
  INV_X1    g248(.A(G15gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n447_), .A2(new_n448_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n451_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n362_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n445_), .B(new_n446_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n451_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n458_), .A2(new_n363_), .A3(new_n452_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n455_), .A2(KEYINPUT90), .A3(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n264_), .B(KEYINPUT31), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n442_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n410_), .A2(new_n463_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n432_), .A2(new_n462_), .A3(new_n441_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n462_), .B1(new_n432_), .B2(new_n441_), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n380_), .A2(new_n384_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(KEYINPUT27), .A3(new_n404_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT27), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n470_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n472_), .A2(new_n275_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n467_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n464_), .A2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G29gat), .B(G36gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G43gat), .B(G50gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT15), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G1gat), .B(G8gat), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n480_), .A2(KEYINPUT75), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(KEYINPUT75), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G15gat), .B(G22gat), .ZN(new_n484_));
  INV_X1    g283(.A(G1gat), .ZN(new_n485_));
  INV_X1    g284(.A(G8gat), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT14), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n484_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n483_), .A2(new_n488_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n481_), .A2(new_n487_), .A3(new_n484_), .A4(new_n482_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n479_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n489_), .A2(new_n478_), .A3(new_n490_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G229gat), .A2(G233gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n492_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n494_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n493_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n478_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n496_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G113gat), .B(G141gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G169gat), .B(G197gat), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n500_), .B(new_n501_), .Z(new_n502_));
  AND3_X1   g301(.A1(new_n495_), .A2(new_n499_), .A3(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n502_), .B1(new_n495_), .B2(new_n499_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n505_), .B(KEYINPUT82), .Z(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n475_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G232gat), .A2(G233gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT34), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT35), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n478_), .B(KEYINPUT15), .Z(new_n515_));
  NAND2_X1  g314(.A1(G99gat), .A2(G106gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT6), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT7), .ZN(new_n518_));
  INV_X1    g317(.A(G99gat), .ZN(new_n519_));
  INV_X1    g318(.A(G106gat), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .A4(KEYINPUT66), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n519_), .A2(new_n520_), .A3(KEYINPUT66), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT7), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n517_), .A2(new_n521_), .A3(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(G85gat), .B(G92gat), .Z(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT8), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT8), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n524_), .A2(new_n528_), .A3(new_n525_), .ZN(new_n529_));
  OR2_X1    g328(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT64), .ZN(new_n531_));
  NAND2_X1  g330(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n530_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n531_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n520_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT65), .ZN(new_n537_));
  INV_X1    g336(.A(G85gat), .ZN(new_n538_));
  INV_X1    g337(.A(G92gat), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n537_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n540_), .A2(KEYINPUT9), .B1(new_n538_), .B2(new_n539_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT9), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n537_), .B(new_n542_), .C1(new_n538_), .C2(new_n539_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n536_), .A2(new_n517_), .A3(new_n544_), .ZN(new_n545_));
  AOI22_X1  g344(.A1(new_n527_), .A2(new_n529_), .B1(new_n545_), .B2(KEYINPUT68), .ZN(new_n546_));
  INV_X1    g345(.A(new_n517_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT10), .B(G99gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT64), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(new_n533_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n547_), .B1(new_n550_), .B2(new_n520_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT68), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(new_n552_), .A3(new_n544_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n515_), .B1(new_n546_), .B2(new_n553_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n524_), .A2(new_n528_), .A3(new_n525_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n528_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n545_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n478_), .ZN(new_n558_));
  OAI22_X1  g357(.A1(new_n557_), .A2(new_n558_), .B1(KEYINPUT35), .B2(new_n510_), .ZN(new_n559_));
  NOR3_X1   g358(.A1(new_n554_), .A2(new_n559_), .A3(KEYINPUT70), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT70), .ZN(new_n561_));
  AOI22_X1  g360(.A1(new_n527_), .A2(new_n529_), .B1(new_n544_), .B2(new_n551_), .ZN(new_n562_));
  AOI22_X1  g361(.A1(new_n562_), .A2(new_n478_), .B1(new_n512_), .B2(new_n511_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n527_), .A2(new_n529_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n545_), .A2(KEYINPUT68), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n564_), .A2(new_n565_), .A3(new_n553_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(new_n479_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n561_), .B1(new_n563_), .B2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n514_), .B1(new_n560_), .B2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(KEYINPUT70), .B1(new_n554_), .B2(new_n559_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n563_), .A2(new_n567_), .A3(new_n561_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n570_), .A2(new_n571_), .A3(new_n513_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G190gat), .B(G218gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G134gat), .B(G162gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT36), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n569_), .A2(new_n572_), .A3(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(KEYINPUT74), .B(KEYINPUT37), .Z(new_n580_));
  NAND2_X1  g379(.A1(new_n569_), .A2(new_n572_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT36), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n577_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(KEYINPUT73), .B1(new_n581_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT73), .ZN(new_n586_));
  AOI211_X1 g385(.A(new_n586_), .B(new_n583_), .C1(new_n569_), .C2(new_n572_), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n579_), .B(new_n580_), .C1(new_n585_), .C2(new_n587_), .ZN(new_n588_));
  XOR2_X1   g387(.A(G127gat), .B(G155gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT16), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G183gat), .B(G211gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT17), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n593_), .A2(KEYINPUT78), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n592_), .A2(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n596_), .B1(new_n593_), .B2(new_n592_), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n489_), .A2(KEYINPUT76), .A3(new_n490_), .ZN(new_n598_));
  AOI21_X1  g397(.A(KEYINPUT76), .B1(new_n489_), .B2(new_n490_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(G231gat), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n600_), .B1(new_n601_), .B2(new_n423_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G57gat), .B(G64gat), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n603_), .A2(KEYINPUT11), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(KEYINPUT11), .ZN(new_n605_));
  XOR2_X1   g404(.A(G71gat), .B(G78gat), .Z(new_n606_));
  NAND3_X1  g405(.A1(new_n604_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n605_), .A2(new_n606_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n609_), .B(KEYINPUT77), .Z(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  OAI211_X1 g410(.A(G231gat), .B(G233gat), .C1(new_n598_), .C2(new_n599_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n602_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n611_), .B1(new_n602_), .B2(new_n612_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n597_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n602_), .A2(new_n612_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(new_n610_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n618_), .A2(new_n596_), .A3(new_n613_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT79), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n616_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n620_), .B1(new_n616_), .B2(new_n619_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n579_), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n570_), .A2(new_n513_), .A3(new_n571_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n513_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n584_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n586_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n581_), .A2(KEYINPUT73), .A3(new_n584_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n624_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(KEYINPUT74), .A2(KEYINPUT37), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n588_), .B(new_n623_), .C1(new_n630_), .C2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(KEYINPUT80), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT67), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n562_), .A2(new_n635_), .A3(new_n609_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n609_), .ZN(new_n637_));
  OAI21_X1  g436(.A(KEYINPUT67), .B1(new_n557_), .B2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n557_), .A2(new_n637_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n636_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(G230gat), .A2(G233gat), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT12), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n639_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n607_), .A2(KEYINPUT12), .A3(new_n608_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n566_), .A2(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n642_), .B1(new_n562_), .B2(new_n609_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n645_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n643_), .A2(new_n650_), .ZN(new_n651_));
  XOR2_X1   g450(.A(G120gat), .B(G148gat), .Z(new_n652_));
  XNOR2_X1  g451(.A(G176gat), .B(G204gat), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n651_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n643_), .A2(new_n650_), .A3(new_n656_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT13), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n658_), .A2(KEYINPUT13), .A3(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n579_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(new_n631_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT80), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n667_), .A2(new_n668_), .A3(new_n588_), .A4(new_n623_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n634_), .A2(new_n665_), .A3(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n508_), .B1(new_n670_), .B2(KEYINPUT81), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT81), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n634_), .A2(new_n672_), .A3(new_n665_), .A4(new_n669_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n675_), .A2(new_n485_), .A3(new_n275_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n616_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n619_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n505_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n665_), .A2(new_n681_), .A3(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n475_), .A2(KEYINPUT105), .A3(new_n666_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n685_));
  AOI22_X1  g484(.A1(new_n410_), .A2(new_n463_), .B1(new_n467_), .B2(new_n473_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n685_), .B1(new_n686_), .B2(new_n630_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n683_), .B1(new_n684_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n275_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G1gat), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n676_), .A2(new_n677_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n678_), .A2(new_n691_), .A3(new_n692_), .ZN(G1324gat));
  XNOR2_X1  g492(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT39), .ZN(new_n695_));
  AOI211_X1 g494(.A(new_n695_), .B(new_n486_), .C1(new_n688_), .C2(new_n472_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n684_), .A2(new_n687_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n683_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n697_), .A2(new_n472_), .A3(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(KEYINPUT39), .B1(new_n699_), .B2(G8gat), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n696_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n670_), .A2(KEYINPUT81), .ZN(new_n702_));
  INV_X1    g501(.A(new_n508_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n472_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n704_), .A2(G8gat), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n702_), .A2(new_n673_), .A3(new_n703_), .A4(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT106), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n671_), .A2(KEYINPUT106), .A3(new_n673_), .A4(new_n705_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n694_), .B1(new_n701_), .B2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n699_), .A2(G8gat), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n695_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n699_), .A2(KEYINPUT39), .A3(G8gat), .ZN(new_n714_));
  AND4_X1   g513(.A1(new_n710_), .A2(new_n713_), .A3(new_n714_), .A4(new_n694_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n711_), .A2(new_n715_), .ZN(G1325gat));
  NAND3_X1  g515(.A1(new_n675_), .A2(new_n450_), .A3(new_n462_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n688_), .A2(new_n462_), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT41), .B1(new_n718_), .B2(G15gat), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT41), .ZN(new_n720_));
  AOI211_X1 g519(.A(new_n720_), .B(new_n450_), .C1(new_n688_), .C2(new_n462_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n719_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT108), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n717_), .B(new_n724_), .C1(new_n719_), .C2(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1326gat));
  INV_X1    g525(.A(new_n442_), .ZN(new_n727_));
  OR3_X1    g526(.A1(new_n674_), .A2(G22gat), .A3(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(G22gat), .B1(new_n689_), .B2(new_n727_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n729_), .A2(KEYINPUT42), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(KEYINPUT42), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n728_), .B1(new_n730_), .B2(new_n731_), .ZN(G1327gat));
  NOR3_X1   g531(.A1(new_n666_), .A2(new_n623_), .A3(new_n664_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n463_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n406_), .A2(new_n407_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n396_), .A2(new_n397_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n736_), .B2(KEYINPUT100), .ZN(new_n737_));
  INV_X1    g536(.A(new_n399_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n270_), .B1(new_n273_), .B2(new_n208_), .ZN(new_n739_));
  AOI21_X1  g538(.A(KEYINPUT33), .B1(new_n739_), .B2(new_n207_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n738_), .A2(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n737_), .A2(new_n741_), .A3(new_n398_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n734_), .B1(new_n742_), .B2(new_n394_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n465_), .A2(new_n466_), .ZN(new_n744_));
  NOR3_X1   g543(.A1(new_n744_), .A2(new_n275_), .A3(new_n472_), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n507_), .B(new_n733_), .C1(new_n743_), .C2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT109), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n475_), .A2(KEYINPUT109), .A3(new_n507_), .A4(new_n733_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(G29gat), .B1(new_n750_), .B2(new_n275_), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n623_), .A2(new_n664_), .A3(new_n505_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n630_), .A2(new_n632_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n588_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n755_), .A2(new_n686_), .A3(KEYINPUT43), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT43), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n667_), .A2(new_n588_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n475_), .B2(new_n758_), .ZN(new_n759_));
  OAI211_X1 g558(.A(KEYINPUT44), .B(new_n752_), .C1(new_n756_), .C2(new_n759_), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n760_), .A2(G29gat), .A3(new_n275_), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT43), .B1(new_n755_), .B2(new_n686_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n475_), .A2(new_n757_), .A3(new_n758_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(KEYINPUT44), .B1(new_n764_), .B2(new_n752_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n751_), .B1(new_n761_), .B2(new_n766_), .ZN(G1328gat));
  NAND2_X1  g566(.A1(new_n760_), .A2(new_n472_), .ZN(new_n768_));
  OAI21_X1  g567(.A(G36gat), .B1(new_n768_), .B2(new_n765_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n704_), .A2(G36gat), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n748_), .A2(new_n749_), .A3(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT110), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n748_), .A2(new_n749_), .A3(new_n774_), .A4(new_n770_), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n772_), .A2(new_n773_), .A3(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n773_), .B1(new_n772_), .B2(new_n775_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n769_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT46), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n769_), .B(KEYINPUT46), .C1(new_n776_), .C2(new_n777_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(G1329gat));
  AND2_X1   g581(.A1(new_n750_), .A2(new_n462_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n760_), .A2(G43gat), .A3(new_n462_), .ZN(new_n784_));
  OAI22_X1  g583(.A1(new_n783_), .A2(G43gat), .B1(new_n784_), .B2(new_n765_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g585(.A(G50gat), .B1(new_n750_), .B2(new_n442_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n760_), .A2(G50gat), .A3(new_n442_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n787_), .B1(new_n788_), .B2(new_n766_), .ZN(G1331gat));
  NAND3_X1  g588(.A1(new_n623_), .A2(new_n664_), .A3(new_n506_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n684_), .B2(new_n687_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(G57gat), .B1(new_n792_), .B2(new_n690_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n634_), .A2(new_n664_), .A3(new_n669_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n795_));
  OR2_X1    g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n686_), .A2(new_n682_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n794_), .A2(new_n795_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n796_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n799_));
  OR2_X1    g598(.A1(new_n690_), .A2(G57gat), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n793_), .B1(new_n799_), .B2(new_n800_), .ZN(G1332gat));
  OR3_X1    g600(.A1(new_n799_), .A2(G64gat), .A3(new_n704_), .ZN(new_n802_));
  OAI21_X1  g601(.A(G64gat), .B1(new_n792_), .B2(new_n704_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n803_), .A2(KEYINPUT48), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n803_), .A2(KEYINPUT48), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n802_), .B1(new_n804_), .B2(new_n805_), .ZN(G1333gat));
  XNOR2_X1  g605(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n791_), .A2(new_n462_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n807_), .B1(new_n808_), .B2(G71gat), .ZN(new_n809_));
  INV_X1    g608(.A(G71gat), .ZN(new_n810_));
  INV_X1    g609(.A(new_n807_), .ZN(new_n811_));
  AOI211_X1 g610(.A(new_n810_), .B(new_n811_), .C1(new_n791_), .C2(new_n462_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n462_), .A2(new_n810_), .ZN(new_n813_));
  OAI22_X1  g612(.A1(new_n809_), .A2(new_n812_), .B1(new_n799_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT113), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT113), .ZN(new_n816_));
  OAI221_X1 g615(.A(new_n816_), .B1(new_n799_), .B2(new_n813_), .C1(new_n809_), .C2(new_n812_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(G1334gat));
  OAI21_X1  g617(.A(G78gat), .B1(new_n792_), .B2(new_n727_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n819_), .A2(KEYINPUT50), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n819_), .A2(KEYINPUT50), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n727_), .A2(G78gat), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(KEYINPUT114), .ZN(new_n823_));
  OAI22_X1  g622(.A1(new_n820_), .A2(new_n821_), .B1(new_n799_), .B2(new_n823_), .ZN(G1335gat));
  INV_X1    g623(.A(new_n623_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(new_n664_), .A3(new_n505_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n826_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(G85gat), .B1(new_n828_), .B2(new_n690_), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n665_), .A2(new_n666_), .A3(new_n623_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n797_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(new_n538_), .A3(new_n275_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n829_), .A2(new_n833_), .ZN(G1336gat));
  AOI21_X1  g633(.A(G92gat), .B1(new_n832_), .B2(new_n472_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n472_), .A2(G92gat), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(KEYINPUT115), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n835_), .B1(new_n827_), .B2(new_n837_), .ZN(G1337gat));
  INV_X1    g637(.A(new_n462_), .ZN(new_n839_));
  OAI21_X1  g638(.A(G99gat), .B1(new_n828_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n462_), .A2(new_n550_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n831_), .A2(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n842_), .A2(KEYINPUT116), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n831_), .A2(new_n844_), .A3(new_n841_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n840_), .B1(new_n843_), .B2(new_n845_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g646(.A1(new_n832_), .A2(new_n520_), .A3(new_n442_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT117), .B(KEYINPUT52), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n827_), .A2(new_n442_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(G106gat), .ZN(new_n852_));
  AOI211_X1 g651(.A(new_n520_), .B(new_n849_), .C1(new_n827_), .C2(new_n442_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n848_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(KEYINPUT53), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n856_), .B(new_n848_), .C1(new_n852_), .C2(new_n853_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(G1339gat));
  NOR2_X1   g657(.A1(new_n472_), .A2(new_n690_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n465_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n492_), .A2(new_n493_), .A3(new_n496_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n491_), .A2(new_n558_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n496_), .B1(new_n862_), .B2(new_n493_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n863_), .A2(new_n864_), .A3(new_n502_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n494_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n502_), .ZN(new_n867_));
  AOI21_X1  g666(.A(KEYINPUT121), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n861_), .B1(new_n865_), .B2(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n503_), .B1(new_n869_), .B2(KEYINPUT122), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT122), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n871_), .B(new_n861_), .C1(new_n865_), .C2(new_n868_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n659_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT119), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT55), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n650_), .B2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n645_), .A2(new_n648_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n636_), .A2(new_n638_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n642_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n650_), .A2(new_n877_), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n644_), .A2(new_n639_), .B1(new_n566_), .B2(new_n647_), .ZN(new_n883_));
  NAND4_X1  g682(.A1(new_n883_), .A2(KEYINPUT119), .A3(KEYINPUT55), .A4(new_n649_), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n878_), .A2(new_n881_), .A3(new_n882_), .A4(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n885_), .A2(KEYINPUT56), .A3(new_n657_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(KEYINPUT56), .B1(new_n885_), .B2(new_n657_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n875_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT58), .ZN(new_n890_));
  AOI22_X1  g689(.A1(new_n667_), .A2(new_n588_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  OR2_X1    g690(.A1(new_n889_), .A2(new_n890_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT57), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n885_), .A2(new_n657_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT56), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n897_), .A2(KEYINPUT120), .A3(new_n886_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n885_), .A2(new_n899_), .A3(KEYINPUT56), .A4(new_n657_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n874_), .A2(new_n505_), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n898_), .A2(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n873_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n905_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n894_), .B1(new_n906_), .B2(new_n666_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n904_), .B1(new_n898_), .B2(new_n902_), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n908_), .A2(KEYINPUT57), .A3(new_n630_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n893_), .B1(new_n907_), .B2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n681_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  AND3_X1   g711(.A1(new_n506_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n667_), .A2(new_n588_), .A3(new_n913_), .A4(new_n623_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n914_), .B(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n860_), .B1(new_n912_), .B2(new_n916_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n917_), .A2(new_n211_), .A3(new_n682_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT59), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n906_), .A2(new_n894_), .A3(new_n666_), .ZN(new_n920_));
  OAI21_X1  g719(.A(KEYINPUT57), .B1(new_n908_), .B2(new_n630_), .ZN(new_n921_));
  AOI22_X1  g720(.A1(new_n920_), .A2(new_n921_), .B1(new_n892_), .B2(new_n891_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n916_), .B1(new_n922_), .B2(new_n681_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n860_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n919_), .B1(new_n923_), .B2(new_n924_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n919_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n910_), .A2(new_n825_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n926_), .B1(new_n927_), .B2(new_n916_), .ZN(new_n928_));
  NOR3_X1   g727(.A1(new_n925_), .A2(new_n928_), .A3(new_n506_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n918_), .B1(new_n929_), .B2(new_n211_), .ZN(G1340gat));
  NOR3_X1   g729(.A1(new_n925_), .A2(new_n928_), .A3(new_n665_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n923_), .A2(new_n924_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n209_), .B1(new_n665_), .B2(KEYINPUT60), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n933_), .B1(KEYINPUT60), .B2(new_n209_), .ZN(new_n934_));
  OAI22_X1  g733(.A1(new_n931_), .A2(new_n209_), .B1(new_n932_), .B2(new_n934_), .ZN(G1341gat));
  INV_X1    g734(.A(KEYINPUT123), .ZN(new_n936_));
  INV_X1    g735(.A(G127gat), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n911_), .A2(new_n937_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n938_), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n925_), .A2(new_n928_), .A3(new_n939_), .ZN(new_n940_));
  AOI21_X1  g739(.A(G127gat), .B1(new_n917_), .B2(new_n623_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n936_), .B1(new_n940_), .B2(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n927_), .A2(new_n916_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n860_), .A2(KEYINPUT59), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n943_), .A2(new_n944_), .ZN(new_n945_));
  OAI211_X1 g744(.A(new_n945_), .B(new_n938_), .C1(new_n919_), .C2(new_n917_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n937_), .B1(new_n932_), .B2(new_n825_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n946_), .A2(new_n947_), .A3(KEYINPUT123), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n942_), .A2(new_n948_), .ZN(G1342gat));
  INV_X1    g748(.A(G134gat), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n917_), .A2(new_n950_), .A3(new_n630_), .ZN(new_n951_));
  NOR3_X1   g750(.A1(new_n925_), .A2(new_n928_), .A3(new_n755_), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n951_), .B1(new_n952_), .B2(new_n950_), .ZN(G1343gat));
  AND2_X1   g752(.A1(new_n923_), .A2(new_n466_), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n954_), .A2(new_n682_), .A3(new_n859_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(KEYINPUT124), .B(G141gat), .ZN(new_n956_));
  XNOR2_X1  g755(.A(new_n955_), .B(new_n956_), .ZN(G1344gat));
  NAND3_X1  g756(.A1(new_n954_), .A2(new_n664_), .A3(new_n859_), .ZN(new_n958_));
  XNOR2_X1  g757(.A(KEYINPUT125), .B(G148gat), .ZN(new_n959_));
  XNOR2_X1  g758(.A(new_n958_), .B(new_n959_), .ZN(G1345gat));
  NAND3_X1  g759(.A1(new_n954_), .A2(new_n623_), .A3(new_n859_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(KEYINPUT61), .B(G155gat), .ZN(new_n962_));
  XNOR2_X1  g761(.A(new_n961_), .B(new_n962_), .ZN(G1346gat));
  NAND2_X1  g762(.A1(new_n954_), .A2(new_n859_), .ZN(new_n964_));
  OAI21_X1  g763(.A(G162gat), .B1(new_n964_), .B2(new_n755_), .ZN(new_n965_));
  OR2_X1    g764(.A1(new_n666_), .A2(G162gat), .ZN(new_n966_));
  OAI21_X1  g765(.A(new_n965_), .B1(new_n964_), .B2(new_n966_), .ZN(G1347gat));
  NOR2_X1   g766(.A1(new_n704_), .A2(new_n275_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n968_), .A2(new_n462_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(new_n969_), .A2(new_n442_), .ZN(new_n970_));
  NAND3_X1  g769(.A1(new_n943_), .A2(new_n682_), .A3(new_n970_), .ZN(new_n971_));
  INV_X1    g770(.A(KEYINPUT62), .ZN(new_n972_));
  AND3_X1   g771(.A1(new_n971_), .A2(new_n972_), .A3(G169gat), .ZN(new_n973_));
  AOI21_X1  g772(.A(new_n972_), .B1(new_n971_), .B2(G169gat), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n943_), .A2(new_n970_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n682_), .A2(new_n330_), .ZN(new_n976_));
  XOR2_X1   g775(.A(new_n976_), .B(KEYINPUT126), .Z(new_n977_));
  OAI22_X1  g776(.A1(new_n973_), .A2(new_n974_), .B1(new_n975_), .B2(new_n977_), .ZN(G1348gat));
  INV_X1    g777(.A(new_n975_), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n979_), .A2(new_n664_), .ZN(new_n980_));
  AOI21_X1  g779(.A(new_n442_), .B1(new_n912_), .B2(new_n916_), .ZN(new_n981_));
  INV_X1    g780(.A(G176gat), .ZN(new_n982_));
  NOR3_X1   g781(.A1(new_n969_), .A2(new_n982_), .A3(new_n665_), .ZN(new_n983_));
  AOI22_X1  g782(.A1(new_n980_), .A2(new_n329_), .B1(new_n981_), .B2(new_n983_), .ZN(G1349gat));
  NAND4_X1  g783(.A1(new_n981_), .A2(new_n623_), .A3(new_n462_), .A4(new_n968_), .ZN(new_n985_));
  NOR3_X1   g784(.A1(new_n911_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n986_));
  AOI22_X1  g785(.A1(new_n985_), .A2(new_n311_), .B1(new_n979_), .B2(new_n986_), .ZN(G1350gat));
  NAND3_X1  g786(.A1(new_n979_), .A2(new_n630_), .A3(new_n358_), .ZN(new_n988_));
  NAND3_X1  g787(.A1(new_n943_), .A2(new_n758_), .A3(new_n970_), .ZN(new_n989_));
  AND3_X1   g788(.A1(new_n989_), .A2(KEYINPUT127), .A3(G190gat), .ZN(new_n990_));
  AOI21_X1  g789(.A(KEYINPUT127), .B1(new_n989_), .B2(G190gat), .ZN(new_n991_));
  OAI21_X1  g790(.A(new_n988_), .B1(new_n990_), .B2(new_n991_), .ZN(G1351gat));
  NAND3_X1  g791(.A1(new_n954_), .A2(new_n682_), .A3(new_n968_), .ZN(new_n993_));
  XNOR2_X1  g792(.A(new_n993_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g793(.A1(new_n954_), .A2(new_n664_), .A3(new_n968_), .ZN(new_n995_));
  XNOR2_X1  g794(.A(new_n995_), .B(G204gat), .ZN(G1353gat));
  XNOR2_X1  g795(.A(KEYINPUT63), .B(G211gat), .ZN(new_n997_));
  NAND4_X1  g796(.A1(new_n954_), .A2(new_n681_), .A3(new_n968_), .A4(new_n997_), .ZN(new_n998_));
  NAND2_X1  g797(.A1(new_n954_), .A2(new_n968_), .ZN(new_n999_));
  NOR2_X1   g798(.A1(new_n999_), .A2(new_n911_), .ZN(new_n1000_));
  NOR2_X1   g799(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1001_));
  OAI21_X1  g800(.A(new_n998_), .B1(new_n1000_), .B2(new_n1001_), .ZN(G1354gat));
  OAI21_X1  g801(.A(G218gat), .B1(new_n999_), .B2(new_n755_), .ZN(new_n1003_));
  OR2_X1    g802(.A1(new_n666_), .A2(G218gat), .ZN(new_n1004_));
  OAI21_X1  g803(.A(new_n1003_), .B1(new_n999_), .B2(new_n1004_), .ZN(G1355gat));
endmodule


