//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 0 1 0 1 1 0 1 0 0 0 0 1 0 0 1 1 1 1 0 1 1 0 1 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n822_, new_n823_, new_n825_, new_n826_, new_n827_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n947_, new_n948_,
    new_n949_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n980_, new_n981_, new_n983_,
    new_n984_, new_n985_, new_n986_, new_n987_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n993_, new_n995_, new_n996_,
    new_n998_, new_n999_, new_n1000_, new_n1002_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1009_, new_n1010_, new_n1011_, new_n1012_,
    new_n1013_, new_n1014_, new_n1015_, new_n1016_;
  INV_X1    g000(.A(KEYINPUT93), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT21), .ZN(new_n203_));
  INV_X1    g002(.A(G211gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(G218gat), .ZN(new_n205_));
  INV_X1    g004(.A(G218gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(G211gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n203_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G197gat), .B(G204gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n206_), .A2(G211gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n204_), .A2(G218gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n211_), .A2(new_n212_), .A3(KEYINPUT21), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n208_), .A2(new_n210_), .A3(new_n213_), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n209_), .A2(KEYINPUT21), .A3(new_n211_), .A4(new_n212_), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT23), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n219_), .A2(G183gat), .A3(G190gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n218_), .A2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n221_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(G183gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT25), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT25), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(G183gat), .ZN(new_n230_));
  INV_X1    g029(.A(G190gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT26), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT26), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(G190gat), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n228_), .A2(new_n230_), .A3(new_n232_), .A4(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(G169gat), .ZN(new_n236_));
  INV_X1    g035(.A(G176gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G169gat), .A2(G176gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(KEYINPUT24), .A3(new_n239_), .ZN(new_n240_));
  AND3_X1   g039(.A1(new_n235_), .A2(KEYINPUT92), .A3(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(KEYINPUT92), .B1(new_n235_), .B2(new_n240_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n226_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n239_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT22), .B(G169gat), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n244_), .B1(new_n245_), .B2(new_n237_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT80), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n218_), .A2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n217_), .A2(KEYINPUT80), .A3(KEYINPUT23), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT81), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n220_), .A2(new_n250_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n219_), .A2(KEYINPUT81), .A3(G183gat), .A4(G190gat), .ZN(new_n252_));
  AOI22_X1  g051(.A1(new_n248_), .A2(new_n249_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n227_), .A2(new_n231_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n246_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n216_), .B1(new_n243_), .B2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n221_), .A2(new_n254_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n246_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT79), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n239_), .A2(KEYINPUT24), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n260_), .B1(new_n261_), .B2(new_n222_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n238_), .A2(KEYINPUT79), .A3(KEYINPUT24), .A4(new_n239_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n262_), .A2(new_n235_), .A3(new_n263_), .A4(new_n224_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n259_), .B1(new_n264_), .B2(new_n253_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n214_), .A2(new_n215_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT20), .ZN(new_n268_));
  NOR3_X1   g067(.A1(new_n257_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G226gat), .A2(G233gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT19), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n202_), .B1(new_n269_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n235_), .A2(new_n240_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT92), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n235_), .A2(KEYINPUT92), .A3(new_n240_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n225_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n246_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n248_), .A2(new_n249_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n251_), .A2(new_n252_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n279_), .B1(new_n282_), .B2(new_n254_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n266_), .B1(new_n278_), .B2(new_n283_), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n216_), .B(new_n259_), .C1(new_n253_), .C2(new_n264_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n284_), .A2(KEYINPUT20), .A3(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n286_), .A2(KEYINPUT93), .A3(new_n271_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n243_), .A2(new_n216_), .A3(new_n256_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n265_), .A2(new_n266_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(KEYINPUT20), .A3(new_n289_), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n290_), .A2(new_n271_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n273_), .A2(new_n287_), .A3(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G8gat), .B(G36gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT18), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(G64gat), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n295_), .A2(G92gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(G92gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n292_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n298_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n273_), .A2(new_n300_), .A3(new_n287_), .A4(new_n291_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT27), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT96), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n269_), .A2(new_n305_), .A3(new_n272_), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n284_), .A2(KEYINPUT20), .A3(new_n285_), .A4(new_n272_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT96), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n290_), .A2(new_n271_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n306_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(new_n298_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n311_), .A2(KEYINPUT27), .A3(new_n301_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n304_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT98), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT98), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n304_), .A2(new_n315_), .A3(new_n312_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n318_));
  NAND3_X1  g117(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT2), .ZN(new_n321_));
  INV_X1    g120(.A(G141gat), .ZN(new_n322_));
  INV_X1    g121(.A(G148gat), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n321_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  NOR4_X1   g123(.A1(KEYINPUT85), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT85), .ZN(new_n326_));
  NOR2_X1   g125(.A1(G141gat), .A2(G148gat), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT3), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n326_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n320_), .B(new_n324_), .C1(new_n325_), .C2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT86), .ZN(new_n331_));
  AND2_X1   g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332_));
  NOR2_X1   g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n331_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  OR2_X1    g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(KEYINPUT86), .A3(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n330_), .A2(new_n334_), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT1), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n333_), .B1(new_n332_), .B2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n336_), .A2(KEYINPUT1), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT83), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT83), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n336_), .A2(new_n343_), .A3(KEYINPUT1), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n340_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n322_), .A2(new_n323_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n346_), .A2(new_n327_), .ZN(new_n347_));
  AND3_X1   g146(.A1(new_n345_), .A2(KEYINPUT84), .A3(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT84), .B1(new_n345_), .B2(new_n347_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n338_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n216_), .B1(new_n350_), .B2(KEYINPUT29), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G228gat), .A2(G233gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT88), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT87), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n337_), .A2(new_n334_), .ZN(new_n356_));
  NOR3_X1   g155(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(new_n326_), .ZN(new_n358_));
  AND3_X1   g157(.A1(new_n324_), .A2(new_n319_), .A3(new_n318_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n356_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT84), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n335_), .B1(KEYINPUT1), .B2(new_n336_), .ZN(new_n362_));
  AND3_X1   g161(.A1(new_n336_), .A2(new_n343_), .A3(KEYINPUT1), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n343_), .B1(new_n336_), .B2(KEYINPUT1), .ZN(new_n364_));
  NOR3_X1   g163(.A1(new_n362_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n347_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n361_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n345_), .A2(KEYINPUT84), .A3(new_n347_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n360_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT29), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n355_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n350_), .A2(KEYINPUT87), .A3(KEYINPUT29), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n266_), .A2(new_n353_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n371_), .A2(new_n372_), .A3(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT89), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n350_), .A2(KEYINPUT29), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n373_), .B1(new_n378_), .B2(new_n355_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(KEYINPUT89), .A3(new_n372_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n354_), .B1(new_n377_), .B2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G78gat), .B(G106gat), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n369_), .A2(new_n370_), .ZN(new_n384_));
  XOR2_X1   g183(.A(G22gat), .B(G50gat), .Z(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT28), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n384_), .B(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n387_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n383_), .A2(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n375_), .A2(new_n376_), .ZN(new_n390_));
  AOI21_X1  g189(.A(KEYINPUT89), .B1(new_n379_), .B2(new_n372_), .ZN(new_n391_));
  OAI22_X1  g190(.A1(new_n390_), .A2(new_n391_), .B1(new_n353_), .B2(new_n351_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n382_), .A2(KEYINPUT90), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n387_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n395_));
  AOI211_X1 g194(.A(new_n354_), .B(new_n394_), .C1(new_n377_), .C2(new_n380_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n395_), .A2(KEYINPUT91), .A3(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT91), .ZN(new_n399_));
  INV_X1    g198(.A(new_n387_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n400_), .B1(new_n381_), .B2(new_n393_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n399_), .B1(new_n401_), .B2(new_n396_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n389_), .B1(new_n398_), .B2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G1gat), .B(G29gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(KEYINPUT0), .ZN(new_n405_));
  INV_X1    g204(.A(G57gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(G85gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G225gat), .A2(G233gat), .ZN(new_n410_));
  XOR2_X1   g209(.A(G127gat), .B(G134gat), .Z(new_n411_));
  XOR2_X1   g210(.A(G113gat), .B(G120gat), .Z(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n350_), .A2(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n415_), .A2(KEYINPUT4), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n338_), .B(new_n413_), .C1(new_n348_), .C2(new_n349_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n415_), .A2(KEYINPUT4), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT94), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n415_), .A2(KEYINPUT94), .A3(KEYINPUT4), .A4(new_n417_), .ZN(new_n421_));
  AOI211_X1 g220(.A(new_n410_), .B(new_n416_), .C1(new_n420_), .C2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n415_), .A2(new_n417_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n410_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n409_), .B1(new_n422_), .B2(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n416_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n424_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n425_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n409_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n426_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n265_), .B(KEYINPUT30), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G227gat), .A2(G233gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT82), .ZN(new_n436_));
  XOR2_X1   g235(.A(G71gat), .B(G99gat), .Z(new_n437_));
  XOR2_X1   g236(.A(new_n436_), .B(new_n437_), .Z(new_n438_));
  XNOR2_X1  g237(.A(new_n434_), .B(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(new_n414_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G15gat), .B(G43gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT31), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n440_), .B(new_n442_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n317_), .A2(new_n403_), .A3(new_n433_), .A4(new_n443_), .ZN(new_n444_));
  OR2_X1    g243(.A1(new_n383_), .A2(new_n388_), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT91), .B1(new_n395_), .B2(new_n397_), .ZN(new_n446_));
  NOR3_X1   g245(.A1(new_n401_), .A2(new_n399_), .A3(new_n396_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n445_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n433_), .A2(new_n304_), .A3(new_n312_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT33), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n302_), .B1(new_n451_), .B2(new_n431_), .ZN(new_n452_));
  AOI211_X1 g251(.A(new_n425_), .B(new_n409_), .C1(new_n427_), .C2(new_n424_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n409_), .B1(new_n423_), .B2(new_n410_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n454_), .B1(new_n427_), .B2(new_n410_), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT33), .B1(new_n453_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n452_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n398_), .A2(new_n402_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n296_), .A2(KEYINPUT32), .A3(new_n297_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n273_), .A2(new_n287_), .A3(new_n291_), .A4(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT95), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n459_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n310_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT95), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n462_), .B1(new_n465_), .B2(new_n460_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n432_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n457_), .A2(new_n458_), .A3(new_n467_), .A4(new_n445_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n443_), .ZN(new_n469_));
  AND4_X1   g268(.A1(KEYINPUT97), .A2(new_n450_), .A3(new_n468_), .A4(new_n469_), .ZN(new_n470_));
  AOI22_X1  g269(.A1(new_n452_), .A2(new_n456_), .B1(new_n466_), .B2(new_n432_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n443_), .B1(new_n471_), .B2(new_n403_), .ZN(new_n472_));
  AOI21_X1  g271(.A(KEYINPUT97), .B1(new_n472_), .B2(new_n450_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n444_), .B1(new_n470_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G229gat), .A2(G233gat), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G29gat), .B(G36gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(G43gat), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT68), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(G50gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  OR2_X1    g281(.A1(new_n478_), .A2(new_n479_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n478_), .A2(new_n479_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(G50gat), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n482_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT76), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G15gat), .B(G22gat), .Z(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT74), .B(G8gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(G1gat), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n489_), .B1(new_n491_), .B2(KEYINPUT14), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(G1gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(G8gat), .ZN(new_n494_));
  INV_X1    g293(.A(G1gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n492_), .B(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(G8gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n494_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n482_), .A2(KEYINPUT76), .A3(new_n485_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n488_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n501_), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT76), .B1(new_n482_), .B2(new_n485_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n499_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT77), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n488_), .A2(new_n501_), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT77), .B1(new_n508_), .B2(new_n499_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n476_), .B(new_n502_), .C1(new_n507_), .C2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G113gat), .B(G141gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(G197gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT78), .B(G169gat), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n512_), .B(new_n513_), .Z(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n505_), .A2(new_n506_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n508_), .A2(KEYINPUT77), .A3(new_n499_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT15), .ZN(new_n518_));
  INV_X1    g317(.A(new_n485_), .ZN(new_n519_));
  AOI21_X1  g318(.A(G50gat), .B1(new_n483_), .B2(new_n484_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n518_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n482_), .A2(KEYINPUT15), .A3(new_n485_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  AOI22_X1  g322(.A1(new_n516_), .A2(new_n517_), .B1(new_n500_), .B2(new_n523_), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n510_), .B(new_n515_), .C1(new_n476_), .C2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n523_), .A2(new_n500_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n527_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(new_n475_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n515_), .B1(new_n529_), .B2(new_n510_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n526_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G120gat), .B(G148gat), .ZN(new_n532_));
  INV_X1    g331(.A(G204gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT5), .B(G176gat), .ZN(new_n535_));
  XOR2_X1   g334(.A(new_n534_), .B(new_n535_), .Z(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G99gat), .A2(G106gat), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT6), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT64), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n538_), .B(KEYINPUT6), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT64), .ZN(new_n544_));
  NOR2_X1   g343(.A1(G99gat), .A2(G106gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT7), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n542_), .A2(new_n544_), .A3(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(G85gat), .B(G92gat), .Z(new_n548_));
  INV_X1    g347(.A(KEYINPUT8), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n547_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n546_), .A2(new_n543_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(new_n548_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT8), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n551_), .A2(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n542_), .A2(new_n544_), .ZN(new_n556_));
  XOR2_X1   g355(.A(KEYINPUT10), .B(G99gat), .Z(new_n557_));
  INV_X1    g356(.A(G106gat), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n548_), .A2(KEYINPUT9), .ZN(new_n560_));
  INV_X1    g359(.A(G92gat), .ZN(new_n561_));
  OR3_X1    g360(.A1(new_n408_), .A2(new_n561_), .A3(KEYINPUT9), .ZN(new_n562_));
  AND3_X1   g361(.A1(new_n559_), .A2(new_n560_), .A3(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n556_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n555_), .A2(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(G71gat), .B(G78gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(G57gat), .B(G64gat), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n566_), .B1(KEYINPUT11), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(KEYINPUT11), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(KEYINPUT65), .A2(KEYINPUT12), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n565_), .A2(new_n570_), .A3(new_n572_), .ZN(new_n573_));
  AOI22_X1  g372(.A1(new_n551_), .A2(new_n554_), .B1(new_n556_), .B2(new_n563_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n570_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  AND2_X1   g375(.A1(KEYINPUT65), .A2(KEYINPUT12), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n577_), .A2(new_n571_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n573_), .B1(new_n576_), .B2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT66), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n574_), .A2(new_n575_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G230gat), .A2(G233gat), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n580_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n582_), .ZN(new_n585_));
  AOI211_X1 g384(.A(KEYINPUT66), .B(new_n585_), .C1(new_n574_), .C2(new_n575_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n579_), .B1(new_n584_), .B2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n565_), .A2(new_n570_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n582_), .B1(new_n589_), .B2(new_n581_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n537_), .B1(new_n588_), .B2(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n589_), .B1(new_n577_), .B2(new_n571_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n592_), .B(new_n573_), .C1(new_n583_), .C2(new_n586_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n590_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n593_), .A2(new_n594_), .A3(new_n536_), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n591_), .A2(KEYINPUT13), .A3(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(KEYINPUT13), .B1(new_n591_), .B2(new_n595_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n531_), .A2(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n474_), .A2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n521_), .A2(new_n565_), .A3(new_n522_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G232gat), .A2(G233gat), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n603_), .B(KEYINPUT67), .Z(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT34), .ZN(new_n605_));
  OAI21_X1  g404(.A(KEYINPUT70), .B1(new_n605_), .B2(KEYINPUT35), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n606_), .B1(new_n486_), .B2(new_n574_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n602_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n605_), .A2(KEYINPUT35), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G190gat), .B(G218gat), .ZN(new_n612_));
  INV_X1    g411(.A(G134gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT69), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n615_), .A2(G162gat), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT36), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(G162gat), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n616_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n602_), .A2(new_n609_), .A3(new_n607_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n611_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT71), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n611_), .A2(KEYINPUT71), .A3(new_n620_), .A4(new_n621_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n621_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n609_), .B1(new_n602_), .B2(new_n607_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n617_), .B1(new_n616_), .B2(new_n618_), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT72), .B1(new_n620_), .B2(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n615_), .B(G162gat), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT36), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT72), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n633_), .A2(new_n634_), .A3(new_n619_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n631_), .A2(new_n635_), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n629_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n626_), .A2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n638_), .A2(KEYINPUT73), .A3(KEYINPUT37), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT73), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n636_), .B1(new_n611_), .B2(new_n621_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n641_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT37), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n640_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  OAI211_X1 g443(.A(new_n619_), .B(new_n633_), .C1(new_n627_), .C2(new_n628_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n626_), .A2(new_n643_), .A3(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n639_), .A2(new_n644_), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(G127gat), .B(G155gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT16), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(G183gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(G211gat), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT17), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n499_), .B1(G231gat), .B2(G233gat), .ZN(new_n655_));
  NAND2_X1  g454(.A1(G231gat), .A2(G233gat), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n656_), .B1(new_n494_), .B2(new_n498_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n575_), .B1(new_n655_), .B2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n500_), .A2(new_n656_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n657_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n659_), .A2(new_n570_), .A3(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT17), .B1(new_n658_), .B2(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n654_), .B1(new_n662_), .B2(new_n652_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n658_), .A2(new_n661_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT75), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n663_), .A2(new_n666_), .ZN(new_n667_));
  OAI211_X1 g466(.A(new_n665_), .B(new_n654_), .C1(new_n662_), .C2(new_n652_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n648_), .A2(new_n670_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n601_), .A2(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n672_), .A2(new_n495_), .A3(new_n432_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT38), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n444_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT97), .ZN(new_n677_));
  OAI211_X1 g476(.A(new_n301_), .B(new_n299_), .C1(new_n453_), .C2(KEYINPUT33), .ZN(new_n678_));
  INV_X1    g477(.A(new_n455_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n451_), .B1(new_n431_), .B2(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n467_), .B1(new_n678_), .B2(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n469_), .B1(new_n681_), .B2(new_n448_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n313_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n403_), .B1(new_n433_), .B2(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n677_), .B1(new_n682_), .B2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n472_), .A2(KEYINPUT97), .A3(new_n450_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n676_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n626_), .A2(new_n645_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT100), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n687_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n600_), .A2(new_n669_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT99), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G1gat), .B1(new_n694_), .B2(new_n433_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n673_), .A2(new_n674_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n675_), .A2(new_n695_), .A3(new_n696_), .ZN(G1324gat));
  INV_X1    g496(.A(new_n490_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n317_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n672_), .A2(new_n698_), .A3(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n691_), .A2(new_n699_), .A3(new_n693_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT39), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n701_), .A2(new_n702_), .A3(G8gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n701_), .B2(G8gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n700_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT101), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT101), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n700_), .B(new_n707_), .C1(new_n703_), .C2(new_n704_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n706_), .A2(KEYINPUT40), .A3(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT40), .B1(new_n706_), .B2(new_n708_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1325gat));
  OAI21_X1  g510(.A(G15gat), .B1(new_n694_), .B2(new_n469_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT102), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n712_), .A2(KEYINPUT102), .ZN(new_n715_));
  OAI21_X1  g514(.A(KEYINPUT103), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n712_), .A2(KEYINPUT102), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT103), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n717_), .A2(new_n718_), .A3(new_n713_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n716_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT41), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(G15gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n672_), .A2(new_n723_), .A3(new_n443_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n716_), .A2(new_n719_), .A3(KEYINPUT41), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n722_), .A2(new_n724_), .A3(new_n725_), .ZN(G1326gat));
  OAI21_X1  g525(.A(G22gat), .B1(new_n694_), .B2(new_n403_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT42), .ZN(new_n728_));
  INV_X1    g527(.A(G22gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n672_), .A2(new_n729_), .A3(new_n448_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(G1327gat));
  OAI21_X1  g530(.A(KEYINPUT43), .B1(new_n687_), .B2(new_n647_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n474_), .A2(new_n733_), .A3(new_n648_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n600_), .A2(new_n670_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT44), .B1(new_n735_), .B2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT44), .ZN(new_n739_));
  AOI211_X1 g538(.A(new_n739_), .B(new_n736_), .C1(new_n732_), .C2(new_n734_), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n738_), .A2(new_n740_), .A3(new_n433_), .ZN(new_n741_));
  INV_X1    g540(.A(G29gat), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n669_), .A2(new_n688_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT104), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n601_), .A2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n432_), .A2(new_n742_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT105), .ZN(new_n747_));
  OAI22_X1  g546(.A1(new_n741_), .A2(new_n742_), .B1(new_n745_), .B2(new_n747_), .ZN(G1328gat));
  INV_X1    g547(.A(KEYINPUT46), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT106), .ZN(new_n750_));
  OR2_X1    g549(.A1(new_n749_), .A2(KEYINPUT106), .ZN(new_n751_));
  INV_X1    g550(.A(G36gat), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n738_), .A2(new_n740_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n753_), .B2(new_n699_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n601_), .A2(new_n744_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n755_), .A2(KEYINPUT45), .A3(new_n752_), .A4(new_n699_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n699_), .A2(new_n752_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n745_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n756_), .A2(new_n759_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n750_), .B(new_n751_), .C1(new_n754_), .C2(new_n760_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n687_), .A2(KEYINPUT43), .A3(new_n647_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n733_), .B1(new_n474_), .B2(new_n648_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n737_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n739_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n735_), .A2(KEYINPUT44), .A3(new_n737_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n765_), .A2(new_n699_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(G36gat), .ZN(new_n768_));
  INV_X1    g567(.A(new_n760_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n768_), .A2(new_n769_), .A3(KEYINPUT106), .A4(new_n749_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n761_), .A2(new_n770_), .ZN(G1329gat));
  INV_X1    g570(.A(G43gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n772_), .B1(new_n745_), .B2(new_n469_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT108), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n469_), .A2(new_n772_), .ZN(new_n775_));
  AOI21_X1  g574(.A(KEYINPUT107), .B1(new_n753_), .B2(new_n775_), .ZN(new_n776_));
  AND4_X1   g575(.A1(KEYINPUT107), .A2(new_n765_), .A3(new_n766_), .A4(new_n775_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n774_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT47), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT47), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n780_), .B(new_n774_), .C1(new_n776_), .C2(new_n777_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1330gat));
  AOI21_X1  g581(.A(G50gat), .B1(new_n755_), .B2(new_n448_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n403_), .A2(new_n481_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n753_), .B2(new_n784_), .ZN(G1331gat));
  INV_X1    g584(.A(new_n510_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n516_), .A2(new_n517_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n476_), .B1(new_n787_), .B2(new_n527_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n514_), .B1(new_n786_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(new_n525_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n790_), .A2(new_n598_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n687_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n671_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n794_), .A2(KEYINPUT109), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n432_), .B1(new_n794_), .B2(KEYINPUT109), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n406_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n792_), .A2(new_n670_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n691_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n432_), .A2(G57gat), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n797_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT110), .ZN(G1332gat));
  OAI21_X1  g601(.A(G64gat), .B1(new_n799_), .B2(new_n317_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(KEYINPUT48), .ZN(new_n804_));
  OR2_X1    g603(.A1(new_n317_), .A2(G64gat), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n794_), .B2(new_n805_), .ZN(G1333gat));
  OR3_X1    g605(.A1(new_n794_), .A2(G71gat), .A3(new_n469_), .ZN(new_n807_));
  OAI21_X1  g606(.A(G71gat), .B1(new_n799_), .B2(new_n469_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n808_), .A2(KEYINPUT49), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n808_), .A2(KEYINPUT49), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n807_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(KEYINPUT111), .ZN(G1334gat));
  OAI21_X1  g611(.A(G78gat), .B1(new_n799_), .B2(new_n403_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT50), .ZN(new_n814_));
  OR2_X1    g613(.A1(new_n403_), .A2(G78gat), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n814_), .B1(new_n794_), .B2(new_n815_), .ZN(G1335gat));
  AND2_X1   g615(.A1(new_n793_), .A2(new_n744_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n817_), .A2(new_n408_), .A3(new_n432_), .ZN(new_n818_));
  AOI211_X1 g617(.A(new_n669_), .B(new_n792_), .C1(new_n732_), .C2(new_n734_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n819_), .A2(new_n432_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n818_), .B1(new_n820_), .B2(new_n408_), .ZN(G1336gat));
  NAND3_X1  g620(.A1(new_n817_), .A2(new_n561_), .A3(new_n699_), .ZN(new_n822_));
  AND2_X1   g621(.A1(new_n819_), .A2(new_n699_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n823_), .B2(new_n561_), .ZN(G1337gat));
  AND3_X1   g623(.A1(new_n817_), .A2(new_n557_), .A3(new_n443_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n819_), .A2(new_n443_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(G99gat), .ZN(new_n827_));
  XOR2_X1   g626(.A(new_n827_), .B(KEYINPUT51), .Z(G1338gat));
  NAND4_X1  g627(.A1(new_n735_), .A2(new_n670_), .A3(new_n448_), .A4(new_n791_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT113), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n830_), .A3(G106gat), .ZN(new_n831_));
  XNOR2_X1  g630(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n830_), .B1(new_n829_), .B2(G106gat), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n829_), .A2(new_n830_), .A3(G106gat), .A4(new_n832_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n817_), .A2(new_n558_), .A3(new_n448_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(KEYINPUT53), .B1(new_n836_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n839_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n841_), .B(new_n842_), .C1(new_n835_), .C2(new_n834_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n840_), .A2(new_n843_), .ZN(G1339gat));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n789_), .A2(new_n667_), .A3(new_n668_), .A4(new_n525_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(new_n599_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n531_), .A2(new_n669_), .A3(KEYINPUT114), .A4(new_n598_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n849_), .A2(new_n850_), .A3(new_n647_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n850_), .B1(new_n849_), .B2(new_n647_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n514_), .B1(new_n524_), .B2(new_n476_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n787_), .A2(new_n502_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n475_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n789_), .A2(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n859_), .B1(new_n591_), .B2(new_n595_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT55), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n592_), .A2(new_n581_), .A3(new_n573_), .ZN(new_n862_));
  AOI22_X1  g661(.A1(new_n593_), .A2(new_n861_), .B1(new_n862_), .B2(new_n585_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n588_), .A2(KEYINPUT55), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n536_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT115), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT56), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n870_));
  OAI21_X1  g669(.A(KEYINPUT116), .B1(new_n868_), .B2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n862_), .A2(new_n585_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n872_), .B1(new_n588_), .B2(KEYINPUT55), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n593_), .A2(new_n861_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n537_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT115), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n876_), .A2(new_n877_), .A3(new_n867_), .A4(new_n869_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n865_), .A2(KEYINPUT56), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n871_), .A2(new_n878_), .A3(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n790_), .A2(new_n595_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n860_), .B1(new_n880_), .B2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n688_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n854_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n789_), .A2(new_n858_), .A3(new_n595_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n875_), .A2(new_n869_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n879_), .ZN(new_n888_));
  AOI21_X1  g687(.A(KEYINPUT58), .B1(new_n886_), .B2(new_n888_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n889_), .A2(new_n647_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n888_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n789_), .A2(new_n858_), .A3(new_n595_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(KEYINPUT117), .B1(new_n893_), .B2(KEYINPUT58), .ZN(new_n894_));
  AND4_X1   g693(.A1(KEYINPUT117), .A2(new_n886_), .A3(KEYINPUT58), .A4(new_n888_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n890_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n879_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n876_), .A2(new_n869_), .A3(new_n867_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n897_), .B1(new_n898_), .B2(KEYINPUT116), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n881_), .B1(new_n899_), .B2(new_n878_), .ZN(new_n900_));
  OAI211_X1 g699(.A(KEYINPUT57), .B(new_n688_), .C1(new_n900_), .C2(new_n860_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n885_), .A2(new_n896_), .A3(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n853_), .B1(new_n902_), .B2(new_n670_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n699_), .A2(new_n433_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n443_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n903_), .A2(new_n448_), .A3(new_n905_), .ZN(new_n906_));
  INV_X1    g705(.A(G113gat), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n906_), .A2(new_n907_), .A3(new_n790_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT59), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n906_), .A2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n906_), .A2(new_n909_), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n911_), .A2(new_n912_), .A3(new_n531_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n908_), .B1(new_n913_), .B2(new_n907_), .ZN(G1340gat));
  INV_X1    g713(.A(KEYINPUT60), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n915_), .B1(new_n598_), .B2(G120gat), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n598_), .B1(new_n906_), .B2(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n902_), .A2(new_n670_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n853_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  NAND4_X1  g719(.A1(new_n920_), .A2(new_n403_), .A3(new_n443_), .A4(new_n904_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(KEYINPUT59), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n917_), .A2(new_n922_), .A3(new_n910_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(G120gat), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n906_), .A2(new_n915_), .A3(new_n916_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(G1341gat));
  AOI21_X1  g725(.A(G127gat), .B1(new_n906_), .B2(new_n669_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n911_), .A2(new_n912_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n669_), .A2(G127gat), .ZN(new_n929_));
  XOR2_X1   g728(.A(new_n929_), .B(KEYINPUT118), .Z(new_n930_));
  AOI21_X1  g729(.A(new_n927_), .B1(new_n928_), .B2(new_n930_), .ZN(G1342gat));
  AOI21_X1  g730(.A(G134gat), .B1(new_n906_), .B2(new_n690_), .ZN(new_n932_));
  XOR2_X1   g731(.A(KEYINPUT119), .B(G134gat), .Z(new_n933_));
  NOR2_X1   g732(.A1(new_n647_), .A2(new_n933_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n932_), .B1(new_n928_), .B2(new_n934_), .ZN(G1343gat));
  NOR2_X1   g734(.A1(new_n903_), .A2(new_n443_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT120), .ZN(new_n937_));
  NOR3_X1   g736(.A1(new_n699_), .A2(new_n403_), .A3(new_n433_), .ZN(new_n938_));
  AND3_X1   g737(.A1(new_n936_), .A2(new_n937_), .A3(new_n938_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n937_), .B1(new_n936_), .B2(new_n938_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n790_), .B1(new_n939_), .B2(new_n940_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(KEYINPUT121), .B(G141gat), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n941_), .A2(new_n942_), .ZN(new_n943_));
  INV_X1    g742(.A(new_n942_), .ZN(new_n944_));
  OAI211_X1 g743(.A(new_n790_), .B(new_n944_), .C1(new_n939_), .C2(new_n940_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n943_), .A2(new_n945_), .ZN(G1344gat));
  OAI21_X1  g745(.A(new_n599_), .B1(new_n939_), .B2(new_n940_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(G148gat), .ZN(new_n948_));
  OAI211_X1 g747(.A(new_n323_), .B(new_n599_), .C1(new_n939_), .C2(new_n940_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n948_), .A2(new_n949_), .ZN(G1345gat));
  OAI21_X1  g749(.A(new_n669_), .B1(new_n939_), .B2(new_n940_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(KEYINPUT61), .B(G155gat), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n951_), .A2(new_n952_), .ZN(new_n953_));
  INV_X1    g752(.A(new_n952_), .ZN(new_n954_));
  OAI211_X1 g753(.A(new_n669_), .B(new_n954_), .C1(new_n939_), .C2(new_n940_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n953_), .A2(new_n955_), .ZN(G1346gat));
  INV_X1    g755(.A(new_n940_), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n936_), .A2(new_n937_), .A3(new_n938_), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n647_), .B1(new_n957_), .B2(new_n958_), .ZN(new_n959_));
  INV_X1    g758(.A(G162gat), .ZN(new_n960_));
  NOR2_X1   g759(.A1(new_n939_), .A2(new_n940_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n690_), .A2(new_n960_), .ZN(new_n962_));
  OAI22_X1  g761(.A1(new_n959_), .A2(new_n960_), .B1(new_n961_), .B2(new_n962_), .ZN(G1347gat));
  AOI21_X1  g762(.A(new_n236_), .B1(KEYINPUT123), .B2(KEYINPUT62), .ZN(new_n964_));
  NAND3_X1  g763(.A1(new_n699_), .A2(new_n433_), .A3(new_n443_), .ZN(new_n965_));
  XNOR2_X1  g764(.A(new_n965_), .B(KEYINPUT122), .ZN(new_n966_));
  INV_X1    g765(.A(new_n966_), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n920_), .A2(new_n403_), .A3(new_n967_), .ZN(new_n968_));
  OAI21_X1  g767(.A(new_n964_), .B1(new_n968_), .B2(new_n531_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n970_));
  OR2_X1    g769(.A1(new_n969_), .A2(new_n970_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n969_), .A2(new_n970_), .ZN(new_n972_));
  INV_X1    g771(.A(KEYINPUT124), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n968_), .A2(new_n973_), .ZN(new_n974_));
  NOR3_X1   g773(.A1(new_n903_), .A2(new_n448_), .A3(new_n966_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n975_), .A2(KEYINPUT124), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n974_), .A2(new_n976_), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n790_), .A2(new_n245_), .ZN(new_n978_));
  OAI211_X1 g777(.A(new_n971_), .B(new_n972_), .C1(new_n977_), .C2(new_n978_), .ZN(G1348gat));
  NOR3_X1   g778(.A1(new_n968_), .A2(new_n237_), .A3(new_n598_), .ZN(new_n980_));
  NAND3_X1  g779(.A1(new_n974_), .A2(new_n976_), .A3(new_n599_), .ZN(new_n981_));
  AOI21_X1  g780(.A(new_n980_), .B1(new_n981_), .B2(new_n237_), .ZN(G1349gat));
  AOI21_X1  g781(.A(new_n448_), .B1(new_n918_), .B2(new_n919_), .ZN(new_n983_));
  AOI21_X1  g782(.A(KEYINPUT124), .B1(new_n983_), .B2(new_n967_), .ZN(new_n984_));
  NOR4_X1   g783(.A1(new_n903_), .A2(new_n973_), .A3(new_n448_), .A4(new_n966_), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n228_), .A2(new_n230_), .ZN(new_n986_));
  NAND2_X1  g785(.A1(new_n669_), .A2(new_n986_), .ZN(new_n987_));
  NOR3_X1   g786(.A1(new_n984_), .A2(new_n985_), .A3(new_n987_), .ZN(new_n988_));
  AOI21_X1  g787(.A(G183gat), .B1(new_n975_), .B2(new_n669_), .ZN(new_n989_));
  OAI21_X1  g788(.A(KEYINPUT125), .B1(new_n988_), .B2(new_n989_), .ZN(new_n990_));
  INV_X1    g789(.A(KEYINPUT125), .ZN(new_n991_));
  OAI21_X1  g790(.A(new_n227_), .B1(new_n968_), .B2(new_n670_), .ZN(new_n992_));
  OAI211_X1 g791(.A(new_n991_), .B(new_n992_), .C1(new_n977_), .C2(new_n987_), .ZN(new_n993_));
  NAND2_X1  g792(.A1(new_n990_), .A2(new_n993_), .ZN(G1350gat));
  OAI21_X1  g793(.A(G190gat), .B1(new_n977_), .B2(new_n647_), .ZN(new_n995_));
  NAND3_X1  g794(.A1(new_n690_), .A2(new_n232_), .A3(new_n234_), .ZN(new_n996_));
  OAI21_X1  g795(.A(new_n995_), .B1(new_n977_), .B2(new_n996_), .ZN(G1351gat));
  NOR3_X1   g796(.A1(new_n317_), .A2(new_n403_), .A3(new_n432_), .ZN(new_n998_));
  NAND2_X1  g797(.A1(new_n936_), .A2(new_n998_), .ZN(new_n999_));
  NOR2_X1   g798(.A1(new_n999_), .A2(new_n531_), .ZN(new_n1000_));
  XOR2_X1   g799(.A(new_n1000_), .B(G197gat), .Z(G1352gat));
  NOR2_X1   g800(.A1(new_n999_), .A2(new_n598_), .ZN(new_n1002_));
  XNOR2_X1  g801(.A(new_n1002_), .B(new_n533_), .ZN(G1353gat));
  NAND3_X1  g802(.A1(new_n936_), .A2(new_n669_), .A3(new_n998_), .ZN(new_n1004_));
  XNOR2_X1  g803(.A(KEYINPUT63), .B(G211gat), .ZN(new_n1005_));
  NOR2_X1   g804(.A1(new_n1004_), .A2(new_n1005_), .ZN(new_n1006_));
  NOR2_X1   g805(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1007_));
  AOI21_X1  g806(.A(new_n1006_), .B1(new_n1004_), .B2(new_n1007_), .ZN(G1354gat));
  AND3_X1   g807(.A1(new_n936_), .A2(new_n690_), .A3(new_n998_), .ZN(new_n1009_));
  XNOR2_X1  g808(.A(KEYINPUT126), .B(G218gat), .ZN(new_n1010_));
  INV_X1    g809(.A(new_n1010_), .ZN(new_n1011_));
  NAND2_X1  g810(.A1(new_n648_), .A2(new_n1011_), .ZN(new_n1012_));
  OAI22_X1  g811(.A1(new_n1009_), .A2(new_n1011_), .B1(new_n999_), .B2(new_n1012_), .ZN(new_n1013_));
  NAND2_X1  g812(.A1(new_n1013_), .A2(KEYINPUT127), .ZN(new_n1014_));
  INV_X1    g813(.A(KEYINPUT127), .ZN(new_n1015_));
  OAI221_X1 g814(.A(new_n1015_), .B1(new_n999_), .B2(new_n1012_), .C1(new_n1009_), .C2(new_n1011_), .ZN(new_n1016_));
  NAND2_X1  g815(.A1(new_n1014_), .A2(new_n1016_), .ZN(G1355gat));
endmodule


