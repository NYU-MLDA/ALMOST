//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 0 1 0 1 0 0 0 0 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 0 1 0 0 1 1 1 0 1 1 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n765_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n927_, new_n929_, new_n930_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n947_, new_n948_, new_n949_;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(new_n202_), .A2(KEYINPUT21), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(KEYINPUT21), .ZN(new_n204_));
  XOR2_X1   g003(.A(G197gat), .B(G204gat), .Z(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n204_), .A2(new_n205_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT82), .ZN(new_n210_));
  INV_X1    g009(.A(G141gat), .ZN(new_n211_));
  INV_X1    g010(.A(G148gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(KEYINPUT83), .A3(KEYINPUT3), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G141gat), .A2(G148gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT2), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT2), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(G141gat), .A3(G148gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  NOR3_X1   g018(.A1(KEYINPUT82), .A2(G141gat), .A3(G148gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT83), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G141gat), .A2(G148gat), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n223_), .B1(new_n224_), .B2(new_n221_), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n214_), .B(new_n219_), .C1(new_n222_), .C2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT84), .ZN(new_n227_));
  NOR3_X1   g026(.A1(KEYINPUT83), .A2(G141gat), .A3(G148gat), .ZN(new_n228_));
  OAI22_X1  g027(.A1(new_n221_), .A2(new_n220_), .B1(new_n228_), .B2(new_n223_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT84), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n229_), .A2(new_n230_), .A3(new_n214_), .A4(new_n219_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n227_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(G155gat), .ZN(new_n233_));
  INV_X1    g032(.A(G162gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(G155gat), .A2(G162gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT81), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n232_), .A2(new_n236_), .A3(new_n238_), .ZN(new_n239_));
  OR2_X1    g038(.A1(new_n236_), .A2(KEYINPUT1), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n236_), .A2(KEYINPUT1), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n240_), .A2(new_n238_), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n224_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n242_), .A2(new_n243_), .A3(new_n215_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n239_), .A2(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n209_), .B1(new_n245_), .B2(KEYINPUT29), .ZN(new_n246_));
  XOR2_X1   g045(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  OR2_X1    g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n248_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n245_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT29), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G78gat), .B(G106gat), .ZN(new_n254_));
  XOR2_X1   g053(.A(new_n254_), .B(KEYINPUT86), .Z(new_n255_));
  NAND3_X1  g054(.A1(new_n252_), .A2(new_n253_), .A3(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n255_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n257_), .B1(new_n245_), .B2(KEYINPUT29), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G22gat), .B(G50gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G228gat), .A2(G233gat), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n259_), .B(new_n260_), .Z(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n256_), .A2(new_n258_), .A3(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n262_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n251_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n258_), .ZN(new_n267_));
  NOR3_X1   g066(.A1(new_n245_), .A2(KEYINPUT29), .A3(new_n257_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n261_), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n269_), .A2(new_n249_), .A3(new_n250_), .A4(new_n263_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n266_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G15gat), .B(G43gat), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G227gat), .A2(G233gat), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G169gat), .A2(G176gat), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G183gat), .A2(G190gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT23), .ZN(new_n280_));
  OR2_X1    g079(.A1(G183gat), .A2(G190gat), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n278_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(G176gat), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT22), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT78), .B1(new_n284_), .B2(G169gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT22), .B(G169gat), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n283_), .B(new_n285_), .C1(new_n286_), .C2(KEYINPUT78), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n282_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT30), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT25), .B(G183gat), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT77), .ZN(new_n291_));
  INV_X1    g090(.A(G190gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT26), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n292_), .A2(KEYINPUT26), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n290_), .B(new_n293_), .C1(new_n294_), .C2(new_n291_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(G169gat), .A2(G176gat), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n297_), .A2(KEYINPUT24), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n297_), .A2(KEYINPUT24), .A3(new_n277_), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n295_), .A2(new_n280_), .A3(new_n298_), .A4(new_n299_), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n288_), .A2(new_n289_), .A3(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n289_), .B1(new_n288_), .B2(new_n300_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n276_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n288_), .A2(new_n300_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT30), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n288_), .A2(new_n289_), .A3(new_n300_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n305_), .A2(new_n306_), .A3(new_n275_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G71gat), .B(G99gat), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n303_), .A2(new_n307_), .A3(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n309_), .B1(new_n303_), .B2(new_n307_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n274_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n303_), .A2(new_n307_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n308_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n303_), .A2(new_n307_), .A3(new_n309_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(new_n273_), .A3(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n312_), .A2(new_n316_), .A3(KEYINPUT80), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G127gat), .B(G134gat), .ZN(new_n318_));
  INV_X1    g117(.A(G113gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(G120gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n317_), .A2(new_n325_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n312_), .A2(new_n316_), .A3(KEYINPUT80), .A4(new_n324_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n272_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT0), .B(G57gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(G85gat), .ZN(new_n332_));
  XOR2_X1   g131(.A(G1gat), .B(G29gat), .Z(new_n333_));
  XOR2_X1   g132(.A(new_n332_), .B(new_n333_), .Z(new_n334_));
  XNOR2_X1  g133(.A(new_n320_), .B(G120gat), .ZN(new_n335_));
  INV_X1    g134(.A(new_n238_), .ZN(new_n336_));
  AOI211_X1 g135(.A(new_n235_), .B(new_n336_), .C1(new_n227_), .C2(new_n231_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n244_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n335_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT91), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n239_), .A2(new_n322_), .A3(new_n244_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n245_), .A2(KEYINPUT91), .A3(new_n335_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT4), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT92), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT4), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n245_), .A2(new_n347_), .A3(new_n335_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G225gat), .A2(G233gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n345_), .A2(new_n346_), .A3(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n347_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT92), .B1(new_n354_), .B2(new_n351_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT93), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n357_), .B1(new_n344_), .B2(new_n349_), .ZN(new_n358_));
  AOI211_X1 g157(.A(KEYINPUT93), .B(new_n350_), .C1(new_n342_), .C2(new_n343_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n334_), .B1(new_n356_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n344_), .A2(new_n349_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT93), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n344_), .A2(new_n357_), .A3(new_n349_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n334_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n365_), .A2(new_n366_), .A3(new_n353_), .A4(new_n355_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n361_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G226gat), .A2(G233gat), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n369_), .B(KEYINPUT19), .Z(new_n370_));
  NAND2_X1  g169(.A1(new_n286_), .A2(new_n283_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n282_), .A2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT26), .B(G190gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n290_), .A2(new_n373_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n298_), .A2(new_n374_), .A3(new_n280_), .A4(new_n299_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n209_), .A2(new_n372_), .A3(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(KEYINPUT96), .B1(new_n376_), .B2(KEYINPUT20), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n377_), .B1(new_n304_), .B2(new_n208_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n376_), .A2(KEYINPUT96), .A3(KEYINPUT20), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n370_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT20), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n288_), .A2(new_n300_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n381_), .B1(new_n382_), .B2(new_n209_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n372_), .A2(new_n375_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n208_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT88), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n384_), .A2(KEYINPUT88), .A3(new_n208_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n383_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n370_), .B(KEYINPUT87), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n380_), .A2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT18), .B(G64gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(G92gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G8gat), .B(G36gat), .ZN(new_n395_));
  XOR2_X1   g194(.A(new_n394_), .B(new_n395_), .Z(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT32), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n392_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT89), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n389_), .A2(new_n400_), .A3(new_n390_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n400_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT95), .ZN(new_n405_));
  OR2_X1    g204(.A1(new_n376_), .A2(KEYINPUT90), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n381_), .B1(new_n376_), .B2(KEYINPUT90), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n304_), .A2(new_n208_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n406_), .A2(new_n407_), .A3(new_n370_), .A4(new_n408_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n404_), .A2(new_n405_), .A3(new_n409_), .A4(new_n397_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n389_), .A2(new_n390_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT89), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n412_), .A2(new_n401_), .A3(new_n409_), .A4(new_n397_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT95), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n368_), .A2(new_n399_), .A3(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT33), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n367_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n412_), .A2(new_n401_), .A3(new_n409_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n396_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n412_), .A2(new_n396_), .A3(new_n401_), .A4(new_n409_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n345_), .A2(new_n349_), .A3(new_n348_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n344_), .A2(new_n350_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n425_), .A2(KEYINPUT94), .A3(new_n334_), .A4(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT94), .ZN(new_n428_));
  INV_X1    g227(.A(new_n348_), .ZN(new_n429_));
  NOR3_X1   g228(.A1(new_n354_), .A2(new_n350_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n426_), .A2(new_n334_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n428_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n424_), .B1(new_n427_), .B2(new_n432_), .ZN(new_n433_));
  AND2_X1   g232(.A1(new_n353_), .A2(new_n355_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n434_), .A2(KEYINPUT33), .A3(new_n366_), .A4(new_n365_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n419_), .A2(new_n433_), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n330_), .B1(new_n417_), .B2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n328_), .A2(new_n271_), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n326_), .A2(new_n327_), .B1(new_n266_), .B2(new_n270_), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n361_), .B(new_n367_), .C1(new_n438_), .C2(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n421_), .B1(new_n380_), .B2(new_n391_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n441_), .A2(KEYINPUT27), .A3(new_n423_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT27), .ZN(new_n443_));
  AOI21_X1  g242(.A(KEYINPUT97), .B1(new_n424_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT97), .ZN(new_n445_));
  AOI211_X1 g244(.A(new_n445_), .B(KEYINPUT27), .C1(new_n422_), .C2(new_n423_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n442_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n440_), .A2(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n437_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT74), .ZN(new_n450_));
  XNOR2_X1  g249(.A(KEYINPUT16), .B(G183gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(G211gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G127gat), .B(G155gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n450_), .B1(new_n454_), .B2(KEYINPUT17), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G231gat), .A2(G233gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G15gat), .B(G22gat), .ZN(new_n458_));
  XOR2_X1   g257(.A(KEYINPUT72), .B(G1gat), .Z(new_n459_));
  INV_X1    g258(.A(KEYINPUT14), .ZN(new_n460_));
  OAI211_X1 g259(.A(G8gat), .B(new_n458_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n458_), .A2(new_n460_), .ZN(new_n462_));
  INV_X1    g261(.A(G8gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n461_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT73), .B(G1gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n461_), .A2(new_n466_), .A3(new_n464_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n457_), .B(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G57gat), .B(G64gat), .ZN(new_n473_));
  OR2_X1    g272(.A1(new_n473_), .A2(KEYINPUT11), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(KEYINPUT11), .ZN(new_n475_));
  XOR2_X1   g274(.A(G71gat), .B(G78gat), .Z(new_n476_));
  NAND3_X1  g275(.A1(new_n474_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n475_), .A2(new_n476_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n472_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n454_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT17), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n472_), .A2(new_n480_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n481_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n449_), .A2(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G113gat), .B(G141gat), .Z(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(G169gat), .ZN(new_n490_));
  INV_X1    g289(.A(G197gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G229gat), .A2(G233gat), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT75), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G29gat), .B(G36gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(G43gat), .ZN(new_n496_));
  INV_X1    g295(.A(G50gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n495_), .A2(G43gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n495_), .A2(G43gat), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n499_), .A2(G50gat), .A3(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n498_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n502_), .A2(new_n469_), .A3(new_n468_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n502_), .B1(new_n469_), .B2(new_n468_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n494_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n498_), .A2(new_n501_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n470_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n508_), .A2(KEYINPUT75), .A3(new_n503_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n493_), .B1(new_n506_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n493_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT15), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n502_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n498_), .A2(KEYINPUT15), .A3(new_n501_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  AOI211_X1 g314(.A(new_n511_), .B(new_n505_), .C1(new_n515_), .C2(new_n471_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n492_), .B1(new_n510_), .B2(new_n516_), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n508_), .A2(KEYINPUT75), .A3(new_n503_), .ZN(new_n518_));
  AOI21_X1  g317(.A(KEYINPUT75), .B1(new_n508_), .B2(new_n503_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n511_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n505_), .B1(new_n515_), .B2(new_n471_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(new_n493_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n492_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n520_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n517_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT76), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT70), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT35), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G232gat), .A2(G233gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT34), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT6), .ZN(new_n533_));
  INV_X1    g332(.A(G99gat), .ZN(new_n534_));
  INV_X1    g333(.A(G106gat), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n533_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT9), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n539_), .A2(G85gat), .A3(G92gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G85gat), .B(G92gat), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n538_), .B(new_n540_), .C1(new_n539_), .C2(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(KEYINPUT10), .B(G99gat), .Z(new_n543_));
  AND2_X1   g342(.A1(new_n543_), .A2(new_n535_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n534_), .A2(new_n535_), .A3(KEYINPUT64), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT64), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n547_), .B1(G99gat), .B2(G106gat), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT7), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n546_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT65), .ZN(new_n551_));
  OAI21_X1  g350(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n536_), .A2(new_n537_), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT65), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n546_), .A2(new_n548_), .A3(new_n554_), .A4(new_n549_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n551_), .A2(new_n553_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT8), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n541_), .A2(KEYINPUT66), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n556_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n557_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n507_), .B(new_n545_), .C1(new_n559_), .C2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT68), .ZN(new_n562_));
  AOI211_X1 g361(.A(new_n529_), .B(new_n532_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n545_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT67), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT67), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n566_), .B(new_n545_), .C1(new_n559_), .C2(new_n560_), .ZN(new_n567_));
  AOI22_X1  g366(.A1(new_n565_), .A2(new_n567_), .B1(new_n514_), .B2(new_n513_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n532_), .A2(new_n529_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n561_), .A2(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n563_), .B1(new_n568_), .B2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n542_), .A2(new_n544_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n556_), .A2(new_n558_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT8), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n556_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n572_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n576_), .A2(new_n566_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n567_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n515_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n561_), .A2(new_n562_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n580_), .A2(KEYINPUT35), .A3(new_n531_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n570_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n579_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n571_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT71), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G190gat), .B(G218gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(G134gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(new_n234_), .ZN(new_n588_));
  XOR2_X1   g387(.A(new_n588_), .B(KEYINPUT36), .Z(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT71), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n571_), .A2(new_n583_), .A3(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n585_), .A2(new_n590_), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT37), .ZN(new_n594_));
  XNOR2_X1  g393(.A(KEYINPUT69), .B(KEYINPUT36), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n583_), .A2(new_n571_), .A3(new_n588_), .A4(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n593_), .A2(new_n594_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n596_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n589_), .B1(new_n571_), .B2(new_n583_), .ZN(new_n599_));
  OAI21_X1  g398(.A(KEYINPUT37), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n528_), .B1(new_n597_), .B2(new_n600_), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n600_), .A2(new_n528_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT12), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n479_), .A2(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n605_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n545_), .B(new_n479_), .C1(new_n559_), .C2(new_n560_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n564_), .A2(new_n480_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n608_), .B1(new_n604_), .B2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G230gat), .A2(G233gat), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n606_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n609_), .A2(new_n607_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n611_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G120gat), .B(G148gat), .ZN(new_n617_));
  INV_X1    g416(.A(G204gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT5), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(new_n283_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n616_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n612_), .A2(new_n615_), .A3(new_n621_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT13), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT13), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n623_), .A2(new_n627_), .A3(new_n624_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n603_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n488_), .A2(new_n527_), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT98), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n459_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n368_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT99), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT99), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n368_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n634_), .A2(new_n635_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT38), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n525_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n626_), .B2(new_n628_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(new_n486_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT100), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n646_), .B(new_n647_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n419_), .A2(new_n433_), .A3(new_n435_), .ZN(new_n649_));
  AOI211_X1 g448(.A(new_n398_), .B(new_n415_), .C1(new_n361_), .C2(new_n367_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n329_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n440_), .A2(new_n447_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n593_), .A2(KEYINPUT101), .A3(new_n596_), .ZN(new_n654_));
  AOI21_X1  g453(.A(KEYINPUT101), .B1(new_n593_), .B2(new_n596_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n648_), .A2(new_n653_), .A3(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G1gat), .B1(new_n657_), .B2(new_n636_), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n634_), .A2(KEYINPUT38), .A3(new_n635_), .A4(new_n640_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n643_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT102), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n643_), .A2(KEYINPUT102), .A3(new_n658_), .A4(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1324gat));
  NAND3_X1  g463(.A1(new_n634_), .A2(new_n463_), .A3(new_n447_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n447_), .ZN(new_n666_));
  OAI21_X1  g465(.A(KEYINPUT103), .B1(new_n657_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n656_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n449_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT103), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n669_), .A2(new_n670_), .A3(new_n447_), .A4(new_n648_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT39), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n667_), .A2(new_n671_), .A3(G8gat), .A4(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n672_), .A2(KEYINPUT39), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n675_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n665_), .A2(new_n676_), .A3(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n678_), .B(new_n679_), .ZN(G1325gat));
  INV_X1    g479(.A(new_n328_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G15gat), .B1(new_n657_), .B2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT41), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n632_), .A2(G15gat), .A3(new_n681_), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1326gat));
  OAI21_X1  g484(.A(G22gat), .B1(new_n657_), .B2(new_n271_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT42), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n632_), .A2(G22gat), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n687_), .B1(new_n271_), .B2(new_n688_), .ZN(G1327gat));
  NOR2_X1   g488(.A1(new_n449_), .A2(new_n656_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(new_n629_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n486_), .A2(new_n526_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G29gat), .B1(new_n695_), .B2(new_n368_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n640_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698_));
  INV_X1    g497(.A(new_n603_), .ZN(new_n699_));
  OAI21_X1  g498(.A(KEYINPUT43), .B1(new_n449_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n701_));
  OAI211_X1 g500(.A(new_n701_), .B(new_n603_), .C1(new_n437_), .C2(new_n448_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n645_), .A2(new_n487_), .ZN(new_n704_));
  AOI211_X1 g503(.A(KEYINPUT106), .B(new_n698_), .C1(new_n703_), .C2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n698_), .A2(KEYINPUT106), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(KEYINPUT44), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n703_), .A2(new_n704_), .A3(new_n707_), .A4(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n697_), .B1(new_n706_), .B2(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n696_), .B1(new_n711_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g511(.A(G36gat), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n692_), .A2(new_n713_), .A3(new_n447_), .A4(new_n693_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT45), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n666_), .B1(new_n706_), .B2(new_n710_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n715_), .B1(new_n716_), .B2(new_n713_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT46), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n715_), .B(KEYINPUT46), .C1(new_n716_), .C2(new_n713_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1329gat));
  NOR3_X1   g520(.A1(new_n694_), .A2(G43gat), .A3(new_n681_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n710_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n328_), .B1(new_n705_), .B2(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n722_), .B1(new_n724_), .B2(G43gat), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g525(.A(new_n272_), .B1(new_n705_), .B2(new_n723_), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n727_), .A2(KEYINPUT107), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(KEYINPUT107), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n728_), .A2(G50gat), .A3(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n695_), .A2(new_n497_), .A3(new_n272_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1331gat));
  AND2_X1   g531(.A1(new_n486_), .A2(new_n526_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n669_), .A2(new_n630_), .A3(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(G57gat), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n734_), .A2(new_n735_), .A3(new_n636_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT110), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n488_), .A2(new_n644_), .A3(new_n630_), .A4(new_n699_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT108), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT109), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(new_n640_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n737_), .B1(new_n741_), .B2(new_n735_), .ZN(G1332gat));
  OAI21_X1  g541(.A(G64gat), .B1(new_n734_), .B2(new_n666_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT48), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n666_), .A2(G64gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n744_), .B1(new_n739_), .B2(new_n745_), .ZN(G1333gat));
  OR3_X1    g545(.A1(new_n739_), .A2(G71gat), .A3(new_n681_), .ZN(new_n747_));
  OAI21_X1  g546(.A(G71gat), .B1(new_n734_), .B2(new_n681_), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n748_), .A2(KEYINPUT111), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(KEYINPUT111), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n749_), .A2(KEYINPUT49), .A3(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(KEYINPUT49), .B1(new_n749_), .B2(new_n750_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n747_), .B1(new_n751_), .B2(new_n752_), .ZN(G1334gat));
  OAI21_X1  g552(.A(G78gat), .B1(new_n734_), .B2(new_n271_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT50), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n271_), .A2(G78gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n755_), .B1(new_n739_), .B2(new_n756_), .ZN(G1335gat));
  NOR3_X1   g556(.A1(new_n629_), .A2(new_n486_), .A3(new_n525_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n690_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(G85gat), .B1(new_n760_), .B2(new_n640_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n703_), .A2(new_n758_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n762_), .A2(new_n636_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n761_), .B1(new_n763_), .B2(G85gat), .ZN(G1336gat));
  INV_X1    g563(.A(G92gat), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n762_), .A2(new_n765_), .A3(new_n666_), .ZN(new_n766_));
  AOI21_X1  g565(.A(G92gat), .B1(new_n760_), .B2(new_n447_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(new_n767_), .ZN(G1337gat));
  OAI21_X1  g567(.A(G99gat), .B1(new_n762_), .B2(new_n681_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n760_), .A2(new_n543_), .A3(new_n328_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n772_), .A2(KEYINPUT112), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n771_), .B(new_n773_), .ZN(G1338gat));
  AOI21_X1  g573(.A(new_n701_), .B1(new_n653_), .B2(new_n603_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n702_), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n272_), .B(new_n758_), .C1(new_n775_), .C2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT113), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n703_), .A2(KEYINPUT113), .A3(new_n272_), .A4(new_n758_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(G106gat), .A3(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT52), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n779_), .A2(new_n783_), .A3(new_n780_), .A4(G106gat), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n760_), .A2(new_n535_), .A3(new_n272_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT53), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT53), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n785_), .A2(new_n789_), .A3(new_n786_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(G1339gat));
  OAI211_X1 g590(.A(new_n733_), .B(new_n629_), .C1(new_n601_), .C2(new_n602_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n792_), .B(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n525_), .A2(new_n624_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT114), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT114), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n525_), .A2(new_n624_), .A3(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT56), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n612_), .A2(KEYINPUT115), .A3(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT115), .B1(new_n612_), .B2(new_n801_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n606_), .A2(new_n610_), .A3(KEYINPUT55), .A4(new_n611_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n604_), .B1(new_n576_), .B2(new_n479_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n607_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n605_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n565_), .B2(new_n567_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n614_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n804_), .A2(new_n809_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n802_), .A2(new_n803_), .A3(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n800_), .B1(new_n811_), .B2(new_n621_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n612_), .A2(new_n801_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT115), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n804_), .A2(new_n809_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n612_), .A2(KEYINPUT115), .A3(new_n801_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n815_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n818_), .A2(KEYINPUT56), .A3(new_n622_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n799_), .B1(new_n812_), .B2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n493_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n521_), .A2(new_n511_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n821_), .A2(new_n492_), .A3(new_n822_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n823_), .A2(new_n524_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n625_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  OAI211_X1 g625(.A(KEYINPUT57), .B(new_n656_), .C1(new_n820_), .C2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT116), .ZN(new_n828_));
  AND3_X1   g627(.A1(new_n818_), .A2(KEYINPUT56), .A3(new_n622_), .ZN(new_n829_));
  AOI21_X1  g628(.A(KEYINPUT56), .B1(new_n818_), .B2(new_n622_), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n624_), .B(new_n824_), .C1(new_n829_), .C2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n812_), .A2(new_n819_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n834_), .A2(KEYINPUT58), .A3(new_n624_), .A4(new_n824_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n833_), .A2(new_n603_), .A3(new_n835_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n796_), .A2(new_n798_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n825_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT116), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n839_), .A2(new_n840_), .A3(KEYINPUT57), .A4(new_n656_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n656_), .B1(new_n820_), .B2(new_n826_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT57), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n828_), .A2(new_n836_), .A3(new_n841_), .A4(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n794_), .B1(new_n845_), .B2(new_n487_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n640_), .A2(new_n666_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n847_), .A2(new_n681_), .A3(new_n272_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n846_), .A2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(G113gat), .B1(new_n850_), .B2(new_n525_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(KEYINPUT117), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT59), .B1(new_n848_), .B2(new_n853_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n828_), .A2(new_n841_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n836_), .A2(new_n844_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n486_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n852_), .B(new_n854_), .C1(new_n857_), .C2(new_n794_), .ZN(new_n858_));
  OAI21_X1  g657(.A(KEYINPUT59), .B1(new_n846_), .B2(new_n849_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n860_), .A2(new_n526_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n851_), .B1(new_n861_), .B2(G113gat), .ZN(G1340gat));
  NAND3_X1  g661(.A1(new_n858_), .A2(new_n630_), .A3(new_n859_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(G120gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n321_), .B1(new_n629_), .B2(KEYINPUT60), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n850_), .B(new_n865_), .C1(KEYINPUT60), .C2(new_n321_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(KEYINPUT118), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT118), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n864_), .A2(new_n869_), .A3(new_n866_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n870_), .ZN(G1341gat));
  INV_X1    g670(.A(G127gat), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n860_), .A2(new_n872_), .A3(new_n487_), .ZN(new_n873_));
  AOI21_X1  g672(.A(G127gat), .B1(new_n850_), .B2(new_n486_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1342gat));
  NOR3_X1   g674(.A1(new_n846_), .A2(new_n656_), .A3(new_n849_), .ZN(new_n876_));
  OR2_X1    g675(.A1(new_n876_), .A2(G134gat), .ZN(new_n877_));
  XOR2_X1   g676(.A(KEYINPUT119), .B(G134gat), .Z(new_n878_));
  NAND2_X1  g677(.A1(new_n603_), .A2(new_n878_), .ZN(new_n879_));
  XOR2_X1   g678(.A(new_n879_), .B(KEYINPUT120), .Z(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n877_), .B1(new_n860_), .B2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT121), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n877_), .B(KEYINPUT121), .C1(new_n860_), .C2(new_n881_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1343gat));
  NAND2_X1  g685(.A1(new_n845_), .A2(new_n487_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n794_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n847_), .A2(new_n328_), .A3(new_n271_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n889_), .A2(new_n890_), .A3(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n891_), .ZN(new_n893_));
  OAI21_X1  g692(.A(KEYINPUT122), .B1(new_n846_), .B2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(new_n525_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n630_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(KEYINPUT123), .B(G148gat), .ZN(new_n899_));
  XOR2_X1   g698(.A(new_n898_), .B(new_n899_), .Z(G1345gat));
  NAND2_X1  g699(.A1(new_n895_), .A2(new_n486_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT61), .B(G155gat), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n901_), .B(new_n902_), .ZN(G1346gat));
  AOI211_X1 g702(.A(new_n234_), .B(new_n699_), .C1(new_n892_), .C2(new_n894_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n656_), .B1(new_n892_), .B2(new_n894_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT124), .ZN(new_n906_));
  OR3_X1    g705(.A1(new_n905_), .A2(new_n906_), .A3(G162gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n905_), .B2(G162gat), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n904_), .B1(new_n907_), .B2(new_n908_), .ZN(G1347gat));
  NAND3_X1  g708(.A1(new_n697_), .A2(new_n328_), .A3(new_n447_), .ZN(new_n910_));
  AND2_X1   g709(.A1(new_n910_), .A2(KEYINPUT125), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n910_), .A2(KEYINPUT125), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n911_), .A2(new_n912_), .A3(new_n272_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n889_), .A2(new_n913_), .ZN(new_n914_));
  OAI21_X1  g713(.A(G169gat), .B1(new_n914_), .B2(new_n644_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(KEYINPUT126), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT126), .ZN(new_n917_));
  OAI211_X1 g716(.A(new_n917_), .B(G169gat), .C1(new_n914_), .C2(new_n644_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n916_), .A2(KEYINPUT62), .A3(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n914_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n920_), .A2(new_n286_), .A3(new_n525_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n915_), .A2(KEYINPUT126), .A3(new_n922_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n919_), .A2(new_n921_), .A3(new_n923_), .ZN(G1348gat));
  NOR2_X1   g723(.A1(new_n914_), .A2(new_n629_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(new_n283_), .ZN(G1349gat));
  NOR2_X1   g725(.A1(new_n914_), .A2(new_n487_), .ZN(new_n927_));
  MUX2_X1   g726(.A(G183gat), .B(new_n290_), .S(new_n927_), .Z(G1350gat));
  OAI21_X1  g727(.A(G190gat), .B1(new_n914_), .B2(new_n699_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n668_), .A2(new_n373_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n914_), .B2(new_n930_), .ZN(G1351gat));
  NOR2_X1   g730(.A1(new_n846_), .A2(new_n368_), .ZN(new_n932_));
  AND2_X1   g731(.A1(new_n447_), .A2(new_n438_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n934_), .A2(new_n644_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(new_n491_), .ZN(G1352gat));
  NOR2_X1   g735(.A1(new_n934_), .A2(new_n629_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(new_n618_), .ZN(G1353gat));
  NOR2_X1   g737(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n939_));
  AND2_X1   g738(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n940_));
  NOR4_X1   g739(.A1(new_n934_), .A2(new_n487_), .A3(new_n939_), .A4(new_n940_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n939_), .B1(new_n934_), .B2(new_n487_), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT127), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(new_n944_));
  OAI211_X1 g743(.A(KEYINPUT127), .B(new_n939_), .C1(new_n934_), .C2(new_n487_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n941_), .B1(new_n944_), .B2(new_n945_), .ZN(G1354gat));
  INV_X1    g745(.A(G218gat), .ZN(new_n947_));
  NOR3_X1   g746(.A1(new_n934_), .A2(new_n947_), .A3(new_n699_), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n932_), .A2(new_n668_), .A3(new_n933_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n948_), .B1(new_n947_), .B2(new_n949_), .ZN(G1355gat));
endmodule


