//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 1 0 0 1 0 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 1 1 1 1 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n824_, new_n825_,
    new_n826_, new_n828_, new_n829_, new_n830_, new_n832_, new_n833_,
    new_n834_, new_n836_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_;
  INV_X1    g000(.A(G183gat), .ZN(new_n202_));
  INV_X1    g001(.A(G190gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT23), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT86), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  OR3_X1    g005(.A1(new_n202_), .A2(new_n203_), .A3(KEYINPUT23), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT24), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n208_), .A2(new_n211_), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n212_), .A2(KEYINPUT87), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(KEYINPUT87), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  OR3_X1    g015(.A1(new_n216_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n202_), .A2(KEYINPUT25), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n218_), .B(KEYINPUT85), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n202_), .A2(KEYINPUT84), .A3(KEYINPUT25), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT26), .B(G190gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n202_), .A2(KEYINPUT25), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT84), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .A4(new_n224_), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n213_), .A2(new_n214_), .A3(new_n217_), .A4(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(G176gat), .ZN(new_n227_));
  INV_X1    g026(.A(G169gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT22), .B1(new_n228_), .B2(KEYINPUT88), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n228_), .A2(KEYINPUT22), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n227_), .B(new_n229_), .C1(new_n230_), .C2(KEYINPUT88), .ZN(new_n231_));
  XOR2_X1   g030(.A(new_n231_), .B(KEYINPUT89), .Z(new_n232_));
  NAND2_X1  g031(.A1(new_n207_), .A2(new_n204_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n233_), .B1(G183gat), .B2(G190gat), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n216_), .B1(new_n234_), .B2(KEYINPUT90), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n232_), .B(new_n235_), .C1(KEYINPUT90), .C2(new_n234_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n226_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G71gat), .B(G99gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(G43gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n237_), .B(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(KEYINPUT92), .B(KEYINPUT31), .Z(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT91), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G127gat), .B(G134gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G113gat), .B(G120gat), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n243_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(new_n244_), .B(new_n245_), .Z(new_n247_));
  OAI21_X1  g046(.A(new_n246_), .B1(new_n247_), .B2(new_n243_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G227gat), .A2(G233gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(G15gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT30), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n248_), .B(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n242_), .B(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(G197gat), .B(G204gat), .Z(new_n254_));
  OR2_X1    g053(.A1(new_n254_), .A2(KEYINPUT21), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(KEYINPUT21), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G211gat), .B(G218gat), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n256_), .A2(new_n257_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(G141gat), .ZN(new_n262_));
  INV_X1    g061(.A(G148gat), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n263_), .ZN(new_n265_));
  AOI22_X1  g064(.A1(new_n264_), .A2(KEYINPUT2), .B1(new_n265_), .B2(KEYINPUT3), .ZN(new_n266_));
  NOR2_X1   g065(.A1(G141gat), .A2(G148gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT3), .ZN(new_n268_));
  AOI21_X1  g067(.A(KEYINPUT93), .B1(new_n267_), .B2(new_n268_), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n267_), .A2(KEYINPUT93), .A3(new_n268_), .ZN(new_n270_));
  OAI221_X1 g069(.A(new_n266_), .B1(KEYINPUT2), .B2(new_n264_), .C1(new_n269_), .C2(new_n270_), .ZN(new_n271_));
  OR2_X1    g070(.A1(G155gat), .A2(G162gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G155gat), .A2(G162gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n274_), .B(KEYINPUT94), .Z(new_n275_));
  NAND2_X1  g074(.A1(new_n271_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT95), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n272_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n279_), .B1(KEYINPUT1), .B2(new_n273_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n280_), .B1(KEYINPUT1), .B2(new_n273_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n264_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n281_), .A2(new_n265_), .A3(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n278_), .A2(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n261_), .B1(new_n284_), .B2(KEYINPUT29), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G228gat), .A2(G233gat), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n285_), .B1(KEYINPUT96), .B2(new_n286_), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n286_), .B(KEYINPUT96), .Z(new_n288_));
  OAI21_X1  g087(.A(new_n287_), .B1(new_n285_), .B2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G78gat), .B(G106gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT97), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n284_), .A2(KEYINPUT29), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G22gat), .B(G50gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT28), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n293_), .B(new_n295_), .Z(new_n296_));
  NAND2_X1  g095(.A1(new_n292_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n289_), .B(new_n290_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n289_), .A2(new_n290_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n292_), .A2(new_n300_), .A3(new_n291_), .A4(new_n296_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT101), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n278_), .A2(new_n283_), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n304_), .A2(new_n248_), .ZN(new_n305_));
  XOR2_X1   g104(.A(new_n247_), .B(KEYINPUT99), .Z(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n305_), .A2(KEYINPUT4), .A3(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT100), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G225gat), .A2(G233gat), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n304_), .A2(new_n248_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT4), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n310_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n308_), .A2(new_n309_), .A3(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n311_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n310_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G1gat), .B(G29gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(G85gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT0), .B(G57gat), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n319_), .B(new_n320_), .Z(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n309_), .B1(new_n308_), .B2(new_n313_), .ZN(new_n323_));
  NOR3_X1   g122(.A1(new_n317_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n303_), .B1(new_n324_), .B2(KEYINPUT33), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n226_), .A2(new_n261_), .A3(new_n236_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT20), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n208_), .B1(G183gat), .B2(G190gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT22), .B(G169gat), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n216_), .B1(new_n329_), .B2(new_n227_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n221_), .A2(new_n218_), .A3(new_n222_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n233_), .A2(new_n217_), .A3(new_n332_), .A4(new_n211_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n327_), .B1(new_n334_), .B2(new_n260_), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n326_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G226gat), .A2(G233gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT19), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n338_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n261_), .B1(new_n226_), .B2(new_n236_), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT20), .B1(new_n334_), .B2(new_n260_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n340_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G8gat), .B(G36gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT18), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G64gat), .B(G92gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n345_), .B(new_n346_), .Z(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n339_), .A2(new_n343_), .A3(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n348_), .B1(new_n339_), .B2(new_n343_), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT98), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n351_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT98), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(new_n354_), .A3(new_n349_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n315_), .A2(G225gat), .A3(G233gat), .ZN(new_n356_));
  INV_X1    g155(.A(new_n308_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n310_), .B1(new_n305_), .B2(KEYINPUT4), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n356_), .B(new_n322_), .C1(new_n357_), .C2(new_n358_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n352_), .A2(new_n355_), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n324_), .A2(KEYINPUT33), .ZN(new_n361_));
  INV_X1    g160(.A(new_n323_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n362_), .A2(new_n321_), .A3(new_n316_), .A4(new_n314_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT33), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n363_), .A2(KEYINPUT101), .A3(new_n364_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n325_), .A2(new_n360_), .A3(new_n361_), .A4(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n322_), .B1(new_n317_), .B2(new_n323_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(new_n363_), .ZN(new_n368_));
  AOI22_X1  g167(.A1(new_n339_), .A2(new_n343_), .B1(KEYINPUT32), .B2(new_n347_), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n369_), .B(KEYINPUT102), .Z(new_n370_));
  AOI21_X1  g169(.A(new_n260_), .B1(new_n334_), .B2(KEYINPUT104), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n371_), .B1(KEYINPUT104), .B2(new_n334_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT103), .B(KEYINPUT20), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(KEYINPUT105), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n341_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(KEYINPUT105), .B1(new_n372_), .B2(new_n373_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n338_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n336_), .A2(new_n340_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n347_), .A2(KEYINPUT32), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n368_), .B(new_n370_), .C1(new_n380_), .C2(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n302_), .B1(new_n366_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n368_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n302_), .ZN(new_n385_));
  OAI211_X1 g184(.A(KEYINPUT27), .B(new_n353_), .C1(new_n380_), .C2(new_n347_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT27), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n387_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n385_), .A2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n253_), .B1(new_n383_), .B2(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n389_), .A2(new_n302_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n368_), .A2(new_n253_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n391_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT69), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G99gat), .A2(G106gat), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT66), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n398_), .A2(KEYINPUT6), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT6), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n400_), .A2(KEYINPUT66), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n397_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(KEYINPUT66), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n398_), .A2(KEYINPUT6), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n403_), .A2(new_n404_), .A3(G99gat), .A4(G106gat), .ZN(new_n405_));
  OR2_X1    g204(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n406_));
  INV_X1    g205(.A(G106gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n406_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n402_), .A2(new_n405_), .A3(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT64), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(KEYINPUT64), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(G92gat), .B1(KEYINPUT9), .B2(G85gat), .ZN(new_n416_));
  NOR2_X1   g215(.A1(KEYINPUT9), .A2(G85gat), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n415_), .A2(KEYINPUT65), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT65), .B1(new_n415_), .B2(new_n418_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n410_), .B(KEYINPUT67), .C1(new_n419_), .C2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n422_));
  OR3_X1    g221(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n402_), .A2(new_n405_), .A3(new_n422_), .A4(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT8), .ZN(new_n425_));
  INV_X1    g224(.A(G92gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(G85gat), .ZN(new_n427_));
  INV_X1    g226(.A(G85gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(G92gat), .ZN(new_n429_));
  AOI21_X1  g228(.A(KEYINPUT68), .B1(new_n427_), .B2(new_n429_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n424_), .A2(new_n425_), .A3(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n425_), .B1(new_n424_), .B2(new_n430_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n421_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n415_), .A2(new_n418_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT65), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n415_), .A2(KEYINPUT65), .A3(new_n418_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(KEYINPUT67), .B1(new_n438_), .B2(new_n410_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n396_), .B1(new_n433_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n424_), .A2(new_n430_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT8), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n424_), .A2(new_n425_), .A3(new_n430_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n410_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT67), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n444_), .A2(new_n447_), .A3(KEYINPUT69), .A4(new_n421_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n440_), .A2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G57gat), .B(G64gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT11), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT70), .ZN(new_n452_));
  XOR2_X1   g251(.A(G71gat), .B(G78gat), .Z(new_n453_));
  OAI21_X1  g252(.A(new_n453_), .B1(KEYINPUT11), .B2(new_n450_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n452_), .B(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n449_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT12), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n455_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n440_), .A2(new_n448_), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(G230gat), .ZN(new_n461_));
  INV_X1    g260(.A(G233gat), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n460_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT71), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n466_), .B1(new_n433_), .B2(new_n439_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n444_), .A2(new_n447_), .A3(KEYINPUT71), .A4(new_n421_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n467_), .A2(KEYINPUT12), .A3(new_n468_), .A4(new_n455_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n458_), .A2(new_n465_), .A3(KEYINPUT72), .A4(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT72), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n459_), .B1(new_n440_), .B2(new_n448_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n469_), .B1(new_n472_), .B2(KEYINPUT12), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n460_), .A2(new_n464_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n471_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n456_), .A2(new_n460_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(new_n463_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n470_), .A2(new_n475_), .A3(new_n477_), .ZN(new_n478_));
  XOR2_X1   g277(.A(G120gat), .B(G148gat), .Z(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT74), .ZN(new_n480_));
  XOR2_X1   g279(.A(G176gat), .B(G204gat), .Z(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n483_));
  XOR2_X1   g282(.A(new_n482_), .B(new_n483_), .Z(new_n484_));
  NAND2_X1  g283(.A1(new_n478_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n484_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n470_), .A2(new_n475_), .A3(new_n477_), .A4(new_n486_), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n485_), .A2(KEYINPUT13), .A3(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(KEYINPUT13), .B1(new_n485_), .B2(new_n487_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  XOR2_X1   g290(.A(G29gat), .B(G36gat), .Z(new_n492_));
  XOR2_X1   g291(.A(G43gat), .B(G50gat), .Z(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT15), .ZN(new_n495_));
  INV_X1    g294(.A(G1gat), .ZN(new_n496_));
  INV_X1    g295(.A(G8gat), .ZN(new_n497_));
  OAI21_X1  g296(.A(KEYINPUT14), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT78), .B(G15gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n499_), .A2(G22gat), .ZN(new_n500_));
  INV_X1    g299(.A(G15gat), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n501_), .A2(KEYINPUT78), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n501_), .A2(KEYINPUT78), .ZN(new_n503_));
  INV_X1    g302(.A(G22gat), .ZN(new_n504_));
  NOR3_X1   g303(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n498_), .B1(new_n500_), .B2(new_n505_), .ZN(new_n506_));
  XOR2_X1   g305(.A(G1gat), .B(G8gat), .Z(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n507_), .B(new_n498_), .C1(new_n500_), .C2(new_n505_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n495_), .A2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n509_), .A2(new_n494_), .A3(new_n510_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G229gat), .A2(G233gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT82), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n512_), .A2(new_n513_), .A3(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT83), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT81), .ZN(new_n519_));
  INV_X1    g318(.A(new_n513_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n494_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n519_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n521_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n523_), .A2(KEYINPUT81), .A3(new_n513_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n522_), .A2(new_n524_), .A3(G229gat), .A4(G233gat), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n520_), .B1(new_n495_), .B2(new_n511_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n526_), .A2(KEYINPUT83), .A3(new_n515_), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n518_), .A2(new_n525_), .A3(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G113gat), .B(G141gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G169gat), .B(G197gat), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n529_), .B(new_n530_), .Z(new_n531_));
  XNOR2_X1  g330(.A(new_n528_), .B(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n491_), .A2(new_n533_), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n395_), .A2(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(new_n511_), .B(KEYINPUT79), .Z(new_n536_));
  NAND2_X1  g335(.A1(G231gat), .A2(G233gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(new_n459_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G127gat), .B(G155gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT16), .ZN(new_n541_));
  XOR2_X1   g340(.A(G183gat), .B(G211gat), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT17), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n539_), .A2(new_n545_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n538_), .A2(new_n455_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n538_), .A2(new_n455_), .ZN(new_n548_));
  OAI22_X1  g347(.A1(new_n547_), .A2(new_n548_), .B1(new_n544_), .B2(new_n543_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n546_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n467_), .A2(new_n468_), .A3(new_n495_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n440_), .A2(new_n494_), .A3(new_n448_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G232gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT34), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n555_), .B(KEYINPUT35), .Z(new_n556_));
  NAND4_X1  g355(.A1(new_n552_), .A2(new_n553_), .A3(KEYINPUT76), .A4(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n552_), .A2(new_n553_), .A3(new_n556_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT76), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n555_), .A2(KEYINPUT35), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n561_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n557_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G190gat), .B(G218gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G134gat), .B(G162gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT75), .B(KEYINPUT36), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n563_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n566_), .B(KEYINPUT36), .Z(new_n570_));
  OAI211_X1 g369(.A(new_n557_), .B(new_n570_), .C1(new_n560_), .C2(new_n562_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT77), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n569_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n572_), .A2(new_n574_), .A3(KEYINPUT37), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT37), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n569_), .B(new_n571_), .C1(new_n573_), .C2(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n551_), .B1(new_n575_), .B2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT80), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n535_), .A2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n580_), .A2(new_n496_), .A3(new_n368_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT38), .ZN(new_n582_));
  INV_X1    g381(.A(new_n572_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n583_), .B1(new_n391_), .B2(new_n394_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n584_), .A2(new_n550_), .A3(new_n534_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT106), .ZN(new_n586_));
  OAI21_X1  g385(.A(G1gat), .B1(new_n586_), .B2(new_n384_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n582_), .A2(new_n587_), .ZN(G1324gat));
  INV_X1    g387(.A(new_n389_), .ZN(new_n589_));
  OAI21_X1  g388(.A(G8gat), .B1(new_n585_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT107), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n591_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n592_), .A2(KEYINPUT39), .A3(new_n593_), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n593_), .A2(KEYINPUT39), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n580_), .A2(new_n497_), .A3(new_n389_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n594_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT40), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n594_), .A2(new_n595_), .A3(KEYINPUT40), .A4(new_n596_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(G1325gat));
  INV_X1    g400(.A(new_n253_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n580_), .A2(new_n501_), .A3(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(G15gat), .B1(new_n586_), .B2(new_n253_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT41), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n604_), .A2(new_n605_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n603_), .B1(new_n606_), .B2(new_n607_), .ZN(G1326gat));
  NAND3_X1  g407(.A1(new_n580_), .A2(new_n504_), .A3(new_n302_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n302_), .ZN(new_n610_));
  OAI21_X1  g409(.A(G22gat), .B1(new_n586_), .B2(new_n610_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n611_), .A2(KEYINPUT42), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(KEYINPUT42), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n609_), .B1(new_n612_), .B2(new_n613_), .ZN(G1327gat));
  NAND2_X1  g413(.A1(new_n534_), .A2(new_n551_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT108), .Z(new_n616_));
  INV_X1    g415(.A(KEYINPUT43), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n575_), .A2(new_n577_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n617_), .B1(new_n395_), .B2(new_n619_), .ZN(new_n620_));
  AOI211_X1 g419(.A(KEYINPUT43), .B(new_n618_), .C1(new_n391_), .C2(new_n394_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n616_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT44), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  OAI211_X1 g423(.A(KEYINPUT44), .B(new_n616_), .C1(new_n620_), .C2(new_n621_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(new_n368_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(G29gat), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n550_), .A2(new_n572_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n535_), .A2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n384_), .A2(G29gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT109), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n628_), .B1(new_n630_), .B2(new_n632_), .ZN(G1328gat));
  NAND3_X1  g432(.A1(new_n624_), .A2(new_n389_), .A3(new_n625_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(G36gat), .ZN(new_n635_));
  INV_X1    g434(.A(new_n630_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n589_), .A2(G36gat), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT45), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT45), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n636_), .A2(new_n640_), .A3(new_n637_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n635_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT46), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n635_), .A2(new_n642_), .A3(KEYINPUT46), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(G1329gat));
  NAND4_X1  g446(.A1(new_n624_), .A2(G43gat), .A3(new_n602_), .A4(new_n625_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n630_), .A2(new_n253_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n648_), .B1(G43gat), .B2(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g450(.A(G50gat), .B1(new_n636_), .B2(new_n302_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n302_), .A2(G50gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n652_), .B1(new_n626_), .B2(new_n653_), .ZN(G1331gat));
  NOR2_X1   g453(.A1(new_n490_), .A2(new_n532_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(new_n550_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  AND4_X1   g456(.A1(G57gat), .A2(new_n584_), .A3(new_n368_), .A4(new_n657_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n579_), .A2(new_n491_), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n659_), .A2(KEYINPUT110), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n532_), .B1(new_n391_), .B2(new_n394_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(KEYINPUT110), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n660_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT111), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n384_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n665_), .B1(new_n664_), .B2(new_n663_), .ZN(new_n666_));
  INV_X1    g465(.A(G57gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n658_), .B1(new_n666_), .B2(new_n667_), .ZN(G1332gat));
  OR3_X1    g467(.A1(new_n663_), .A2(G64gat), .A3(new_n589_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n584_), .A2(new_n389_), .A3(new_n657_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(G64gat), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n671_), .A2(KEYINPUT113), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(KEYINPUT113), .ZN(new_n673_));
  XNOR2_X1  g472(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n672_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n669_), .B1(new_n675_), .B2(new_n676_), .ZN(G1333gat));
  NAND3_X1  g476(.A1(new_n584_), .A2(new_n602_), .A3(new_n657_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(KEYINPUT114), .B(KEYINPUT49), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n678_), .A2(G71gat), .A3(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n678_), .B2(G71gat), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n253_), .A2(G71gat), .ZN(new_n682_));
  OAI22_X1  g481(.A1(new_n680_), .A2(new_n681_), .B1(new_n663_), .B2(new_n682_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT115), .Z(G1334gat));
  INV_X1    g483(.A(KEYINPUT50), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n584_), .A2(new_n302_), .A3(new_n657_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(G78gat), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT116), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n687_), .A2(KEYINPUT116), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n685_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n690_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n692_), .A2(KEYINPUT50), .A3(new_n688_), .ZN(new_n693_));
  OR3_X1    g492(.A1(new_n663_), .A2(G78gat), .A3(new_n610_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n691_), .A2(new_n693_), .A3(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(KEYINPUT117), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT117), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n691_), .A2(new_n693_), .A3(new_n697_), .A4(new_n694_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(G1335gat));
  NAND2_X1  g498(.A1(new_n655_), .A2(new_n551_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n701_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G85gat), .B1(new_n702_), .B2(new_n384_), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n490_), .A2(new_n572_), .A3(new_n550_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n661_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n706_), .A2(new_n428_), .A3(new_n368_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n703_), .A2(new_n707_), .ZN(G1336gat));
  OAI21_X1  g507(.A(G92gat), .B1(new_n702_), .B2(new_n589_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n706_), .A2(new_n426_), .A3(new_n389_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1337gat));
  OAI21_X1  g510(.A(G99gat), .B1(new_n702_), .B2(new_n253_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n406_), .A2(new_n408_), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n253_), .A2(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n712_), .B1(new_n705_), .B2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g515(.A1(new_n706_), .A2(new_n407_), .A3(new_n302_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n302_), .B(new_n701_), .C1(new_n620_), .C2(new_n621_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT52), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n718_), .A2(new_n719_), .A3(G106gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n718_), .B2(G106gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g522(.A1(new_n392_), .A2(new_n368_), .A3(new_n602_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n485_), .A2(new_n487_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n518_), .A2(new_n525_), .A3(new_n527_), .A4(new_n531_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n522_), .A2(new_n524_), .A3(new_n515_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT119), .ZN(new_n728_));
  INV_X1    g527(.A(new_n531_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n727_), .A2(new_n728_), .A3(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n515_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n526_), .A2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n728_), .B1(new_n727_), .B2(new_n729_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n726_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT120), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT120), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n737_), .B(new_n726_), .C1(new_n733_), .C2(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n725_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT121), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n725_), .A2(KEYINPUT121), .A3(new_n739_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n532_), .A2(new_n487_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT55), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n470_), .A2(new_n475_), .A3(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n473_), .A2(new_n474_), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n460_), .B(new_n469_), .C1(new_n472_), .C2(KEYINPUT12), .ZN(new_n749_));
  AOI22_X1  g548(.A1(new_n748_), .A2(KEYINPUT55), .B1(new_n463_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n747_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(new_n484_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT56), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n751_), .A2(KEYINPUT56), .A3(new_n484_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n745_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  OAI211_X1 g555(.A(KEYINPUT57), .B(new_n572_), .C1(new_n744_), .C2(new_n756_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n739_), .A2(new_n487_), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT56), .B1(new_n751_), .B2(new_n484_), .ZN(new_n759_));
  AOI211_X1 g558(.A(new_n753_), .B(new_n486_), .C1(new_n747_), .C2(new_n750_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n758_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT58), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n758_), .B(KEYINPUT58), .C1(new_n759_), .C2(new_n760_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n763_), .A2(new_n619_), .A3(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n757_), .A2(new_n765_), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n725_), .A2(KEYINPUT121), .A3(new_n739_), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT121), .B1(new_n725_), .B2(new_n739_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n532_), .B(new_n487_), .C1(new_n759_), .C2(new_n760_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n583_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n771_), .A2(KEYINPUT57), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n551_), .B1(new_n766_), .B2(new_n772_), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n488_), .A2(new_n489_), .A3(new_n532_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT54), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n578_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT118), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n578_), .A2(new_n774_), .A3(KEYINPUT118), .A4(new_n775_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n578_), .A2(new_n774_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT54), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n778_), .A2(new_n779_), .A3(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  AOI211_X1 g582(.A(KEYINPUT59), .B(new_n724_), .C1(new_n773_), .C2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(G113gat), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n533_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT123), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT122), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n789_), .B1(new_n771_), .B2(KEYINPUT57), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n572_), .B1(new_n744_), .B2(new_n756_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(KEYINPUT122), .A3(new_n792_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n790_), .A2(new_n793_), .A3(new_n757_), .A4(new_n765_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n551_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n788_), .B1(new_n795_), .B2(new_n783_), .ZN(new_n796_));
  AOI211_X1 g595(.A(KEYINPUT123), .B(new_n782_), .C1(new_n794_), .C2(new_n551_), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n796_), .A2(new_n797_), .A3(new_n724_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT59), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n785_), .B(new_n787_), .C1(new_n798_), .C2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT122), .B1(new_n791_), .B2(new_n792_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n801_), .A2(new_n766_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n550_), .B1(new_n802_), .B2(new_n793_), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT123), .B1(new_n803_), .B2(new_n782_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n795_), .A2(new_n788_), .A3(new_n783_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n724_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n804_), .A2(new_n532_), .A3(new_n805_), .A4(new_n806_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n807_), .A2(KEYINPUT124), .A3(new_n786_), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT124), .B1(new_n807_), .B2(new_n786_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n800_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT125), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT125), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n800_), .B(new_n812_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n813_), .ZN(G1340gat));
  NOR2_X1   g613(.A1(new_n796_), .A2(new_n797_), .ZN(new_n815_));
  INV_X1    g614(.A(G120gat), .ZN(new_n816_));
  OR2_X1    g615(.A1(new_n816_), .A2(KEYINPUT60), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n816_), .B1(new_n490_), .B2(KEYINPUT60), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n815_), .A2(new_n806_), .A3(new_n817_), .A4(new_n818_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(KEYINPUT126), .ZN(new_n820_));
  INV_X1    g619(.A(new_n798_), .ZN(new_n821_));
  AOI211_X1 g620(.A(new_n490_), .B(new_n784_), .C1(new_n821_), .C2(KEYINPUT59), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n820_), .B1(new_n822_), .B2(new_n816_), .ZN(G1341gat));
  INV_X1    g622(.A(G127gat), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n798_), .A2(new_n824_), .A3(new_n550_), .ZN(new_n825_));
  AOI211_X1 g624(.A(new_n551_), .B(new_n784_), .C1(new_n821_), .C2(KEYINPUT59), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(new_n824_), .ZN(G1342gat));
  INV_X1    g626(.A(G134gat), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n798_), .A2(new_n828_), .A3(new_n583_), .ZN(new_n829_));
  AOI211_X1 g628(.A(new_n618_), .B(new_n784_), .C1(new_n821_), .C2(KEYINPUT59), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(new_n828_), .ZN(G1343gat));
  NOR3_X1   g630(.A1(new_n610_), .A2(new_n384_), .A3(new_n602_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n815_), .A2(new_n589_), .A3(new_n832_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n833_), .A2(new_n533_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(new_n262_), .ZN(G1344gat));
  NOR2_X1   g634(.A1(new_n833_), .A2(new_n490_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(new_n263_), .ZN(G1345gat));
  NOR2_X1   g636(.A1(new_n833_), .A2(new_n551_), .ZN(new_n838_));
  XOR2_X1   g637(.A(KEYINPUT61), .B(G155gat), .Z(new_n839_));
  XNOR2_X1  g638(.A(new_n838_), .B(new_n839_), .ZN(G1346gat));
  OAI21_X1  g639(.A(G162gat), .B1(new_n833_), .B2(new_n618_), .ZN(new_n841_));
  OR2_X1    g640(.A1(new_n572_), .A2(G162gat), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n833_), .B2(new_n842_), .ZN(G1347gat));
  AOI21_X1  g642(.A(new_n302_), .B1(new_n773_), .B2(new_n783_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n393_), .A2(new_n389_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(KEYINPUT127), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n844_), .A2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n532_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n848_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n849_));
  INV_X1    g648(.A(new_n329_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n849_), .B1(new_n850_), .B2(new_n848_), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT62), .B1(new_n848_), .B2(G169gat), .ZN(new_n852_));
  OR2_X1    g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1348gat));
  AOI21_X1  g652(.A(G176gat), .B1(new_n847_), .B2(new_n491_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n796_), .A2(new_n797_), .A3(new_n302_), .ZN(new_n855_));
  AND3_X1   g654(.A1(new_n846_), .A2(G176gat), .A3(new_n491_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n854_), .B1(new_n855_), .B2(new_n856_), .ZN(G1349gat));
  AND2_X1   g656(.A1(new_n846_), .A2(new_n550_), .ZN(new_n858_));
  AOI21_X1  g657(.A(G183gat), .B1(new_n855_), .B2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n846_), .A2(new_n550_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n860_), .B1(new_n218_), .B2(new_n222_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n859_), .B1(new_n844_), .B2(new_n861_), .ZN(G1350gat));
  NAND3_X1  g661(.A1(new_n847_), .A2(new_n221_), .A3(new_n583_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n847_), .A2(new_n619_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(new_n203_), .ZN(G1351gat));
  NOR3_X1   g664(.A1(new_n385_), .A2(new_n589_), .A3(new_n602_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n815_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(new_n532_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n491_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g671(.A1(new_n867_), .A2(new_n551_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n873_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n874_));
  XOR2_X1   g673(.A(KEYINPUT63), .B(G211gat), .Z(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n873_), .B2(new_n875_), .ZN(G1354gat));
  OAI21_X1  g675(.A(G218gat), .B1(new_n867_), .B2(new_n618_), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n572_), .A2(G218gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n867_), .B2(new_n878_), .ZN(G1355gat));
endmodule


