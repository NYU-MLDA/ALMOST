//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 1 0 1 0 0 1 0 0 0 1 1 0 1 1 1 0 1 1 1 0 0 0 1 0 1 1 1 1 0 0 1 1 1 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n870_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G29gat), .B(G36gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(new_n210_), .ZN(new_n212_));
  AND2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n208_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G229gat), .A2(G233gat), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n211_), .A2(new_n212_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT15), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(new_n208_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n208_), .B(new_n213_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n215_), .ZN(new_n221_));
  AOI22_X1  g020(.A1(new_n216_), .A2(new_n219_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G113gat), .B(G141gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(KEYINPUT74), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G169gat), .B(G197gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n222_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n222_), .A2(new_n226_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT75), .ZN(new_n232_));
  OR3_X1    g031(.A1(new_n228_), .A2(KEYINPUT75), .A3(new_n229_), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(G228gat), .ZN(new_n235_));
  INV_X1    g034(.A(G233gat), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT84), .ZN(new_n239_));
  INV_X1    g038(.A(G155gat), .ZN(new_n240_));
  INV_X1    g039(.A(G162gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G155gat), .A2(G162gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT1), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT85), .B1(new_n245_), .B2(KEYINPUT1), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT85), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT1), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n248_), .A2(new_n249_), .A3(G155gat), .A4(G162gat), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n244_), .A2(new_n246_), .A3(new_n247_), .A4(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(G141gat), .B(G148gat), .Z(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  OR3_X1    g052(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G141gat), .A2(G148gat), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT2), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n254_), .A2(new_n257_), .A3(new_n258_), .A4(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n260_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n253_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT29), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G197gat), .B(G204gat), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT21), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(G218gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(G211gat), .ZN(new_n268_));
  INV_X1    g067(.A(G211gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(G218gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT89), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n268_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n271_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n264_), .A2(new_n265_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT88), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n266_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n266_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT88), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n279_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n278_), .B(new_n280_), .C1(new_n272_), .C2(new_n273_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n277_), .A2(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n238_), .B1(new_n263_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n263_), .A2(new_n282_), .A3(new_n238_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G78gat), .B(G106gat), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n284_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n285_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n286_), .B1(new_n289_), .B2(new_n283_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT90), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n288_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  OAI211_X1 g091(.A(KEYINPUT90), .B(new_n286_), .C1(new_n289_), .C2(new_n283_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n262_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT29), .ZN(new_n295_));
  XOR2_X1   g094(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n294_), .A2(new_n295_), .A3(new_n297_), .ZN(new_n298_));
  XOR2_X1   g097(.A(G22gat), .B(G50gat), .Z(new_n299_));
  OAI21_X1  g098(.A(new_n296_), .B1(new_n262_), .B2(KEYINPUT29), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n298_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n299_), .B1(new_n298_), .B2(new_n300_), .ZN(new_n303_));
  NOR3_X1   g102(.A1(new_n302_), .A2(new_n303_), .A3(KEYINPUT87), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT87), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n298_), .A2(new_n300_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n299_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n305_), .B1(new_n308_), .B2(new_n301_), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n292_), .B(new_n293_), .C1(new_n304_), .C2(new_n309_), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n288_), .A2(new_n290_), .A3(new_n301_), .A4(new_n308_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G226gat), .A2(G233gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT19), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT22), .B(G169gat), .ZN(new_n318_));
  INV_X1    g117(.A(G176gat), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n317_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G183gat), .A2(G190gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT23), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT23), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n323_), .A2(G183gat), .A3(G190gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(G183gat), .A2(G190gat), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT91), .B1(new_n325_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT91), .ZN(new_n329_));
  AOI211_X1 g128(.A(new_n329_), .B(new_n326_), .C1(new_n322_), .C2(new_n324_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n320_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n322_), .A2(new_n324_), .A3(KEYINPUT79), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT79), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n321_), .A2(new_n333_), .A3(KEYINPUT23), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(G169gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n319_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n337_), .A2(KEYINPUT24), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT25), .B(G183gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(KEYINPUT26), .B(G190gat), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n338_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n337_), .A2(KEYINPUT24), .A3(new_n316_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n335_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n331_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT92), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n282_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n345_), .B1(new_n282_), .B2(new_n344_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n332_), .A2(new_n327_), .A3(new_n334_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT80), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT22), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT77), .B1(new_n352_), .B2(G169gat), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n354_), .A2(new_n336_), .A3(KEYINPUT22), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n353_), .A2(new_n355_), .A3(new_n319_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n357_), .B1(new_n336_), .B2(KEYINPUT22), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n352_), .A2(KEYINPUT78), .A3(G169gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n317_), .B1(new_n356_), .B2(new_n360_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n332_), .A2(KEYINPUT80), .A3(new_n327_), .A4(new_n334_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n351_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n342_), .A2(KEYINPUT76), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n342_), .A2(KEYINPUT76), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n364_), .A2(new_n341_), .A3(new_n325_), .A4(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n363_), .A2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT20), .B1(new_n367_), .B2(new_n282_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n315_), .B1(new_n348_), .B2(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(G8gat), .B(G36gat), .Z(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT18), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G64gat), .B(G92gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n315_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT20), .ZN(new_n375_));
  INV_X1    g174(.A(new_n282_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n344_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n375_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n367_), .A2(KEYINPUT93), .A3(new_n282_), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT93), .B1(new_n367_), .B2(new_n282_), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n374_), .B(new_n378_), .C1(new_n379_), .C2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n369_), .A2(new_n373_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT27), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n282_), .A2(new_n344_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT92), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n282_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n368_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(KEYINPUT96), .B1(new_n388_), .B2(new_n374_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n378_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n315_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n388_), .A2(new_n374_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n389_), .B1(new_n393_), .B2(KEYINPUT96), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n384_), .B1(new_n394_), .B2(new_n373_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n373_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n381_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n386_), .A2(new_n387_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n368_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n374_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n396_), .B1(new_n397_), .B2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n382_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT27), .ZN(new_n403_));
  AOI21_X1  g202(.A(KEYINPUT98), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT98), .ZN(new_n405_));
  AOI211_X1 g204(.A(new_n405_), .B(KEYINPUT27), .C1(new_n401_), .C2(new_n382_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n313_), .B(new_n395_), .C1(new_n404_), .C2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G227gat), .A2(G233gat), .ZN(new_n408_));
  INV_X1    g207(.A(G15gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT30), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n367_), .B(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT81), .B(G43gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(G134gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(G127gat), .ZN(new_n416_));
  INV_X1    g215(.A(G127gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(G134gat), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n416_), .A2(new_n418_), .A3(KEYINPUT82), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT82), .B1(new_n416_), .B2(new_n418_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G113gat), .B(G120gat), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n419_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  XOR2_X1   g221(.A(G113gat), .B(G120gat), .Z(new_n423_));
  INV_X1    g222(.A(KEYINPUT82), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n417_), .A2(G134gat), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n415_), .A2(G127gat), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n424_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n416_), .A2(new_n418_), .A3(KEYINPUT82), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n423_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT83), .B1(new_n422_), .B2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n427_), .A2(new_n428_), .A3(new_n423_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT83), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n430_), .A2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT31), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G71gat), .B(G99gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n435_), .A2(new_n436_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n414_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n414_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n430_), .A2(new_n433_), .A3(new_n262_), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n253_), .B(new_n261_), .C1(new_n422_), .C2(new_n429_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(KEYINPUT4), .A3(new_n444_), .ZN(new_n445_));
  XOR2_X1   g244(.A(KEYINPUT94), .B(KEYINPUT4), .Z(new_n446_));
  NAND4_X1  g245(.A1(new_n430_), .A2(new_n262_), .A3(new_n433_), .A4(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G225gat), .A2(G233gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G1gat), .B(G29gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(G85gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT0), .B(G57gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n450_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n451_), .A2(new_n455_), .A3(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n455_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n449_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n459_), .B1(new_n460_), .B2(new_n456_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n458_), .A2(KEYINPUT97), .A3(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT97), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n451_), .A2(new_n457_), .A3(new_n463_), .A4(new_n455_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n442_), .A2(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n407_), .A2(new_n466_), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n310_), .A2(new_n311_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n395_), .B(new_n468_), .C1(new_n404_), .C2(new_n406_), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n445_), .A2(new_n449_), .A3(new_n447_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n443_), .A2(new_n450_), .A3(new_n444_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n455_), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT33), .B1(new_n470_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(new_n461_), .ZN(new_n474_));
  OAI211_X1 g273(.A(KEYINPUT33), .B(new_n459_), .C1(new_n460_), .C2(new_n456_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n401_), .A2(new_n474_), .A3(new_n382_), .A4(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n373_), .A2(KEYINPUT32), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT93), .ZN(new_n478_));
  AND2_X1   g277(.A1(new_n363_), .A2(new_n366_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n478_), .B1(new_n479_), .B2(new_n376_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n367_), .A2(KEYINPUT93), .A3(new_n282_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n374_), .B1(new_n482_), .B2(new_n378_), .ZN(new_n483_));
  NOR3_X1   g282(.A1(new_n348_), .A2(new_n315_), .A3(new_n368_), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT96), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n389_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n477_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n477_), .B(KEYINPUT95), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n369_), .A2(new_n488_), .A3(new_n381_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n462_), .A2(new_n464_), .A3(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n476_), .B1(new_n487_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(new_n313_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n442_), .B1(new_n469_), .B2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT99), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n467_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n485_), .A2(new_n486_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n383_), .B1(new_n496_), .B2(new_n396_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n312_), .A2(new_n465_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n382_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n373_), .B1(new_n369_), .B2(new_n381_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n403_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(new_n405_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n402_), .A2(KEYINPUT98), .A3(new_n403_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  AOI22_X1  g304(.A1(new_n499_), .A2(new_n505_), .B1(new_n313_), .B2(new_n491_), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT99), .B1(new_n506_), .B2(new_n442_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n234_), .B1(new_n495_), .B2(new_n507_), .ZN(new_n508_));
  OR2_X1    g307(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n509_));
  INV_X1    g308(.A(G106gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n509_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT65), .B(G85gat), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT9), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(G92gat), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n512_), .B1(new_n513_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G99gat), .A2(G106gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT6), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT6), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n519_), .A2(G99gat), .A3(G106gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G85gat), .B(G92gat), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n521_), .B1(new_n522_), .B2(new_n514_), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT66), .B1(new_n516_), .B2(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(G85gat), .B(G92gat), .Z(new_n525_));
  AOI22_X1  g324(.A1(new_n525_), .A2(KEYINPUT9), .B1(new_n518_), .B2(new_n520_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT66), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n513_), .A2(new_n515_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n526_), .A2(new_n527_), .A3(new_n512_), .A4(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT7), .ZN(new_n531_));
  INV_X1    g330(.A(G99gat), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(new_n532_), .A3(new_n510_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n521_), .A2(new_n530_), .A3(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(new_n525_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT8), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT8), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n534_), .A2(new_n537_), .A3(new_n525_), .ZN(new_n538_));
  AOI22_X1  g337(.A1(new_n524_), .A2(new_n529_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G57gat), .B(G64gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT11), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT67), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT67), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n540_), .A2(new_n543_), .A3(KEYINPUT11), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n540_), .A2(KEYINPUT11), .ZN(new_n546_));
  XOR2_X1   g345(.A(G71gat), .B(G78gat), .Z(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n545_), .A2(new_n548_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n542_), .A2(new_n546_), .A3(new_n547_), .A4(new_n544_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n539_), .A2(new_n551_), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n552_), .A2(KEYINPUT68), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G230gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT64), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n539_), .A2(new_n551_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n552_), .A2(KEYINPUT68), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n553_), .B(new_n555_), .C1(new_n556_), .C2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT12), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n559_), .B1(new_n539_), .B2(new_n551_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n551_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n529_), .A2(new_n524_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n536_), .A2(new_n538_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n561_), .A2(new_n564_), .A3(KEYINPUT12), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n555_), .B1(new_n539_), .B2(new_n551_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n560_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n558_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G176gat), .B(G204gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT70), .ZN(new_n570_));
  XOR2_X1   g369(.A(KEYINPUT69), .B(KEYINPUT5), .Z(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G120gat), .B(G148gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n568_), .A2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n558_), .A2(new_n567_), .A3(new_n574_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT13), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT13), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n576_), .A2(new_n580_), .A3(new_n577_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT34), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n584_), .B(KEYINPUT35), .Z(new_n585_));
  NOR2_X1   g384(.A1(new_n564_), .A2(new_n217_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n539_), .A2(new_n218_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n585_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(KEYINPUT71), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT71), .ZN(new_n590_));
  OAI211_X1 g389(.A(new_n590_), .B(new_n585_), .C1(new_n586_), .C2(new_n587_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n586_), .A2(new_n587_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n584_), .A2(KEYINPUT35), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n589_), .B(new_n591_), .C1(new_n592_), .C2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G190gat), .B(G218gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G134gat), .B(G162gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n597_), .B(KEYINPUT36), .Z(new_n598_));
  NAND2_X1  g397(.A1(new_n594_), .A2(new_n598_), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n592_), .A2(new_n593_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n597_), .A2(KEYINPUT36), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n600_), .A2(new_n589_), .A3(new_n591_), .A4(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n599_), .A2(KEYINPUT37), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(KEYINPUT72), .B1(new_n594_), .B2(new_n598_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n594_), .A2(KEYINPUT72), .A3(new_n598_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n606_), .A2(new_n602_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT37), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n604_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(G127gat), .B(G155gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT16), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G183gat), .B(G211gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n614_), .B(KEYINPUT17), .Z(new_n615_));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n208_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(new_n551_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n615_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n614_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n618_), .B1(KEYINPUT17), .B2(new_n621_), .ZN(new_n622_));
  OR3_X1    g421(.A1(new_n620_), .A2(new_n622_), .A3(KEYINPUT73), .ZN(new_n623_));
  OAI21_X1  g422(.A(KEYINPUT73), .B1(new_n620_), .B2(new_n622_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n610_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n508_), .A2(new_n582_), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n465_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(new_n203_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT38), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT100), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n607_), .A2(new_n602_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n634_), .A2(new_n605_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n495_), .B2(new_n507_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n582_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n637_), .A2(new_n230_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n636_), .A2(new_n625_), .A3(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(G1gat), .B1(new_n639_), .B2(new_n465_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n633_), .B(new_n640_), .C1(new_n631_), .C2(new_n630_), .ZN(G1324gat));
  NAND2_X1  g440(.A1(new_n505_), .A2(new_n395_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n628_), .A2(new_n204_), .A3(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n642_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G8gat), .B1(new_n639_), .B2(new_n644_), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n645_), .A2(KEYINPUT101), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT39), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(KEYINPUT101), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n646_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n647_), .B1(new_n646_), .B2(new_n648_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n643_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT40), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  OAI211_X1 g452(.A(KEYINPUT40), .B(new_n643_), .C1(new_n649_), .C2(new_n650_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1325gat));
  INV_X1    g454(.A(new_n442_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G15gat), .B1(new_n639_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT41), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n657_), .B(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n628_), .A2(new_n409_), .A3(new_n442_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT102), .ZN(G1326gat));
  INV_X1    g461(.A(G22gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n628_), .A2(new_n663_), .A3(new_n312_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G22gat), .B1(new_n639_), .B2(new_n313_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n665_), .A2(new_n666_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n664_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT104), .Z(G1327gat));
  NOR3_X1   g469(.A1(new_n637_), .A2(new_n608_), .A3(new_n625_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n508_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(G29gat), .B1(new_n673_), .B2(new_n629_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n495_), .A2(new_n507_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n610_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n676_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  AOI211_X1 g478(.A(KEYINPUT43), .B(new_n610_), .C1(new_n495_), .C2(new_n507_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n625_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n638_), .A2(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n675_), .B1(new_n681_), .B2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n469_), .A2(new_n492_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n685_), .A2(new_n494_), .A3(new_n656_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n467_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n493_), .A2(new_n494_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n678_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT43), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n677_), .A2(new_n676_), .A3(new_n678_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n693_), .A2(KEYINPUT44), .A3(new_n682_), .A4(new_n638_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n684_), .A2(new_n694_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n629_), .A2(G29gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n674_), .B1(new_n695_), .B2(new_n696_), .ZN(G1328gat));
  NOR3_X1   g496(.A1(new_n672_), .A2(G36gat), .A3(new_n644_), .ZN(new_n698_));
  XOR2_X1   g497(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n699_));
  XNOR2_X1  g498(.A(new_n698_), .B(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n684_), .A2(new_n694_), .A3(new_n642_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(G36gat), .B2(new_n701_), .ZN(new_n702_));
  XOR2_X1   g501(.A(KEYINPUT106), .B(KEYINPUT46), .Z(new_n703_));
  OAI21_X1  g502(.A(KEYINPUT107), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n705_));
  INV_X1    g504(.A(new_n703_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n701_), .A2(G36gat), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n705_), .B(new_n706_), .C1(new_n707_), .C2(new_n700_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n702_), .A2(KEYINPUT46), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n704_), .A2(new_n708_), .A3(new_n709_), .ZN(G1329gat));
  NAND4_X1  g509(.A1(new_n684_), .A2(new_n694_), .A3(G43gat), .A4(new_n442_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n672_), .A2(new_n656_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n711_), .B1(G43gat), .B2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g513(.A(G50gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n673_), .A2(new_n715_), .A3(new_n312_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT108), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n695_), .A2(new_n312_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n718_), .B2(G50gat), .ZN(new_n719_));
  AOI211_X1 g518(.A(KEYINPUT108), .B(new_n715_), .C1(new_n695_), .C2(new_n312_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n716_), .B1(new_n719_), .B2(new_n720_), .ZN(G1331gat));
  AND3_X1   g520(.A1(new_n637_), .A2(new_n234_), .A3(new_n625_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n636_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(G57gat), .B1(new_n724_), .B2(new_n465_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n231_), .B1(new_n495_), .B2(new_n507_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n726_), .A2(new_n637_), .A3(new_n627_), .ZN(new_n727_));
  INV_X1    g526(.A(G57gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n727_), .A2(new_n728_), .A3(new_n629_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n725_), .A2(new_n729_), .ZN(G1332gat));
  INV_X1    g529(.A(G64gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(new_n723_), .B2(new_n642_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT48), .Z(new_n733_));
  NAND3_X1  g532(.A1(new_n727_), .A2(new_n731_), .A3(new_n642_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1333gat));
  INV_X1    g534(.A(G71gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n736_), .B1(new_n723_), .B2(new_n442_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT49), .Z(new_n738_));
  NAND3_X1  g537(.A1(new_n727_), .A2(new_n736_), .A3(new_n442_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1334gat));
  INV_X1    g539(.A(G78gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n723_), .B2(new_n312_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n742_), .B(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n727_), .A2(new_n741_), .A3(new_n312_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1335gat));
  AND4_X1   g545(.A1(new_n637_), .A2(new_n726_), .A3(new_n635_), .A4(new_n682_), .ZN(new_n747_));
  AOI21_X1  g546(.A(G85gat), .B1(new_n747_), .B2(new_n629_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n582_), .A2(new_n625_), .A3(new_n231_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n750_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n465_), .A2(new_n513_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(G1336gat));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n642_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n644_), .A2(G92gat), .ZN(new_n755_));
  AOI22_X1  g554(.A1(new_n754_), .A2(G92gat), .B1(new_n747_), .B2(new_n755_), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT110), .Z(G1337gat));
  AOI21_X1  g556(.A(new_n532_), .B1(new_n751_), .B2(new_n442_), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n442_), .A2(new_n509_), .A3(new_n511_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n747_), .B2(new_n759_), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT51), .Z(G1338gat));
  XNOR2_X1  g560(.A(KEYINPUT112), .B(KEYINPUT52), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n312_), .B(new_n749_), .C1(new_n679_), .C2(new_n680_), .ZN(new_n764_));
  OAI21_X1  g563(.A(G106gat), .B1(new_n764_), .B2(KEYINPUT111), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT111), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n751_), .B2(new_n312_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n763_), .B1(new_n765_), .B2(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n751_), .A2(new_n766_), .A3(new_n312_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n764_), .A2(KEYINPUT111), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n769_), .A2(new_n770_), .A3(G106gat), .A4(new_n762_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n768_), .A2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n747_), .A2(new_n510_), .A3(new_n312_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT53), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT53), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n772_), .A2(new_n776_), .A3(new_n773_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(G1339gat));
  INV_X1    g577(.A(KEYINPUT121), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n407_), .A2(new_n656_), .A3(new_n465_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT59), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT57), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n231_), .A2(new_n577_), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n560_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n565_), .A2(new_n560_), .A3(new_n552_), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n785_), .A2(KEYINPUT55), .B1(new_n786_), .B2(new_n555_), .ZN(new_n787_));
  XOR2_X1   g586(.A(KEYINPUT114), .B(KEYINPUT55), .Z(new_n788_));
  NAND2_X1  g587(.A1(new_n567_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT115), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT115), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n567_), .A2(new_n791_), .A3(new_n788_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n787_), .A2(new_n790_), .A3(new_n792_), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n793_), .A2(KEYINPUT56), .A3(new_n575_), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT56), .B1(new_n793_), .B2(new_n575_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n784_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n219_), .A2(new_n214_), .A3(new_n221_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n226_), .B1(new_n220_), .B2(new_n215_), .ZN(new_n798_));
  AOI22_X1  g597(.A1(new_n222_), .A2(new_n226_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n578_), .A2(new_n799_), .ZN(new_n800_));
  AOI211_X1 g599(.A(new_n783_), .B(new_n635_), .C1(new_n796_), .C2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n796_), .A2(new_n800_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT57), .B1(new_n803_), .B2(new_n608_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n577_), .A2(new_n799_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(KEYINPUT116), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n793_), .A2(KEYINPUT56), .A3(new_n575_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n807_), .B1(new_n795_), .B2(KEYINPUT117), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n809_));
  AOI211_X1 g608(.A(new_n809_), .B(KEYINPUT56), .C1(new_n793_), .C2(new_n575_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n806_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT58), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n610_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  OAI211_X1 g612(.A(KEYINPUT58), .B(new_n806_), .C1(new_n808_), .C2(new_n810_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n804_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n802_), .B1(new_n815_), .B2(KEYINPUT120), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT120), .ZN(new_n817_));
  AOI211_X1 g616(.A(new_n817_), .B(new_n804_), .C1(new_n814_), .C2(new_n813_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n682_), .B1(new_n816_), .B2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n582_), .A2(new_n234_), .A3(new_n625_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT113), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n582_), .A2(new_n234_), .A3(new_n822_), .A4(new_n625_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n678_), .B1(new_n821_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n824_), .B(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n782_), .B1(new_n819_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(G113gat), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n234_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n804_), .A2(new_n801_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n811_), .A2(new_n812_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT118), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n832_), .A2(new_n833_), .A3(new_n678_), .A4(new_n814_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n831_), .A2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n833_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n682_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n826_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT119), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n837_), .A2(KEYINPUT119), .A3(new_n826_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n841_), .A3(new_n780_), .ZN(new_n842_));
  AOI211_X1 g641(.A(new_n827_), .B(new_n830_), .C1(new_n842_), .C2(KEYINPUT59), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n840_), .A2(new_n841_), .A3(new_n780_), .ZN(new_n844_));
  AOI21_X1  g643(.A(G113gat), .B1(new_n844_), .B2(new_n231_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n779_), .B1(new_n843_), .B2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n827_), .B1(new_n842_), .B2(KEYINPUT59), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n829_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n828_), .B1(new_n842_), .B2(new_n230_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(KEYINPUT121), .A3(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n846_), .A2(new_n850_), .ZN(G1340gat));
  INV_X1    g650(.A(G120gat), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n852_), .B1(new_n582_), .B2(KEYINPUT60), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n844_), .B(new_n853_), .C1(KEYINPUT60), .C2(new_n852_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n847_), .A2(new_n637_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n852_), .ZN(G1341gat));
  NAND3_X1  g655(.A1(new_n844_), .A2(new_n417_), .A3(new_n625_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n847_), .A2(new_n625_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n417_), .ZN(G1342gat));
  AOI21_X1  g658(.A(G134gat), .B1(new_n844_), .B2(new_n635_), .ZN(new_n860_));
  XOR2_X1   g659(.A(KEYINPUT122), .B(G134gat), .Z(new_n861_));
  NOR2_X1   g660(.A1(new_n610_), .A2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n860_), .B1(new_n847_), .B2(new_n862_), .ZN(G1343gat));
  AND2_X1   g662(.A1(new_n840_), .A2(new_n841_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n442_), .A2(new_n313_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n644_), .A2(new_n629_), .A3(new_n865_), .ZN(new_n866_));
  XOR2_X1   g665(.A(new_n866_), .B(KEYINPUT123), .Z(new_n867_));
  NAND3_X1  g666(.A1(new_n864_), .A2(new_n231_), .A3(new_n867_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g668(.A1(new_n864_), .A2(new_n637_), .A3(new_n867_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g670(.A1(new_n864_), .A2(new_n625_), .A3(new_n867_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(KEYINPUT61), .B(G155gat), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1346gat));
  NAND2_X1  g673(.A1(new_n864_), .A2(new_n867_), .ZN(new_n875_));
  OAI21_X1  g674(.A(G162gat), .B1(new_n875_), .B2(new_n610_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n635_), .A2(new_n241_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n875_), .B2(new_n877_), .ZN(G1347gat));
  INV_X1    g677(.A(KEYINPUT62), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n819_), .A2(new_n826_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n644_), .A2(new_n466_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n313_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n880_), .A2(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n230_), .ZN(new_n885_));
  OAI211_X1 g684(.A(KEYINPUT124), .B(new_n879_), .C1(new_n885_), .C2(new_n336_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n318_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT124), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n336_), .B1(new_n888_), .B2(KEYINPUT62), .ZN(new_n889_));
  OAI221_X1 g688(.A(new_n889_), .B1(new_n888_), .B2(KEYINPUT62), .C1(new_n884_), .C2(new_n230_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n886_), .A2(new_n887_), .A3(new_n890_), .ZN(G1348gat));
  INV_X1    g690(.A(new_n884_), .ZN(new_n892_));
  AOI21_X1  g691(.A(G176gat), .B1(new_n892_), .B2(new_n637_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n864_), .A2(new_n313_), .ZN(new_n894_));
  NOR4_X1   g693(.A1(new_n644_), .A2(new_n319_), .A3(new_n466_), .A4(new_n582_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n893_), .B1(new_n894_), .B2(new_n895_), .ZN(G1349gat));
  NOR3_X1   g695(.A1(new_n884_), .A2(new_n339_), .A3(new_n682_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n894_), .A2(new_n625_), .A3(new_n881_), .ZN(new_n898_));
  INV_X1    g697(.A(G183gat), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n897_), .B1(new_n898_), .B2(new_n899_), .ZN(G1350gat));
  OAI21_X1  g699(.A(G190gat), .B1(new_n884_), .B2(new_n610_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n635_), .A2(new_n340_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n884_), .B2(new_n902_), .ZN(G1351gat));
  AND3_X1   g702(.A1(new_n642_), .A2(new_n465_), .A3(new_n865_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n864_), .A2(new_n231_), .A3(new_n904_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g705(.A1(new_n864_), .A2(new_n637_), .A3(new_n904_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g707(.A(new_n682_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(KEYINPUT125), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n864_), .A2(new_n904_), .A3(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(KEYINPUT126), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n911_), .B(new_n913_), .ZN(G1354gat));
  NAND2_X1  g713(.A1(new_n864_), .A2(new_n904_), .ZN(new_n915_));
  OAI21_X1  g714(.A(G218gat), .B1(new_n915_), .B2(new_n610_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n635_), .A2(new_n267_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n915_), .B2(new_n917_), .ZN(G1355gat));
endmodule


