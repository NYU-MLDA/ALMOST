//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 1 0 0 1 1 1 1 1 0 1 1 0 0 1 1 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n777_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n902_, new_n904_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n927_, new_n929_, new_n930_,
    new_n931_, new_n933_, new_n934_, new_n935_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT93), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT23), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT23), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n206_), .A2(G183gat), .A3(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT24), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n208_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT25), .ZN(new_n213_));
  INV_X1    g012(.A(G183gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n213_), .B1(new_n214_), .B2(KEYINPUT79), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT79), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(KEYINPUT25), .A3(G183gat), .ZN(new_n217_));
  OR2_X1    g016(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n219_));
  AOI22_X1  g018(.A1(new_n215_), .A2(new_n217_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n212_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G169gat), .ZN(new_n222_));
  INV_X1    g021(.A(G176gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(KEYINPUT24), .A3(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(KEYINPUT80), .A2(G169gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT22), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT22), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(KEYINPUT80), .A3(G169gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n230_), .A3(new_n223_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n231_), .A2(new_n225_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n205_), .A2(new_n207_), .A3(KEYINPUT81), .ZN(new_n233_));
  INV_X1    g032(.A(G190gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n214_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT81), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n236_), .A2(new_n206_), .A3(G183gat), .A4(G190gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n233_), .A2(new_n235_), .A3(new_n237_), .ZN(new_n238_));
  AOI22_X1  g037(.A1(new_n221_), .A2(new_n226_), .B1(new_n232_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G197gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(G204gat), .ZN(new_n241_));
  INV_X1    g040(.A(G204gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(G197gat), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT88), .B1(new_n242_), .B2(G197gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT21), .ZN(new_n246_));
  AND2_X1   g045(.A1(G211gat), .A2(G218gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(G211gat), .A2(G218gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n244_), .B1(new_n246_), .B2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G211gat), .B(G218gat), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n251_), .A2(KEYINPUT21), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n241_), .A2(new_n243_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n253_), .A2(new_n251_), .A3(KEYINPUT21), .A4(new_n245_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n250_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n203_), .B1(new_n239_), .B2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT26), .B(G190gat), .ZN(new_n257_));
  AND3_X1   g056(.A1(new_n216_), .A2(KEYINPUT25), .A3(G183gat), .ZN(new_n258_));
  AOI21_X1  g057(.A(KEYINPUT25), .B1(new_n216_), .B2(G183gat), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n257_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n205_), .A2(new_n207_), .B1(new_n210_), .B2(new_n209_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(new_n226_), .A3(new_n261_), .ZN(new_n262_));
  AND3_X1   g061(.A1(new_n233_), .A2(new_n235_), .A3(new_n237_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n231_), .A2(new_n225_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n262_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n250_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(new_n266_), .A3(KEYINPUT93), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n256_), .A2(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(KEYINPUT22), .B(G169gat), .Z(new_n269_));
  NOR2_X1   g068(.A1(new_n269_), .A2(G176gat), .ZN(new_n270_));
  INV_X1    g069(.A(new_n225_), .ZN(new_n271_));
  AOI22_X1  g070(.A1(new_n205_), .A2(new_n207_), .B1(new_n214_), .B2(new_n234_), .ZN(new_n272_));
  NOR3_X1   g071(.A1(new_n270_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n213_), .A2(G183gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n214_), .A2(KEYINPUT25), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT90), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n277_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n257_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n233_), .A2(new_n237_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n210_), .A2(KEYINPUT91), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT91), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT24), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n224_), .A2(new_n282_), .A3(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n271_), .A2(new_n209_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT91), .B(KEYINPUT24), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n285_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n280_), .A2(new_n281_), .A3(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n274_), .A2(new_n255_), .A3(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n268_), .A2(KEYINPUT20), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G226gat), .A2(G233gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT19), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(KEYINPUT89), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n239_), .A2(new_n255_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT92), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n289_), .A2(new_n297_), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n280_), .A2(new_n281_), .A3(new_n288_), .A4(KEYINPUT92), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n273_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  OAI211_X1 g099(.A(KEYINPUT20), .B(new_n296_), .C1(new_n300_), .C2(new_n255_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n294_), .B1(new_n295_), .B2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT18), .B(G64gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(G92gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G8gat), .B(G36gat), .ZN(new_n305_));
  XOR2_X1   g104(.A(new_n304_), .B(new_n305_), .Z(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n202_), .B1(new_n302_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n301_), .A2(new_n295_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n293_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT20), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  AND3_X1   g111(.A1(new_n265_), .A2(KEYINPUT93), .A3(new_n266_), .ZN(new_n313_));
  AOI21_X1  g112(.A(KEYINPUT93), .B1(new_n265_), .B2(new_n266_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n312_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  AOI211_X1 g114(.A(new_n266_), .B(new_n273_), .C1(new_n298_), .C2(new_n299_), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT94), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n311_), .B1(new_n256_), .B2(new_n267_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT94), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n233_), .A2(new_n237_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n214_), .A2(KEYINPUT25), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n213_), .A2(G183gat), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT90), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n320_), .B1(new_n325_), .B2(new_n257_), .ZN(new_n326_));
  AOI21_X1  g125(.A(KEYINPUT92), .B1(new_n326_), .B2(new_n288_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n299_), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n255_), .B(new_n274_), .C1(new_n327_), .C2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n318_), .A2(new_n319_), .A3(new_n329_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n309_), .A2(new_n317_), .A3(new_n330_), .A4(new_n306_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT100), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n331_), .A2(new_n332_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n308_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT101), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  AND4_X1   g136(.A1(new_n319_), .A2(new_n268_), .A3(new_n329_), .A4(new_n312_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n319_), .B1(new_n318_), .B2(new_n329_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n340_), .A2(KEYINPUT100), .A3(new_n309_), .A4(new_n306_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n331_), .A2(new_n332_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n343_), .A2(KEYINPUT101), .A3(new_n308_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n309_), .A2(new_n317_), .A3(new_n330_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(new_n307_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(new_n331_), .ZN(new_n347_));
  AOI22_X1  g146(.A1(new_n337_), .A2(new_n344_), .B1(new_n202_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT95), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G141gat), .A2(G148gat), .ZN(new_n350_));
  INV_X1    g149(.A(G141gat), .ZN(new_n351_));
  INV_X1    g150(.A(G148gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G155gat), .A2(G162gat), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n354_), .A2(KEYINPUT84), .A3(KEYINPUT1), .ZN(new_n355_));
  NOR2_X1   g154(.A1(G155gat), .A2(G162gat), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT1), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n358_), .A2(G155gat), .A3(G162gat), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n355_), .A2(new_n357_), .A3(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(KEYINPUT84), .B1(new_n354_), .B2(KEYINPUT1), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n350_), .B(new_n353_), .C1(new_n360_), .C2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT86), .ZN(new_n363_));
  INV_X1    g162(.A(new_n354_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n363_), .B1(new_n364_), .B2(new_n356_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n357_), .A2(KEYINPUT86), .A3(new_n354_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT3), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n367_), .A2(new_n351_), .A3(new_n352_), .A4(KEYINPUT85), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT85), .ZN(new_n369_));
  OAI22_X1  g168(.A1(new_n369_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT2), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n350_), .A2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n365_), .B(new_n366_), .C1(new_n371_), .C2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(G120gat), .ZN(new_n377_));
  OR2_X1    g176(.A1(G127gat), .A2(G134gat), .ZN(new_n378_));
  INV_X1    g177(.A(G113gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G127gat), .A2(G134gat), .ZN(new_n380_));
  AND3_X1   g179(.A1(new_n378_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n379_), .B1(new_n378_), .B2(new_n380_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n377_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n378_), .A2(new_n380_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(G113gat), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n378_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(G120gat), .A3(new_n386_), .ZN(new_n387_));
  AOI22_X1  g186(.A1(new_n362_), .A2(new_n376_), .B1(new_n383_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT4), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n349_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n362_), .A2(new_n376_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n383_), .A2(new_n387_), .ZN(new_n392_));
  AND4_X1   g191(.A1(new_n349_), .A2(new_n391_), .A3(new_n392_), .A4(new_n389_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n390_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n391_), .A2(new_n392_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n362_), .A2(new_n376_), .A3(new_n383_), .A4(new_n387_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n395_), .A2(KEYINPUT4), .A3(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G225gat), .A2(G233gat), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT96), .B1(new_n394_), .B2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT95), .B1(new_n395_), .B2(KEYINPUT4), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n388_), .A2(new_n349_), .A3(new_n389_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT96), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n404_), .A2(new_n405_), .A3(new_n399_), .A4(new_n397_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n395_), .A2(new_n398_), .A3(new_n396_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n401_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT0), .B(G57gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(G85gat), .ZN(new_n410_));
  XOR2_X1   g209(.A(G1gat), .B(G29gat), .Z(new_n411_));
  XOR2_X1   g210(.A(new_n410_), .B(new_n411_), .Z(new_n412_));
  NAND2_X1  g211(.A1(new_n408_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n412_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n401_), .A2(new_n406_), .A3(new_n414_), .A4(new_n407_), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n413_), .A2(KEYINPUT99), .A3(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(KEYINPUT99), .B1(new_n413_), .B2(new_n415_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n255_), .B1(new_n391_), .B2(KEYINPUT29), .ZN(new_n419_));
  INV_X1    g218(.A(G50gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n391_), .A2(KEYINPUT29), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G78gat), .B(G106gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n421_), .B(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G228gat), .A2(G233gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(G22gat), .ZN(new_n427_));
  XOR2_X1   g226(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n428_));
  XNOR2_X1  g227(.A(new_n427_), .B(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n425_), .B(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n265_), .B(new_n392_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT83), .B(KEYINPUT30), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G71gat), .B(G99gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G227gat), .A2(G233gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G15gat), .B(G43gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n434_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n434_), .A2(new_n442_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n348_), .A2(new_n418_), .A3(new_n431_), .A4(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT102), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n431_), .B1(new_n348_), .B2(new_n418_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n309_), .A2(new_n317_), .A3(new_n330_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n306_), .A2(KEYINPUT32), .ZN(new_n452_));
  AOI22_X1  g251(.A1(new_n413_), .A2(new_n415_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n302_), .A2(KEYINPUT32), .A3(new_n306_), .ZN(new_n454_));
  AOI21_X1  g253(.A(KEYINPUT98), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n395_), .A2(new_n396_), .ZN(new_n457_));
  OR2_X1    g256(.A1(new_n457_), .A2(KEYINPUT97), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(KEYINPUT97), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(new_n399_), .A3(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n404_), .A2(new_n398_), .A3(new_n397_), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n460_), .A2(new_n412_), .A3(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n347_), .A2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n415_), .B(KEYINPUT33), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n430_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n453_), .A2(KEYINPUT98), .A3(new_n454_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n456_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(new_n445_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n449_), .B1(new_n450_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n347_), .A2(new_n202_), .ZN(new_n470_));
  AND3_X1   g269(.A1(new_n343_), .A2(KEYINPUT101), .A3(new_n308_), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT101), .B1(new_n343_), .B2(new_n308_), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n418_), .B(new_n470_), .C1(new_n471_), .C2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(new_n430_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n413_), .A2(new_n415_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n451_), .A2(new_n452_), .ZN(new_n476_));
  AND4_X1   g275(.A1(KEYINPUT98), .A2(new_n475_), .A3(new_n454_), .A4(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n477_), .A2(new_n455_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n446_), .B1(new_n478_), .B2(new_n465_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n474_), .A2(new_n479_), .A3(KEYINPUT102), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n448_), .B1(new_n469_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT77), .ZN(new_n482_));
  XOR2_X1   g281(.A(G15gat), .B(G22gat), .Z(new_n483_));
  NAND2_X1  g282(.A1(G1gat), .A2(G8gat), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n483_), .B1(KEYINPUT14), .B2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT74), .ZN(new_n486_));
  XOR2_X1   g285(.A(G1gat), .B(G8gat), .Z(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G29gat), .B(G36gat), .ZN(new_n489_));
  INV_X1    g288(.A(G43gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(G50gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n489_), .B(G43gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n420_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n488_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n487_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n486_), .B(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n495_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n482_), .B1(new_n496_), .B2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G229gat), .A2(G233gat), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n498_), .A2(new_n499_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n488_), .A2(new_n495_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(new_n505_), .A3(KEYINPUT77), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n501_), .A2(KEYINPUT78), .A3(new_n503_), .A4(new_n506_), .ZN(new_n507_));
  AND3_X1   g306(.A1(new_n501_), .A2(new_n503_), .A3(new_n506_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT78), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT15), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n495_), .B(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n496_), .B1(new_n488_), .B2(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n509_), .B1(new_n512_), .B2(new_n502_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n507_), .B1(new_n508_), .B2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G113gat), .B(G141gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(new_n222_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(new_n240_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n514_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n517_), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n507_), .B(new_n519_), .C1(new_n508_), .C2(new_n513_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT13), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G230gat), .A2(G233gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT64), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G85gat), .B(G92gat), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT66), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G99gat), .A2(G106gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT6), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n532_));
  OR3_X1    g331(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n529_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT8), .ZN(new_n536_));
  AOI21_X1  g335(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n537_), .B1(new_n527_), .B2(KEYINPUT9), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT65), .ZN(new_n539_));
  XNOR2_X1  g338(.A(KEYINPUT10), .B(G99gat), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n539_), .B(new_n531_), .C1(G106gat), .C2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n536_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT67), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  XOR2_X1   g343(.A(G57gat), .B(G64gat), .Z(new_n545_));
  INV_X1    g344(.A(KEYINPUT11), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G71gat), .A2(G78gat), .ZN(new_n548_));
  INV_X1    g347(.A(G71gat), .ZN(new_n549_));
  INV_X1    g348(.A(G78gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n547_), .A2(new_n548_), .A3(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT68), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n545_), .A2(new_n546_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n544_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n542_), .B(KEYINPUT67), .ZN(new_n557_));
  INV_X1    g356(.A(new_n555_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n526_), .B1(new_n556_), .B2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT69), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT69), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n562_), .B(new_n526_), .C1(new_n556_), .C2(new_n559_), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n544_), .A2(new_n555_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT12), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n555_), .A2(KEYINPUT12), .A3(new_n542_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n557_), .A2(new_n558_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n567_), .A2(new_n525_), .A3(new_n568_), .A4(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n564_), .A2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G120gat), .B(G148gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G176gat), .B(G204gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n576_), .B(KEYINPUT71), .Z(new_n577_));
  NAND2_X1  g376(.A1(new_n571_), .A2(new_n577_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n561_), .A2(new_n576_), .A3(new_n563_), .A4(new_n570_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n523_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n577_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n581_), .B1(new_n564_), .B2(new_n570_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n579_), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n582_), .A2(KEYINPUT13), .A3(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n580_), .A2(new_n584_), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n481_), .A2(new_n522_), .A3(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(KEYINPUT73), .A2(KEYINPUT37), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n511_), .A2(new_n542_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT72), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT34), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n590_), .A2(KEYINPUT35), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n589_), .B1(new_n544_), .B2(new_n495_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n593_), .B(new_n589_), .C1(new_n495_), .C2(new_n544_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G190gat), .B(G218gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(G134gat), .ZN(new_n600_));
  INV_X1    g399(.A(G162gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT36), .ZN(new_n604_));
  INV_X1    g403(.A(new_n592_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT35), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n598_), .A2(new_n604_), .A3(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n603_), .A2(KEYINPUT36), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n609_), .ZN(new_n611_));
  AOI22_X1  g410(.A1(new_n596_), .A2(new_n597_), .B1(new_n606_), .B2(new_n605_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n611_), .B1(new_n612_), .B2(new_n604_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n588_), .B1(new_n610_), .B2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n608_), .A2(new_n609_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n612_), .A2(new_n611_), .A3(new_n604_), .ZN(new_n616_));
  XOR2_X1   g415(.A(KEYINPUT73), .B(KEYINPUT37), .Z(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n615_), .A2(new_n616_), .A3(new_n618_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n614_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(G231gat), .A2(G233gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n555_), .B(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(new_n488_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G127gat), .B(G155gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G183gat), .B(G211gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(KEYINPUT17), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n623_), .A2(new_n629_), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n628_), .B(KEYINPUT17), .Z(new_n631_));
  OAI21_X1  g430(.A(new_n630_), .B1(new_n623_), .B2(new_n631_), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n632_), .B(KEYINPUT76), .Z(new_n633_));
  NOR2_X1   g432(.A1(new_n620_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n586_), .A2(new_n634_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT103), .Z(new_n636_));
  INV_X1    g435(.A(G1gat), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n418_), .B(KEYINPUT104), .Z(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n636_), .A2(new_n637_), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT38), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n641_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n610_), .A2(new_n613_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n481_), .A2(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT105), .ZN(new_n646_));
  INV_X1    g445(.A(new_n633_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n585_), .A2(new_n522_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n646_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n418_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n642_), .B(new_n643_), .C1(new_n637_), .C2(new_n651_), .ZN(G1324gat));
  INV_X1    g451(.A(G8gat), .ZN(new_n653_));
  INV_X1    g452(.A(new_n348_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n636_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n646_), .A2(new_n647_), .A3(new_n654_), .A4(new_n648_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT39), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n656_), .A2(new_n657_), .A3(G8gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n656_), .B2(G8gat), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n655_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT40), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n655_), .B(KEYINPUT40), .C1(new_n658_), .C2(new_n659_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1325gat));
  OR3_X1    g463(.A1(new_n635_), .A2(G15gat), .A3(new_n445_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n649_), .A2(new_n446_), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n666_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(KEYINPUT41), .B1(new_n666_), .B2(G15gat), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n665_), .B1(new_n667_), .B2(new_n668_), .ZN(G1326gat));
  OR3_X1    g468(.A1(new_n635_), .A2(G22gat), .A3(new_n431_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n649_), .A2(new_n430_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT42), .ZN(new_n672_));
  AND3_X1   g471(.A1(new_n671_), .A2(new_n672_), .A3(G22gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n671_), .B2(G22gat), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n670_), .B1(new_n673_), .B2(new_n674_), .ZN(G1327gat));
  NOR3_X1   g474(.A1(new_n585_), .A2(new_n647_), .A3(new_n522_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n614_), .A2(KEYINPUT106), .A3(new_n619_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n677_), .A2(KEYINPUT43), .ZN(new_n678_));
  INV_X1    g477(.A(new_n620_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n481_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n677_), .A2(KEYINPUT43), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n474_), .A2(new_n479_), .A3(KEYINPUT102), .ZN(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT102), .B1(new_n474_), .B2(new_n479_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n447_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n681_), .B1(new_n684_), .B2(new_n620_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n676_), .B1(new_n680_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n676_), .B(KEYINPUT44), .C1(new_n680_), .C2(new_n685_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G29gat), .B1(new_n690_), .B2(new_n638_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n644_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n647_), .A2(new_n692_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n586_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(G29gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n694_), .A2(new_n695_), .A3(new_n650_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n691_), .A2(new_n696_), .ZN(G1328gat));
  NAND3_X1  g496(.A1(new_n688_), .A2(new_n654_), .A3(new_n689_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT107), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n688_), .A2(KEYINPUT107), .A3(new_n654_), .A4(new_n689_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n700_), .A2(G36gat), .A3(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(G36gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n694_), .A2(new_n703_), .A3(new_n654_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT45), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n702_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT108), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n707_), .A2(KEYINPUT46), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(new_n709_));
  OAI211_X1 g508(.A(new_n702_), .B(new_n705_), .C1(new_n707_), .C2(KEYINPUT46), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1329gat));
  NAND2_X1  g510(.A1(new_n446_), .A2(G43gat), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n694_), .A2(new_n446_), .ZN(new_n713_));
  OAI22_X1  g512(.A1(new_n690_), .A2(new_n712_), .B1(new_n713_), .B2(G43gat), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g514(.A(G50gat), .B1(new_n690_), .B2(new_n431_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n694_), .A2(new_n420_), .A3(new_n430_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1331gat));
  NOR2_X1   g517(.A1(new_n633_), .A2(new_n521_), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n646_), .A2(new_n585_), .A3(new_n719_), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n720_), .A2(G57gat), .A3(new_n650_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT109), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n722_), .B1(new_n481_), .B2(new_n521_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n684_), .A2(KEYINPUT109), .A3(new_n522_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n585_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(new_n634_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT110), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n638_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n730_), .B1(new_n729_), .B2(new_n728_), .ZN(new_n731_));
  INV_X1    g530(.A(G57gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n721_), .B1(new_n731_), .B2(new_n732_), .ZN(G1332gat));
  INV_X1    g532(.A(KEYINPUT48), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n720_), .A2(new_n654_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n735_), .B2(G64gat), .ZN(new_n736_));
  INV_X1    g535(.A(G64gat), .ZN(new_n737_));
  AOI211_X1 g536(.A(KEYINPUT48), .B(new_n737_), .C1(new_n720_), .C2(new_n654_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n654_), .A2(new_n737_), .ZN(new_n739_));
  OAI22_X1  g538(.A1(new_n736_), .A2(new_n738_), .B1(new_n728_), .B2(new_n739_), .ZN(G1333gat));
  NAND4_X1  g539(.A1(new_n727_), .A2(new_n549_), .A3(new_n446_), .A4(new_n634_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n646_), .A2(new_n446_), .A3(new_n585_), .A4(new_n719_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(KEYINPUT111), .B(KEYINPUT49), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n742_), .A2(G71gat), .A3(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n742_), .B2(G71gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n741_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT112), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n748_), .B(new_n741_), .C1(new_n744_), .C2(new_n745_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1334gat));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n720_), .A2(new_n430_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n752_), .B2(G78gat), .ZN(new_n753_));
  AOI211_X1 g552(.A(KEYINPUT50), .B(new_n550_), .C1(new_n720_), .C2(new_n430_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n430_), .A2(new_n550_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT113), .Z(new_n756_));
  OAI22_X1  g555(.A1(new_n753_), .A2(new_n754_), .B1(new_n728_), .B2(new_n756_), .ZN(G1335gat));
  INV_X1    g556(.A(new_n580_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n584_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n758_), .A2(new_n633_), .A3(new_n759_), .A4(new_n522_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT114), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT114), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n585_), .A2(new_n762_), .A3(new_n633_), .A4(new_n522_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n764_), .B1(new_n680_), .B2(new_n685_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT115), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  OR2_X1    g566(.A1(new_n680_), .A2(new_n685_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n768_), .A2(KEYINPUT115), .A3(new_n764_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n767_), .A2(new_n769_), .A3(G85gat), .A4(new_n650_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n725_), .A2(new_n585_), .A3(new_n693_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n771_), .A2(new_n638_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n770_), .B1(G85gat), .B2(new_n772_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT116), .ZN(G1336gat));
  INV_X1    g573(.A(new_n771_), .ZN(new_n775_));
  AOI21_X1  g574(.A(G92gat), .B1(new_n775_), .B2(new_n654_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n767_), .A2(new_n769_), .A3(new_n654_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(G92gat), .B2(new_n777_), .ZN(G1337gat));
  INV_X1    g577(.A(KEYINPUT117), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n779_), .A2(KEYINPUT51), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n767_), .A2(new_n769_), .A3(new_n446_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(G99gat), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n779_), .A2(KEYINPUT51), .ZN(new_n783_));
  NOR3_X1   g582(.A1(new_n771_), .A2(new_n445_), .A3(new_n540_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  AND4_X1   g584(.A1(new_n780_), .A2(new_n782_), .A3(new_n783_), .A4(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n784_), .B1(new_n781_), .B2(G99gat), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n780_), .B1(new_n787_), .B2(new_n783_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n786_), .A2(new_n788_), .ZN(G1338gat));
  NAND3_X1  g588(.A1(new_n768_), .A2(new_n430_), .A3(new_n764_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(G106gat), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(KEYINPUT118), .A3(new_n792_), .ZN(new_n793_));
  OR3_X1    g592(.A1(new_n771_), .A2(G106gat), .A3(new_n431_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(KEYINPUT118), .ZN(new_n795_));
  OR2_X1    g594(.A1(new_n792_), .A2(KEYINPUT118), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n790_), .A2(G106gat), .A3(new_n795_), .A4(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n793_), .A2(new_n794_), .A3(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT53), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n793_), .A2(new_n794_), .A3(new_n800_), .A4(new_n797_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n799_), .A2(new_n801_), .ZN(G1339gat));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n570_), .A2(new_n803_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n567_), .A2(KEYINPUT55), .A3(new_n568_), .A4(new_n569_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n525_), .A2(KEYINPUT119), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n556_), .B1(new_n566_), .B2(new_n565_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n806_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n808_), .A2(KEYINPUT55), .A3(new_n568_), .A4(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n804_), .A2(new_n807_), .A3(new_n810_), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n811_), .A2(KEYINPUT56), .A3(new_n577_), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT56), .B1(new_n811_), .B2(new_n577_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n501_), .A2(new_n502_), .A3(new_n506_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n512_), .A2(new_n503_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n814_), .A2(new_n517_), .A3(new_n815_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n520_), .A2(new_n816_), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n817_), .A2(KEYINPUT120), .A3(new_n579_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT120), .B1(new_n817_), .B2(new_n579_), .ZN(new_n819_));
  OAI22_X1  g618(.A1(new_n812_), .A2(new_n813_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n820_), .A2(KEYINPUT58), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT58), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n811_), .A2(new_n577_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT56), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n811_), .A2(KEYINPUT56), .A3(new_n577_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n817_), .A2(new_n579_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT120), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n817_), .A2(KEYINPUT120), .A3(new_n579_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n822_), .B1(new_n827_), .B2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n620_), .B1(new_n821_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT121), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n522_), .A2(new_n583_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n817_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT57), .B1(new_n840_), .B2(new_n692_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT57), .ZN(new_n842_));
  AOI211_X1 g641(.A(new_n842_), .B(new_n644_), .C1(new_n838_), .C2(new_n839_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n841_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n820_), .A2(KEYINPUT58), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n827_), .A2(new_n832_), .A3(new_n822_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n679_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT121), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n836_), .A2(new_n844_), .A3(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n633_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n620_), .A2(new_n633_), .A3(new_n521_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n758_), .A2(new_n759_), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n851_), .A2(new_n852_), .A3(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n852_), .B1(new_n851_), .B2(new_n853_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n850_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n348_), .A2(new_n446_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n430_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n639_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n858_), .A2(KEYINPUT122), .A3(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT122), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n856_), .B1(new_n849_), .B2(new_n633_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n861_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n863_), .A2(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(G113gat), .B1(new_n867_), .B2(new_n521_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n844_), .A2(new_n834_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT123), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n869_), .A2(new_n870_), .A3(new_n633_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n847_), .A2(new_n841_), .A3(new_n843_), .ZN(new_n872_));
  OAI21_X1  g671(.A(KEYINPUT123), .B1(new_n872_), .B2(new_n647_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n871_), .A2(new_n873_), .A3(new_n857_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n874_), .A2(new_n875_), .A3(new_n862_), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT59), .B1(new_n865_), .B2(new_n861_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n521_), .A2(G113gat), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(KEYINPUT124), .ZN(new_n879_));
  AND3_X1   g678(.A1(new_n876_), .A2(new_n877_), .A3(new_n879_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n868_), .A2(new_n880_), .ZN(G1340gat));
  XOR2_X1   g680(.A(KEYINPUT125), .B(G120gat), .Z(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n853_), .B2(KEYINPUT60), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n867_), .B(new_n884_), .C1(KEYINPUT60), .C2(new_n883_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n876_), .A2(new_n585_), .A3(new_n877_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n882_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n887_), .ZN(G1341gat));
  OAI21_X1  g687(.A(G127gat), .B1(new_n633_), .B2(KEYINPUT126), .ZN(new_n889_));
  OR2_X1    g688(.A1(KEYINPUT126), .A2(G127gat), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n876_), .A2(new_n877_), .A3(new_n889_), .A4(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n633_), .B1(new_n863_), .B2(new_n866_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(G127gat), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(G1342gat));
  XOR2_X1   g693(.A(KEYINPUT127), .B(G134gat), .Z(new_n895_));
  NAND4_X1  g694(.A1(new_n876_), .A2(new_n620_), .A3(new_n877_), .A4(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n692_), .B1(new_n863_), .B2(new_n866_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n897_), .B2(G134gat), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(G1343gat));
  NOR3_X1   g698(.A1(new_n638_), .A2(new_n431_), .A3(new_n446_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n858_), .A2(new_n348_), .A3(new_n900_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n901_), .A2(new_n522_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(new_n351_), .ZN(G1344gat));
  NOR2_X1   g702(.A1(new_n901_), .A2(new_n853_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(new_n352_), .ZN(G1345gat));
  NOR2_X1   g704(.A1(new_n901_), .A2(new_n633_), .ZN(new_n906_));
  XOR2_X1   g705(.A(KEYINPUT61), .B(G155gat), .Z(new_n907_));
  XNOR2_X1  g706(.A(new_n906_), .B(new_n907_), .ZN(G1346gat));
  NOR3_X1   g707(.A1(new_n901_), .A2(new_n601_), .A3(new_n679_), .ZN(new_n909_));
  OR2_X1    g708(.A1(new_n901_), .A2(new_n692_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(new_n601_), .B2(new_n910_), .ZN(G1347gat));
  NOR3_X1   g710(.A1(new_n639_), .A2(new_n348_), .A3(new_n445_), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n874_), .A2(new_n431_), .A3(new_n521_), .A4(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(G169gat), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT62), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  OR2_X1    g715(.A1(new_n913_), .A2(new_n269_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n913_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n916_), .A2(new_n917_), .A3(new_n918_), .ZN(G1348gat));
  NAND3_X1  g718(.A1(new_n585_), .A2(G176gat), .A3(new_n912_), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n865_), .A2(new_n430_), .A3(new_n920_), .ZN(new_n921_));
  AND2_X1   g720(.A1(new_n874_), .A2(new_n431_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n922_), .A2(new_n585_), .A3(new_n912_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n921_), .B1(new_n923_), .B2(new_n223_), .ZN(G1349gat));
  AND2_X1   g723(.A1(new_n912_), .A2(new_n647_), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n925_), .A2(new_n324_), .A3(new_n323_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n858_), .A2(new_n431_), .A3(new_n925_), .ZN(new_n927_));
  AOI22_X1  g726(.A1(new_n922_), .A2(new_n926_), .B1(new_n927_), .B2(new_n214_), .ZN(G1350gat));
  NAND4_X1  g727(.A1(new_n874_), .A2(new_n431_), .A3(new_n620_), .A4(new_n912_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(G190gat), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n922_), .A2(new_n257_), .A3(new_n912_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n930_), .B1(new_n931_), .B2(new_n692_), .ZN(G1351gat));
  NOR2_X1   g731(.A1(new_n865_), .A2(new_n650_), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n348_), .A2(new_n431_), .A3(new_n446_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n933_), .A2(new_n521_), .A3(new_n934_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g735(.A1(new_n933_), .A2(new_n585_), .A3(new_n934_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g737(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n933_), .A2(new_n934_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n939_), .B1(new_n940_), .B2(new_n633_), .ZN(new_n941_));
  XOR2_X1   g740(.A(KEYINPUT63), .B(G211gat), .Z(new_n942_));
  NAND4_X1  g741(.A1(new_n933_), .A2(new_n647_), .A3(new_n934_), .A4(new_n942_), .ZN(new_n943_));
  AND2_X1   g742(.A1(new_n941_), .A2(new_n943_), .ZN(G1354gat));
  INV_X1    g743(.A(G218gat), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n940_), .A2(new_n945_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n933_), .A2(new_n644_), .A3(new_n934_), .ZN(new_n947_));
  AOI22_X1  g746(.A1(new_n946_), .A2(new_n620_), .B1(new_n945_), .B2(new_n947_), .ZN(G1355gat));
endmodule


