//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n859_, new_n861_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n897_, new_n899_, new_n900_,
    new_n902_, new_n903_, new_n904_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n916_;
  XNOR2_X1  g000(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT88), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G141gat), .A2(G148gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT85), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT3), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT85), .B1(G141gat), .B2(G148gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT86), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT86), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n206_), .A2(new_n211_), .A3(new_n207_), .A4(new_n208_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G141gat), .A2(G148gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT84), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n216_));
  NAND3_X1  g015(.A1(KEYINPUT84), .A2(G141gat), .A3(G148gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n213_), .A2(new_n216_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n204_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n219_), .B1(KEYINPUT3), .B2(new_n220_), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n210_), .A2(new_n212_), .A3(new_n218_), .A4(new_n221_), .ZN(new_n222_));
  AND2_X1   g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n222_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT1), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n215_), .A2(new_n217_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n204_), .B1(new_n223_), .B2(KEYINPUT1), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n226_), .A2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n203_), .B1(new_n232_), .B2(KEYINPUT29), .ZN(new_n233_));
  INV_X1    g032(.A(new_n231_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n234_), .B1(new_n222_), .B2(new_n225_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT29), .ZN(new_n236_));
  INV_X1    g035(.A(new_n203_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n233_), .A2(new_n238_), .ZN(new_n239_));
  XOR2_X1   g038(.A(G22gat), .B(G50gat), .Z(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n233_), .A2(new_n240_), .A3(new_n238_), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  XOR2_X1   g043(.A(G211gat), .B(G218gat), .Z(new_n245_));
  INV_X1    g044(.A(KEYINPUT21), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G197gat), .B(G204gat), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n245_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(G197gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(KEYINPUT89), .A3(G204gat), .ZN(new_n250_));
  XOR2_X1   g049(.A(G197gat), .B(G204gat), .Z(new_n251_));
  OAI211_X1 g050(.A(KEYINPUT21), .B(new_n250_), .C1(new_n251_), .C2(KEYINPUT89), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n247_), .A2(new_n246_), .ZN(new_n253_));
  AOI22_X1  g052(.A1(new_n248_), .A2(new_n252_), .B1(new_n245_), .B2(new_n253_), .ZN(new_n254_));
  AND2_X1   g053(.A1(G228gat), .A2(G233gat), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n256_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT90), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n256_), .B(KEYINPUT90), .C1(new_n236_), .C2(new_n235_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n254_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT91), .B(KEYINPUT29), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n262_), .B1(new_n235_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(new_n255_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G78gat), .B(G106gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n261_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n267_), .B1(new_n261_), .B2(new_n265_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n244_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT92), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT92), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n272_), .B(new_n244_), .C1(new_n268_), .C2(new_n269_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n266_), .A2(KEYINPUT93), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n274_), .B1(new_n261_), .B2(new_n265_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n244_), .A2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n261_), .A2(new_n265_), .A3(new_n274_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n271_), .A2(new_n273_), .A3(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(G8gat), .B(G36gat), .Z(new_n280_));
  XNOR2_X1  g079(.A(G64gat), .B(G92gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT25), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n285_), .A2(KEYINPUT80), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n285_), .A2(KEYINPUT80), .ZN(new_n287_));
  OAI21_X1  g086(.A(G183gat), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT81), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT26), .B(G190gat), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n285_), .A2(G183gat), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT81), .ZN(new_n294_));
  OAI211_X1 g093(.A(new_n294_), .B(G183gat), .C1(new_n286_), .C2(new_n287_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n289_), .A2(new_n293_), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT82), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT23), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n297_), .A2(new_n298_), .A3(G183gat), .A4(G190gat), .ZN(new_n299_));
  INV_X1    g098(.A(G183gat), .ZN(new_n300_));
  INV_X1    g099(.A(G190gat), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT23), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n298_), .A2(G183gat), .A3(G190gat), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n302_), .A2(new_n303_), .A3(KEYINPUT82), .ZN(new_n304_));
  INV_X1    g103(.A(G169gat), .ZN(new_n305_));
  INV_X1    g104(.A(G176gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  OR2_X1    g106(.A1(new_n307_), .A2(KEYINPUT24), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(KEYINPUT24), .A3(new_n309_), .ZN(new_n310_));
  AND4_X1   g109(.A1(new_n299_), .A2(new_n304_), .A3(new_n308_), .A4(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n296_), .A2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n302_), .A2(new_n303_), .A3(KEYINPUT83), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n300_), .A2(new_n301_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT83), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n315_), .B(KEYINPUT23), .C1(new_n300_), .C2(new_n301_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n313_), .A2(new_n314_), .A3(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(G169gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n312_), .A2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT20), .B1(new_n321_), .B2(new_n262_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n304_), .A2(new_n314_), .A3(new_n299_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT97), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT97), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n304_), .A2(new_n325_), .A3(new_n314_), .A4(new_n299_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n309_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT22), .B(G169gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT96), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n328_), .B1(new_n330_), .B2(new_n306_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n327_), .A2(new_n331_), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n313_), .A2(new_n316_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT25), .B(G183gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n290_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT95), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n335_), .A2(new_n336_), .A3(new_n310_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n336_), .B1(new_n335_), .B2(new_n310_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n333_), .B(new_n308_), .C1(new_n337_), .C2(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n254_), .B1(new_n332_), .B2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G226gat), .A2(G233gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  NOR3_X1   g142(.A1(new_n322_), .A2(new_n340_), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n343_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT20), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n346_), .B1(new_n321_), .B2(new_n262_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n332_), .A2(new_n339_), .A3(new_n254_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n345_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n284_), .B1(new_n344_), .B2(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n343_), .B1(new_n322_), .B2(new_n340_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n284_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n347_), .A2(new_n348_), .A3(new_n345_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n350_), .A2(KEYINPUT27), .A3(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT101), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT27), .ZN(new_n357_));
  AND3_X1   g156(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n352_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n357_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT101), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n350_), .A2(new_n361_), .A3(KEYINPUT27), .A4(new_n354_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n356_), .A2(new_n360_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G225gat), .A2(G233gat), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT100), .ZN(new_n365_));
  XOR2_X1   g164(.A(G127gat), .B(G134gat), .Z(new_n366_));
  XOR2_X1   g165(.A(G113gat), .B(G120gat), .Z(new_n367_));
  XOR2_X1   g166(.A(new_n366_), .B(new_n367_), .Z(new_n368_));
  NAND3_X1  g167(.A1(new_n232_), .A2(new_n365_), .A3(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT4), .ZN(new_n370_));
  INV_X1    g169(.A(new_n368_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n370_), .B1(new_n235_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n369_), .A2(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n232_), .A2(new_n365_), .A3(new_n370_), .A4(new_n368_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n364_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G1gat), .B(G29gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(G85gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT0), .B(G57gat), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n377_), .B(new_n378_), .Z(new_n379_));
  NAND2_X1  g178(.A1(new_n232_), .A2(new_n368_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n235_), .A2(new_n371_), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n380_), .A2(new_n381_), .B1(G225gat), .B2(G233gat), .ZN(new_n382_));
  OR3_X1    g181(.A1(new_n375_), .A2(new_n379_), .A3(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n379_), .B1(new_n375_), .B2(new_n382_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  AOI22_X1  g184(.A1(new_n296_), .A2(new_n311_), .B1(new_n317_), .B2(new_n319_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G71gat), .B(G99gat), .ZN(new_n387_));
  INV_X1    g186(.A(G43gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n386_), .B(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n368_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n386_), .B(new_n389_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(new_n371_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G227gat), .A2(G233gat), .ZN(new_n395_));
  INV_X1    g194(.A(G15gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT30), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT31), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n392_), .A2(new_n394_), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n399_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NOR4_X1   g203(.A1(new_n279_), .A2(new_n363_), .A3(new_n385_), .A4(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n344_), .A2(new_n349_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n351_), .A2(new_n353_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n352_), .A2(KEYINPUT32), .ZN(new_n408_));
  MUX2_X1   g207(.A(new_n406_), .B(new_n407_), .S(new_n408_), .Z(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(new_n385_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT33), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n384_), .B(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT99), .B1(new_n358_), .B2(new_n359_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n407_), .A2(new_n284_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT99), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n415_), .A3(new_n354_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n373_), .A2(new_n364_), .A3(new_n374_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n379_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n380_), .A2(new_n381_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n417_), .B(new_n418_), .C1(new_n364_), .C2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n413_), .A2(new_n416_), .A3(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n410_), .B1(new_n412_), .B2(new_n421_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n271_), .A2(new_n273_), .A3(new_n278_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n356_), .A2(new_n360_), .A3(new_n362_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n385_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n279_), .A3(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n424_), .A2(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n405_), .B1(new_n428_), .B2(new_n404_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G113gat), .B(G141gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(KEYINPUT78), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G169gat), .B(G197gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(G22gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n396_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G15gat), .A2(G22gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G1gat), .A2(G8gat), .ZN(new_n437_));
  AOI22_X1  g236(.A1(new_n435_), .A2(new_n436_), .B1(KEYINPUT14), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  OR2_X1    g238(.A1(G1gat), .A2(G8gat), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT72), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(new_n441_), .A3(new_n437_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n441_), .B1(new_n440_), .B2(new_n437_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n439_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n444_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n446_), .A2(new_n438_), .A3(new_n442_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G29gat), .B(G36gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G43gat), .B(G50gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(G29gat), .B(G36gat), .Z(new_n451_));
  XOR2_X1   g250(.A(G43gat), .B(G50gat), .Z(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n445_), .A2(new_n447_), .B1(new_n450_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n450_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT15), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n453_), .A2(KEYINPUT15), .A3(new_n450_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n458_), .A2(new_n459_), .A3(new_n447_), .A4(new_n445_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G229gat), .A2(G233gat), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n455_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT77), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT77), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n455_), .A2(new_n460_), .A3(new_n464_), .A4(new_n461_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT76), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n445_), .A2(new_n447_), .A3(new_n450_), .A4(new_n453_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n467_), .B1(new_n469_), .B2(new_n454_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n455_), .A2(new_n468_), .A3(KEYINPUT76), .ZN(new_n471_));
  INV_X1    g270(.A(new_n461_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n470_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n433_), .B1(new_n466_), .B2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n470_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n433_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n475_), .A2(new_n463_), .A3(new_n465_), .A4(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n474_), .A2(KEYINPUT79), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT79), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n479_), .B(new_n433_), .C1(new_n466_), .C2(new_n473_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n429_), .A2(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(KEYINPUT73), .B(KEYINPUT16), .Z(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT74), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G127gat), .B(G155gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G183gat), .B(G211gat), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n486_), .B(new_n487_), .Z(new_n488_));
  INV_X1    g287(.A(KEYINPUT17), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G57gat), .B(G64gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT65), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n492_), .A2(KEYINPUT65), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT11), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G71gat), .B(G78gat), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n492_), .A2(KEYINPUT65), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT11), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n499_), .A2(new_n500_), .A3(new_n493_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n496_), .A2(new_n498_), .A3(new_n501_), .ZN(new_n502_));
  OAI211_X1 g301(.A(KEYINPUT11), .B(new_n497_), .C1(new_n494_), .C2(new_n495_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G231gat), .A2(G233gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n445_), .A2(new_n447_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n488_), .A2(new_n489_), .ZN(new_n509_));
  NOR3_X1   g308(.A1(new_n491_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n510_), .B1(new_n491_), .B2(new_n508_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G85gat), .A2(G92gat), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n512_), .A2(KEYINPUT9), .ZN(new_n513_));
  OR2_X1    g312(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n514_));
  INV_X1    g313(.A(G106gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n514_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  OR2_X1    g316(.A1(G85gat), .A2(G92gat), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n518_), .A2(KEYINPUT9), .A3(new_n512_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G99gat), .A2(G106gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT6), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT6), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n522_), .A2(G99gat), .A3(G106gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  AND4_X1   g323(.A1(new_n513_), .A2(new_n517_), .A3(new_n519_), .A4(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n518_), .A2(new_n512_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n521_), .A2(new_n523_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT7), .ZN(new_n529_));
  INV_X1    g328(.A(G99gat), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(new_n530_), .A3(new_n515_), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n527_), .B1(new_n528_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT8), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n522_), .B1(G99gat), .B2(G106gat), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n520_), .A2(KEYINPUT6), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n532_), .B(new_n531_), .C1(new_n536_), .C2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT8), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n538_), .A2(new_n539_), .A3(new_n527_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n525_), .B1(new_n535_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n458_), .A2(new_n459_), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT67), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n517_), .A2(new_n519_), .A3(new_n524_), .A4(new_n513_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n532_), .ZN(new_n545_));
  NOR3_X1   g344(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  AOI211_X1 g346(.A(KEYINPUT8), .B(new_n526_), .C1(new_n547_), .C2(new_n524_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n539_), .B1(new_n538_), .B2(new_n527_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n544_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT67), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n550_), .A2(new_n551_), .A3(new_n459_), .A4(new_n458_), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n543_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT68), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n550_), .A2(KEYINPUT64), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT64), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n556_), .B(new_n544_), .C1(new_n548_), .C2(new_n549_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(new_n456_), .A3(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G232gat), .A2(G233gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n553_), .A2(new_n554_), .A3(new_n558_), .A4(new_n562_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n558_), .A2(new_n543_), .A3(new_n554_), .A4(new_n552_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(new_n561_), .ZN(new_n565_));
  AOI21_X1  g364(.A(KEYINPUT35), .B1(new_n553_), .B2(new_n558_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n563_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G190gat), .B(G218gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT69), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G134gat), .B(G162gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT36), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n571_), .A2(new_n572_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n567_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n558_), .A2(new_n543_), .A3(new_n552_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT35), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n578_), .A2(new_n564_), .A3(new_n561_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n579_), .A2(new_n572_), .A3(new_n571_), .A4(new_n563_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT71), .ZN(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT70), .B(KEYINPUT37), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n575_), .A2(new_n580_), .A3(new_n581_), .A4(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n575_), .A2(new_n580_), .A3(new_n582_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT71), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT37), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n586_), .B1(new_n575_), .B2(new_n580_), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n511_), .B(new_n583_), .C1(new_n585_), .C2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G230gat), .A2(G233gat), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n555_), .A2(new_n557_), .A3(new_n504_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n504_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n590_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(G120gat), .B(G148gat), .Z(new_n594_));
  XNOR2_X1  g393(.A(KEYINPUT66), .B(KEYINPUT5), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G176gat), .B(G204gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n555_), .A2(new_n557_), .A3(new_n504_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n550_), .A2(new_n502_), .A3(KEYINPUT12), .A4(new_n503_), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n600_), .B(new_n601_), .C1(new_n592_), .C2(KEYINPUT12), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n593_), .B(new_n599_), .C1(new_n602_), .C2(new_n590_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n600_), .A2(new_n601_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n502_), .A2(new_n503_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n535_), .A2(new_n540_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n556_), .B1(new_n607_), .B2(new_n544_), .ZN(new_n608_));
  AOI211_X1 g407(.A(KEYINPUT64), .B(new_n525_), .C1(new_n535_), .C2(new_n540_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n606_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT12), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n605_), .A2(new_n612_), .A3(new_n589_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n599_), .B1(new_n613_), .B2(new_n593_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n604_), .A2(new_n614_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n615_), .A2(KEYINPUT13), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(KEYINPUT13), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n588_), .A2(new_n618_), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n619_), .A2(KEYINPUT75), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n482_), .A2(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n621_), .B1(KEYINPUT75), .B2(new_n619_), .ZN(new_n622_));
  INV_X1    g421(.A(G1gat), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(new_n623_), .A3(new_n385_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT103), .Z(new_n627_));
  NAND2_X1  g426(.A1(new_n624_), .A2(new_n625_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n575_), .A2(new_n580_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n429_), .A2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n618_), .A2(new_n481_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n631_), .A2(new_n511_), .A3(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G1gat), .B1(new_n633_), .B2(new_n426_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n627_), .A2(new_n628_), .A3(new_n634_), .ZN(G1324gat));
  OAI21_X1  g434(.A(G8gat), .B1(new_n633_), .B2(new_n425_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n636_), .A2(KEYINPUT104), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT39), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n636_), .A2(KEYINPUT104), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n425_), .A2(G8gat), .ZN(new_n642_));
  AOI22_X1  g441(.A1(new_n637_), .A2(new_n638_), .B1(new_n622_), .B2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT40), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(G1325gat));
  OAI21_X1  g445(.A(G15gat), .B1(new_n633_), .B2(new_n404_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n647_), .A2(new_n648_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n622_), .A2(new_n396_), .A3(new_n403_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n649_), .A2(new_n650_), .A3(new_n651_), .ZN(G1326gat));
  OAI21_X1  g451(.A(G22gat), .B1(new_n633_), .B2(new_n423_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT42), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n622_), .A2(new_n434_), .A3(new_n279_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1327gat));
  INV_X1    g455(.A(new_n618_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n511_), .A2(new_n629_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n482_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(G29gat), .B1(new_n660_), .B2(new_n385_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n583_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(KEYINPUT43), .B1(new_n429_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT43), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n403_), .B1(new_n424_), .B2(new_n427_), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n665_), .B(new_n662_), .C1(new_n666_), .C2(new_n405_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n664_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n511_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n632_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(KEYINPUT44), .B1(new_n668_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673_));
  AOI211_X1 g472(.A(new_n673_), .B(new_n670_), .C1(new_n664_), .C2(new_n667_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n672_), .A2(new_n674_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n385_), .A2(G29gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n661_), .B1(new_n675_), .B2(new_n676_), .ZN(G1328gat));
  INV_X1    g476(.A(new_n405_), .ZN(new_n678_));
  AOI22_X1  g477(.A1(new_n270_), .A2(KEYINPUT92), .B1(new_n276_), .B2(new_n277_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n385_), .B1(new_n679_), .B2(new_n273_), .ZN(new_n680_));
  AOI22_X1  g479(.A1(new_n680_), .A2(new_n425_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n678_), .B1(new_n681_), .B2(new_n403_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n665_), .B1(new_n682_), .B2(new_n662_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n667_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n671_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(new_n673_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n668_), .A2(KEYINPUT44), .A3(new_n671_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n686_), .A2(new_n363_), .A3(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n688_), .A2(KEYINPUT106), .A3(G36gat), .ZN(new_n689_));
  INV_X1    g488(.A(G36gat), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n363_), .A2(new_n690_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n659_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT45), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n692_), .B(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n689_), .A2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT106), .B1(new_n688_), .B2(G36gat), .ZN(new_n696_));
  OAI211_X1 g495(.A(KEYINPUT107), .B(KEYINPUT46), .C1(new_n695_), .C2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n672_), .A2(new_n674_), .A3(new_n425_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n699_), .B1(new_n700_), .B2(new_n690_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n701_), .A2(new_n689_), .A3(new_n694_), .ZN(new_n702_));
  AOI21_X1  g501(.A(KEYINPUT46), .B1(new_n702_), .B2(KEYINPUT107), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n698_), .A2(new_n703_), .ZN(G1329gat));
  AOI21_X1  g503(.A(G43gat), .B1(new_n660_), .B2(new_n403_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n404_), .A2(new_n388_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n675_), .B2(new_n706_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g507(.A(G50gat), .B1(new_n660_), .B2(new_n279_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n279_), .A2(G50gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n675_), .B2(new_n710_), .ZN(G1331gat));
  INV_X1    g510(.A(new_n481_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n429_), .A2(new_n657_), .A3(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(new_n663_), .A3(new_n511_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT108), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n426_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n717_));
  AOI21_X1  g516(.A(G57gat), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n657_), .A2(new_n712_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n631_), .A2(new_n511_), .A3(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT109), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n385_), .A2(G57gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n718_), .B1(new_n722_), .B2(new_n723_), .ZN(G1332gat));
  OAI21_X1  g523(.A(G64gat), .B1(new_n721_), .B2(new_n425_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT48), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n425_), .A2(G64gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n714_), .B2(new_n727_), .ZN(G1333gat));
  OR3_X1    g527(.A1(new_n714_), .A2(G71gat), .A3(new_n404_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G71gat), .B1(new_n721_), .B2(new_n404_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n730_), .A2(KEYINPUT49), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n730_), .A2(KEYINPUT49), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n729_), .B1(new_n731_), .B2(new_n732_), .ZN(G1334gat));
  OAI21_X1  g532(.A(G78gat), .B1(new_n721_), .B2(new_n423_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT50), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n423_), .A2(G78gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n735_), .B1(new_n714_), .B2(new_n736_), .ZN(G1335gat));
  NAND2_X1  g536(.A1(new_n713_), .A2(new_n658_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(G85gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(new_n740_), .A3(new_n385_), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n668_), .A2(new_n669_), .A3(new_n719_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n742_), .A2(new_n385_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n741_), .B1(new_n743_), .B2(new_n740_), .ZN(G1336gat));
  AOI21_X1  g543(.A(G92gat), .B1(new_n739_), .B2(new_n363_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n363_), .A2(G92gat), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT110), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n745_), .B1(new_n742_), .B2(new_n747_), .ZN(G1337gat));
  AOI21_X1  g547(.A(new_n530_), .B1(new_n742_), .B2(new_n403_), .ZN(new_n749_));
  AND4_X1   g548(.A1(new_n514_), .A2(new_n739_), .A3(new_n516_), .A4(new_n403_), .ZN(new_n750_));
  OAI22_X1  g549(.A1(new_n749_), .A2(new_n750_), .B1(KEYINPUT111), .B2(KEYINPUT51), .ZN(new_n751_));
  NAND2_X1  g550(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n752_), .B(KEYINPUT112), .Z(new_n753_));
  XNOR2_X1  g552(.A(new_n751_), .B(new_n753_), .ZN(G1338gat));
  NAND3_X1  g553(.A1(new_n739_), .A2(new_n515_), .A3(new_n279_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n515_), .B1(new_n742_), .B2(new_n279_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n756_), .A2(new_n757_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n755_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT53), .ZN(G1339gat));
  OR2_X1    g560(.A1(new_n588_), .A2(new_n618_), .ZN(new_n762_));
  AND2_X1   g561(.A1(KEYINPUT113), .A2(KEYINPUT54), .ZN(new_n763_));
  NOR2_X1   g562(.A1(KEYINPUT113), .A2(KEYINPUT54), .ZN(new_n764_));
  OAI22_X1  g563(.A1(new_n762_), .A2(new_n712_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  OR4_X1    g564(.A1(new_n588_), .A2(new_n618_), .A3(new_n712_), .A4(new_n763_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n470_), .A2(new_n471_), .A3(new_n461_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n455_), .A2(new_n460_), .A3(new_n472_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n768_), .A2(new_n433_), .A3(new_n769_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n477_), .A2(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n771_), .B1(new_n604_), .B2(new_n614_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT116), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  OAI211_X1 g573(.A(KEYINPUT116), .B(new_n771_), .C1(new_n604_), .C2(new_n614_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT55), .B1(new_n589_), .B2(KEYINPUT114), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n777_), .B1(KEYINPUT55), .B2(new_n589_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n605_), .A2(new_n612_), .A3(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n777_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n555_), .A2(new_n557_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT12), .B1(new_n782_), .B2(new_n606_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n600_), .A2(new_n601_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n781_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n780_), .A2(new_n785_), .A3(new_n598_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n786_), .A2(new_n787_), .A3(KEYINPUT56), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT56), .B1(new_n786_), .B2(new_n787_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n478_), .A2(new_n603_), .A3(new_n480_), .ZN(new_n790_));
  NOR3_X1   g589(.A1(new_n788_), .A2(new_n789_), .A3(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n629_), .B1(new_n776_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT57), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n771_), .A2(new_n603_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT56), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n786_), .A2(new_n796_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n780_), .A2(new_n785_), .A3(KEYINPUT56), .A4(new_n598_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n795_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT58), .B1(new_n799_), .B2(KEYINPUT117), .ZN(new_n800_));
  OR3_X1    g599(.A1(new_n799_), .A2(KEYINPUT117), .A3(KEYINPUT58), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n662_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(KEYINPUT57), .B(new_n629_), .C1(new_n776_), .C2(new_n791_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n794_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n669_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n767_), .A2(new_n805_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n279_), .A2(new_n363_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n807_), .A2(new_n385_), .A3(new_n403_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n806_), .A2(new_n809_), .A3(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(G113gat), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n481_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT118), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n804_), .A2(new_n814_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n794_), .A2(new_n802_), .A3(KEYINPUT118), .A4(new_n803_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n669_), .A3(new_n816_), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n817_), .A2(KEYINPUT119), .A3(new_n767_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT119), .B1(new_n817_), .B2(new_n767_), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n818_), .A2(new_n819_), .A3(new_n808_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT59), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n811_), .B(new_n813_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n817_), .A2(new_n767_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n817_), .A2(KEYINPUT119), .A3(new_n767_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n825_), .A2(new_n712_), .A3(new_n826_), .A4(new_n809_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT120), .ZN(new_n828_));
  AND3_X1   g627(.A1(new_n827_), .A2(new_n828_), .A3(new_n812_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n827_), .B2(new_n812_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n822_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT122), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT122), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n833_), .B(new_n822_), .C1(new_n829_), .C2(new_n830_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n834_), .ZN(G1340gat));
  NAND3_X1  g634(.A1(new_n825_), .A2(new_n826_), .A3(new_n809_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT59), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n837_), .A2(new_n618_), .A3(new_n811_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT124), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n837_), .A2(KEYINPUT124), .A3(new_n618_), .A4(new_n811_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(G120gat), .A3(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT60), .ZN(new_n843_));
  AOI21_X1  g642(.A(G120gat), .B1(new_n618_), .B2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT123), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT123), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n846_), .B1(new_n843_), .B2(G120gat), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n820_), .B(new_n845_), .C1(new_n844_), .C2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n842_), .A2(new_n848_), .ZN(G1341gat));
  NAND2_X1  g648(.A1(new_n837_), .A2(new_n811_), .ZN(new_n850_));
  OAI21_X1  g649(.A(G127gat), .B1(new_n850_), .B2(new_n669_), .ZN(new_n851_));
  OR3_X1    g650(.A1(new_n836_), .A2(G127gat), .A3(new_n669_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1342gat));
  OAI21_X1  g652(.A(G134gat), .B1(new_n850_), .B2(new_n663_), .ZN(new_n854_));
  OR3_X1    g653(.A1(new_n836_), .A2(G134gat), .A3(new_n629_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(G1343gat));
  NOR4_X1   g655(.A1(new_n423_), .A2(new_n426_), .A3(new_n363_), .A4(new_n403_), .ZN(new_n857_));
  AND3_X1   g656(.A1(new_n825_), .A2(new_n826_), .A3(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n712_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n618_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g661(.A1(new_n818_), .A2(new_n819_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n857_), .ZN(new_n864_));
  OAI21_X1  g663(.A(KEYINPUT125), .B1(new_n864_), .B2(new_n669_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT125), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n858_), .A2(new_n866_), .A3(new_n511_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n867_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(KEYINPUT61), .B(G155gat), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n870_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n865_), .A2(new_n867_), .A3(new_n869_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(G1346gat));
  OAI21_X1  g672(.A(G162gat), .B1(new_n864_), .B2(new_n663_), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n629_), .A2(G162gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n864_), .B2(new_n875_), .ZN(G1347gat));
  NOR2_X1   g675(.A1(new_n404_), .A2(new_n385_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n363_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n878_), .A2(new_n279_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n806_), .A2(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n305_), .B1(new_n880_), .B2(new_n712_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT126), .ZN(new_n882_));
  OR2_X1    g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n882_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT62), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n883_), .A2(KEYINPUT62), .A3(new_n884_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n880_), .A2(new_n330_), .A3(new_n712_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n887_), .A2(new_n888_), .A3(new_n889_), .ZN(G1348gat));
  AOI21_X1  g689(.A(G176gat), .B1(new_n880_), .B2(new_n618_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n818_), .A2(new_n819_), .A3(new_n279_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n657_), .A2(new_n306_), .A3(new_n878_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n891_), .B1(new_n892_), .B2(new_n893_), .ZN(G1349gat));
  INV_X1    g693(.A(new_n880_), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n895_), .A2(new_n669_), .A3(new_n334_), .ZN(new_n896_));
  NAND4_X1  g695(.A1(new_n892_), .A2(new_n511_), .A3(new_n363_), .A4(new_n877_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n896_), .B1(new_n897_), .B2(new_n300_), .ZN(G1350gat));
  OAI21_X1  g697(.A(G190gat), .B1(new_n895_), .B2(new_n663_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n880_), .A2(new_n630_), .A3(new_n290_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(G1351gat));
  NOR4_X1   g700(.A1(new_n423_), .A2(new_n425_), .A3(new_n385_), .A4(new_n403_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n863_), .A2(new_n902_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n903_), .A2(new_n481_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(new_n249_), .ZN(G1352gat));
  INV_X1    g704(.A(new_n903_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n618_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g707(.A1(new_n903_), .A2(new_n669_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n909_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n910_));
  XOR2_X1   g709(.A(KEYINPUT63), .B(G211gat), .Z(new_n911_));
  AOI21_X1  g710(.A(new_n910_), .B1(new_n909_), .B2(new_n911_), .ZN(G1354gat));
  AND3_X1   g711(.A1(new_n906_), .A2(G218gat), .A3(new_n662_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n903_), .A2(new_n629_), .ZN(new_n914_));
  OR2_X1    g713(.A1(new_n914_), .A2(KEYINPUT127), .ZN(new_n915_));
  AOI21_X1  g714(.A(G218gat), .B1(new_n914_), .B2(KEYINPUT127), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n913_), .B1(new_n915_), .B2(new_n916_), .ZN(G1355gat));
endmodule


