//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 0 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n640_, new_n641_, new_n642_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n841_, new_n842_, new_n843_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n874_, new_n875_, new_n876_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT90), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT2), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT2), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n208_), .A2(KEYINPUT90), .A3(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n210_), .B(new_n212_), .C1(new_n213_), .C2(new_n214_), .ZN(new_n215_));
  AND3_X1   g014(.A1(new_n214_), .A2(KEYINPUT89), .A3(new_n213_), .ZN(new_n216_));
  AOI21_X1  g015(.A(KEYINPUT89), .B1(new_n214_), .B2(new_n213_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n207_), .B1(new_n215_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT1), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n206_), .B1(new_n205_), .B2(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n221_), .B1(new_n220_), .B2(new_n205_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n214_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(new_n208_), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n219_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT29), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G211gat), .B(G218gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT92), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT21), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G197gat), .B(G204gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n227_), .A2(KEYINPUT21), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n234_), .A2(new_n232_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n233_), .B1(new_n231_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n226_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(G228gat), .ZN(new_n238_));
  INV_X1    g037(.A(G233gat), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n237_), .A2(new_n240_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n226_), .B(new_n236_), .C1(new_n238_), .C2(new_n239_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n203_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n241_), .A2(new_n242_), .A3(new_n203_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n225_), .A2(KEYINPUT29), .ZN(new_n247_));
  XOR2_X1   g046(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n248_));
  XNOR2_X1  g047(.A(G22gat), .B(G50gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n247_), .B(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n251_), .B1(new_n243_), .B2(KEYINPUT93), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n246_), .A2(new_n252_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n244_), .A2(new_n251_), .A3(KEYINPUT93), .A4(new_n245_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G227gat), .A2(G233gat), .ZN(new_n257_));
  INV_X1    g056(.A(G15gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT30), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT31), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT83), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G169gat), .A2(G176gat), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT81), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT22), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n264_), .B1(new_n265_), .B2(G169gat), .ZN(new_n266_));
  INV_X1    g065(.A(G176gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT82), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT82), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(G176gat), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n266_), .A2(new_n268_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(G169gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT22), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n265_), .A2(G169gat), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n264_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n262_), .B(new_n263_), .C1(new_n271_), .C2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT84), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G183gat), .A2(G190gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT23), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT23), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n280_), .A2(G183gat), .A3(G190gat), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n277_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT84), .B1(new_n278_), .B2(KEYINPUT23), .ZN(new_n283_));
  OAI22_X1  g082(.A1(new_n282_), .A2(new_n283_), .B1(G183gat), .B2(G190gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n276_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT82), .B(G176gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT22), .B(G169gat), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n266_), .B(new_n286_), .C1(new_n287_), .C2(new_n264_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n262_), .B1(new_n288_), .B2(new_n263_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n285_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(KEYINPUT79), .A2(G190gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT26), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT26), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(KEYINPUT79), .A3(G190gat), .ZN(new_n294_));
  INV_X1    g093(.A(G183gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT25), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT25), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(G183gat), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n292_), .A2(new_n294_), .A3(new_n296_), .A4(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT80), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n272_), .A2(new_n267_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(KEYINPUT24), .A3(new_n263_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n299_), .A2(new_n300_), .A3(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n300_), .B1(new_n299_), .B2(new_n302_), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n301_), .A2(KEYINPUT24), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n279_), .A2(new_n281_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NOR3_X1   g107(.A1(new_n304_), .A2(new_n305_), .A3(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT85), .B1(new_n290_), .B2(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n305_), .A2(new_n308_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n303_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n263_), .B1(new_n271_), .B2(new_n275_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT83), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(new_n284_), .A3(new_n276_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT85), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n312_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n310_), .A2(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(G71gat), .B(G99gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(G43gat), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n318_), .A2(new_n320_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT87), .ZN(new_n324_));
  INV_X1    g123(.A(G134gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(G127gat), .ZN(new_n326_));
  INV_X1    g125(.A(G127gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(G134gat), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n326_), .A2(new_n328_), .A3(KEYINPUT86), .ZN(new_n329_));
  AOI21_X1  g128(.A(KEYINPUT86), .B1(new_n326_), .B2(new_n328_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G113gat), .B(G120gat), .ZN(new_n331_));
  NOR3_X1   g130(.A1(new_n329_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n331_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n326_), .A2(new_n328_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT86), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n326_), .A2(new_n328_), .A3(KEYINPUT86), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n333_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n324_), .B1(new_n332_), .B2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n336_), .A2(new_n337_), .A3(new_n333_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(KEYINPUT87), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n323_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n323_), .A2(new_n343_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n261_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n346_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n261_), .ZN(new_n349_));
  NOR3_X1   g148(.A1(new_n348_), .A2(new_n349_), .A3(new_n344_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT98), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n225_), .A2(new_n339_), .A3(new_n341_), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n219_), .B(new_n224_), .C1(new_n332_), .C2(new_n338_), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n352_), .A2(KEYINPUT4), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT4), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n225_), .A2(new_n339_), .A3(new_n341_), .A4(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G225gat), .A2(G233gat), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n351_), .B1(new_n354_), .B2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n352_), .A2(KEYINPUT4), .A3(new_n353_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n361_), .A2(KEYINPUT98), .A3(new_n358_), .A4(new_n356_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n352_), .A2(new_n353_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n363_), .A2(new_n358_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n360_), .A2(new_n362_), .A3(new_n365_), .ZN(new_n366_));
  XOR2_X1   g165(.A(G1gat), .B(G29gat), .Z(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G57gat), .B(G85gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n366_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n371_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n360_), .A2(new_n373_), .A3(new_n365_), .A4(new_n362_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n347_), .A2(new_n350_), .A3(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G8gat), .B(G36gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT18), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G64gat), .B(G92gat), .ZN(new_n379_));
  XOR2_X1   g178(.A(new_n378_), .B(new_n379_), .Z(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n236_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n382_), .B1(new_n310_), .B2(new_n317_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(G226gat), .A2(G233gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT19), .ZN(new_n385_));
  INV_X1    g184(.A(new_n302_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT26), .B(G190gat), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT94), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n293_), .A2(G190gat), .ZN(new_n390_));
  INV_X1    g189(.A(G190gat), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n391_), .A2(KEYINPUT26), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT94), .B1(new_n390_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n389_), .A2(new_n393_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n296_), .A2(new_n298_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n386_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n306_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT95), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  OAI211_X1 g198(.A(KEYINPUT95), .B(new_n306_), .C1(new_n282_), .C2(new_n283_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n396_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n307_), .B1(G183gat), .B2(G190gat), .ZN(new_n402_));
  XOR2_X1   g201(.A(new_n263_), .B(KEYINPUT96), .Z(new_n403_));
  NAND2_X1  g202(.A1(new_n287_), .A2(new_n286_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n402_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n401_), .A2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT20), .B1(new_n406_), .B2(new_n236_), .ZN(new_n407_));
  NOR3_X1   g206(.A1(new_n383_), .A2(new_n385_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n385_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n310_), .A2(new_n382_), .A3(new_n317_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT20), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n411_), .B1(new_n406_), .B2(new_n236_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n409_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n381_), .B1(new_n408_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(new_n412_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n385_), .ZN(new_n416_));
  NOR3_X1   g215(.A1(new_n290_), .A2(new_n309_), .A3(KEYINPUT85), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n316_), .B1(new_n312_), .B2(new_n315_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n236_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n401_), .A2(new_n405_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n411_), .B1(new_n420_), .B2(new_n382_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n419_), .A2(new_n421_), .A3(new_n409_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n416_), .A2(new_n380_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT97), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n414_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT27), .ZN(new_n426_));
  OAI211_X1 g225(.A(KEYINPUT97), .B(new_n381_), .C1(new_n408_), .C2(new_n413_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n425_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT100), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n425_), .A2(KEYINPUT100), .A3(new_n426_), .A4(new_n427_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n415_), .A2(new_n385_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n409_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  OAI211_X1 g234(.A(KEYINPUT27), .B(new_n423_), .C1(new_n435_), .C2(new_n380_), .ZN(new_n436_));
  AND4_X1   g235(.A1(new_n256_), .A2(new_n376_), .A3(new_n432_), .A4(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT88), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n438_), .B1(new_n347_), .B2(new_n350_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n349_), .B1(new_n348_), .B2(new_n344_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n345_), .A2(new_n261_), .A3(new_n346_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(new_n441_), .A3(KEYINPUT88), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n439_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n375_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n444_), .A2(new_n436_), .A3(new_n255_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n445_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT33), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n374_), .A2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n361_), .A2(new_n358_), .A3(new_n356_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n364_), .B1(new_n449_), .B2(new_n351_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n450_), .A2(KEYINPUT33), .A3(new_n373_), .A4(new_n362_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n361_), .A2(new_n357_), .A3(new_n356_), .ZN(new_n452_));
  OAI211_X1 g251(.A(new_n452_), .B(new_n371_), .C1(new_n363_), .C2(new_n357_), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n448_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n425_), .A2(new_n427_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n380_), .A2(KEYINPUT32), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n416_), .A2(new_n457_), .A3(new_n422_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n375_), .B(new_n458_), .C1(new_n457_), .C2(new_n435_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n255_), .B1(new_n456_), .B2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n443_), .B1(new_n446_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT101), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT101), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n443_), .B(new_n463_), .C1(new_n446_), .C2(new_n460_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n437_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G29gat), .B(G36gat), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n466_), .A2(KEYINPUT72), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(KEYINPUT72), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G43gat), .B(G50gat), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n467_), .A2(new_n468_), .A3(new_n470_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G15gat), .B(G22gat), .ZN(new_n475_));
  INV_X1    g274(.A(G1gat), .ZN(new_n476_));
  INV_X1    g275(.A(G8gat), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT14), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n475_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G1gat), .B(G8gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n474_), .B(new_n481_), .ZN(new_n482_));
  OR2_X1    g281(.A1(new_n482_), .A2(KEYINPUT77), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(KEYINPUT77), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n483_), .A2(G229gat), .A3(G233gat), .A4(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n474_), .B(KEYINPUT15), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(new_n481_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n481_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n474_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G229gat), .A2(G233gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n490_), .B(KEYINPUT78), .Z(new_n491_));
  NAND3_X1  g290(.A1(new_n487_), .A2(new_n489_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n485_), .A2(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(G113gat), .B(G141gat), .Z(new_n494_));
  XNOR2_X1  g293(.A(G169gat), .B(G197gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  XOR2_X1   g295(.A(new_n493_), .B(new_n496_), .Z(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n465_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G57gat), .B(G64gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT11), .ZN(new_n501_));
  XOR2_X1   g300(.A(G71gat), .B(G78gat), .Z(new_n502_));
  OR2_X1    g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n500_), .A2(KEYINPUT11), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n501_), .A2(new_n502_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n503_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT68), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G85gat), .B(G92gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT67), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT66), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT8), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G99gat), .A2(G106gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT6), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n514_));
  OR3_X1    g313(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n513_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n509_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n511_), .A2(new_n517_), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n509_), .B(new_n516_), .C1(new_n510_), .C2(KEYINPUT8), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT65), .B(G85gat), .ZN(new_n521_));
  INV_X1    g320(.A(G92gat), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n520_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(KEYINPUT10), .B(G99gat), .Z(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n525_), .B(new_n513_), .C1(G106gat), .C2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n518_), .A2(new_n519_), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n507_), .A2(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G230gat), .A2(G233gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT64), .ZN(new_n535_));
  INV_X1    g334(.A(new_n529_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT68), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n506_), .B(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n506_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n529_), .A2(KEYINPUT12), .A3(new_n540_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n533_), .A2(new_n535_), .A3(new_n539_), .A4(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n539_), .A2(new_n530_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n535_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n542_), .A2(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(G120gat), .B(G148gat), .Z(new_n547_));
  XNOR2_X1  g346(.A(G176gat), .B(G204gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n546_), .B(new_n552_), .ZN(new_n553_));
  AND2_X1   g352(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n553_), .B1(new_n556_), .B2(new_n554_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  XOR2_X1   g357(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT75), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G127gat), .B(G155gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G183gat), .B(G211gat), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n562_), .B(new_n563_), .Z(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT17), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n481_), .B(new_n566_), .Z(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(new_n540_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n565_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n570_), .A2(KEYINPUT76), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n564_), .A2(KEYINPUT17), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n567_), .A2(new_n538_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n567_), .A2(new_n538_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n572_), .A2(new_n565_), .A3(new_n573_), .A4(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n570_), .A2(KEYINPUT76), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n571_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n536_), .A2(new_n474_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT73), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G232gat), .A2(G233gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT34), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT35), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n579_), .A2(new_n580_), .A3(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n583_), .A2(new_n584_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n486_), .A2(new_n529_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n588_), .A2(new_n585_), .A3(new_n579_), .A4(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G190gat), .B(G218gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G134gat), .B(G162gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n593_), .A2(KEYINPUT36), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n579_), .A2(new_n585_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n589_), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n586_), .B(new_n587_), .C1(new_n595_), .C2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n590_), .A2(new_n594_), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n593_), .B(KEYINPUT36), .Z(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n601_), .B1(new_n590_), .B2(new_n597_), .ZN(new_n602_));
  OAI21_X1  g401(.A(KEYINPUT37), .B1(new_n599_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n602_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT37), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n604_), .A2(new_n605_), .A3(new_n598_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n603_), .A2(new_n606_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n499_), .A2(new_n558_), .A3(new_n578_), .A4(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT102), .Z(new_n609_));
  NAND3_X1  g408(.A1(new_n609_), .A2(new_n476_), .A3(new_n375_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT38), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n558_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n613_), .A2(new_n498_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(new_n578_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT103), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n599_), .A2(new_n602_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n465_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  OAI21_X1  g418(.A(G1gat), .B1(new_n619_), .B2(new_n444_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n610_), .A2(new_n611_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n612_), .A2(new_n620_), .A3(new_n621_), .ZN(G1324gat));
  NAND2_X1  g421(.A1(new_n432_), .A2(new_n436_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n609_), .A2(new_n477_), .A3(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n619_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(new_n623_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n626_), .A2(G8gat), .A3(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n627_), .B1(new_n626_), .B2(G8gat), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n624_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT40), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n624_), .B(KEYINPUT40), .C1(new_n629_), .C2(new_n628_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(G1325gat));
  OAI21_X1  g433(.A(G15gat), .B1(new_n619_), .B2(new_n443_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT41), .Z(new_n636_));
  INV_X1    g435(.A(new_n443_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(new_n258_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n636_), .B1(new_n608_), .B2(new_n638_), .ZN(G1326gat));
  OAI21_X1  g438(.A(G22gat), .B1(new_n619_), .B2(new_n256_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT42), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n256_), .A2(G22gat), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n641_), .B1(new_n608_), .B2(new_n642_), .ZN(G1327gat));
  INV_X1    g442(.A(new_n617_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n644_), .A2(new_n578_), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n499_), .A2(new_n558_), .A3(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(G29gat), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n646_), .A2(new_n647_), .A3(new_n375_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n607_), .B(KEYINPUT105), .Z(new_n649_));
  OAI21_X1  g448(.A(KEYINPUT43), .B1(new_n465_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n437_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n445_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n432_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n456_), .A2(new_n459_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(new_n256_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n463_), .B1(new_n656_), .B2(new_n443_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n464_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n651_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n607_), .A2(KEYINPUT43), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n650_), .A2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n614_), .A2(new_n577_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n663_), .B1(new_n650_), .B2(new_n661_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(KEYINPUT44), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n667_), .A2(new_n375_), .A3(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n670_), .A2(KEYINPUT106), .A3(G29gat), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT106), .B1(new_n670_), .B2(G29gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n648_), .B1(new_n672_), .B2(new_n673_), .ZN(G1328gat));
  INV_X1    g473(.A(G36gat), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n646_), .A2(new_n675_), .A3(new_n623_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT45), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n667_), .A2(new_n623_), .A3(new_n669_), .ZN(new_n678_));
  AOI21_X1  g477(.A(KEYINPUT107), .B1(new_n678_), .B2(G36gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n623_), .B1(new_n668_), .B2(KEYINPUT44), .ZN(new_n680_));
  AOI211_X1 g479(.A(new_n666_), .B(new_n663_), .C1(new_n650_), .C2(new_n661_), .ZN(new_n681_));
  OAI211_X1 g480(.A(KEYINPUT107), .B(G36gat), .C1(new_n680_), .C2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n677_), .B1(new_n679_), .B2(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n677_), .B(new_n685_), .C1(new_n679_), .C2(new_n683_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1329gat));
  NOR2_X1   g488(.A1(new_n347_), .A2(new_n350_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n667_), .A2(G43gat), .A3(new_n690_), .A4(new_n669_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n646_), .A2(new_n637_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n691_), .B1(G43gat), .B2(new_n692_), .ZN(new_n693_));
  XOR2_X1   g492(.A(KEYINPUT109), .B(KEYINPUT47), .Z(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(G1330gat));
  AOI21_X1  g494(.A(G50gat), .B1(new_n646_), .B2(new_n255_), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n667_), .A2(G50gat), .A3(new_n255_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n697_), .B2(new_n669_), .ZN(G1331gat));
  NOR2_X1   g497(.A1(new_n465_), .A2(new_n497_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n699_), .A2(new_n613_), .A3(new_n578_), .A4(new_n607_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT110), .ZN(new_n701_));
  AOI21_X1  g500(.A(G57gat), .B1(new_n701_), .B2(new_n375_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n618_), .A2(new_n498_), .A3(new_n613_), .A4(new_n578_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT111), .ZN(new_n704_));
  INV_X1    g503(.A(G57gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(new_n375_), .B2(KEYINPUT112), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(KEYINPUT112), .B2(new_n705_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n702_), .B1(new_n704_), .B2(new_n707_), .ZN(G1332gat));
  INV_X1    g507(.A(G64gat), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n701_), .A2(new_n709_), .A3(new_n623_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n704_), .A2(new_n623_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(G64gat), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n712_), .A2(KEYINPUT48), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n712_), .A2(KEYINPUT48), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n710_), .B1(new_n713_), .B2(new_n714_), .ZN(G1333gat));
  NOR2_X1   g514(.A1(new_n443_), .A2(G71gat), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT114), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n701_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n704_), .A2(new_n637_), .ZN(new_n719_));
  XOR2_X1   g518(.A(KEYINPUT113), .B(KEYINPUT49), .Z(new_n720_));
  AND3_X1   g519(.A1(new_n719_), .A2(G71gat), .A3(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n719_), .B2(G71gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n718_), .B1(new_n721_), .B2(new_n722_), .ZN(G1334gat));
  INV_X1    g522(.A(G78gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n701_), .A2(new_n724_), .A3(new_n255_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n704_), .A2(new_n255_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(G78gat), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n727_), .A2(KEYINPUT50), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n727_), .A2(KEYINPUT50), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(G1335gat));
  AND3_X1   g529(.A1(new_n699_), .A2(new_n613_), .A3(new_n645_), .ZN(new_n731_));
  AOI21_X1  g530(.A(G85gat), .B1(new_n731_), .B2(new_n375_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n613_), .A2(new_n498_), .A3(new_n577_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n650_), .B2(new_n661_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT115), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n444_), .A2(new_n521_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n732_), .B1(new_n735_), .B2(new_n736_), .ZN(G1336gat));
  NAND3_X1  g536(.A1(new_n731_), .A2(new_n522_), .A3(new_n623_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n735_), .A2(new_n623_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(new_n522_), .ZN(G1337gat));
  NAND2_X1  g539(.A1(new_n734_), .A2(new_n637_), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n347_), .A2(new_n350_), .A3(new_n527_), .ZN(new_n742_));
  AOI22_X1  g541(.A1(new_n741_), .A2(G99gat), .B1(new_n731_), .B2(new_n742_), .ZN(new_n743_));
  XOR2_X1   g542(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n744_));
  XNOR2_X1  g543(.A(new_n743_), .B(new_n744_), .ZN(G1338gat));
  INV_X1    g544(.A(G106gat), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n731_), .A2(new_n746_), .A3(new_n255_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n734_), .A2(new_n255_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n749_), .B2(G106gat), .ZN(new_n750_));
  AOI211_X1 g549(.A(KEYINPUT52), .B(new_n746_), .C1(new_n734_), .C2(new_n255_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n747_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g552(.A(KEYINPUT118), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n539_), .A2(new_n541_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n531_), .B1(new_n507_), .B2(new_n529_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n544_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT55), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n542_), .B2(new_n758_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n542_), .A2(new_n758_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n552_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT56), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n546_), .A2(new_n552_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n485_), .A2(new_n492_), .A3(new_n496_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n487_), .A2(new_n489_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT117), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n491_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n768_), .B1(new_n767_), .B2(new_n766_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n483_), .A2(new_n484_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n496_), .B1(new_n770_), .B2(new_n491_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n765_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT56), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n773_), .B(new_n552_), .C1(new_n759_), .C2(new_n760_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n762_), .A2(new_n764_), .A3(new_n772_), .A4(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT58), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n763_), .B1(new_n761_), .B2(KEYINPUT56), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT58), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n777_), .A2(new_n778_), .A3(new_n772_), .A4(new_n774_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n776_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n607_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n754_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n777_), .A2(new_n497_), .A3(new_n774_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n772_), .A2(new_n553_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT57), .B1(new_n785_), .B2(new_n644_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT57), .ZN(new_n787_));
  AOI211_X1 g586(.A(new_n787_), .B(new_n617_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n782_), .A2(new_n786_), .A3(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n780_), .A2(new_n781_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n790_), .A2(KEYINPUT118), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n578_), .B1(new_n789_), .B2(new_n792_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n558_), .A2(new_n607_), .A3(new_n498_), .A4(new_n578_), .ZN(new_n794_));
  XOR2_X1   g593(.A(new_n794_), .B(KEYINPUT54), .Z(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT119), .B1(new_n793_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n782_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n786_), .A2(new_n788_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n577_), .B1(new_n799_), .B2(new_n791_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT119), .ZN(new_n801_));
  INV_X1    g600(.A(new_n795_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n800_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n623_), .ZN(new_n804_));
  AND4_X1   g603(.A1(new_n256_), .A2(new_n804_), .A3(new_n375_), .A4(new_n690_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n796_), .A2(new_n803_), .A3(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(G113gat), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n808_), .A3(new_n497_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n798_), .A2(new_n790_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n795_), .B1(new_n577_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT59), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n805_), .A2(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n811_), .A2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n814_), .B1(new_n806_), .B2(KEYINPUT59), .ZN(new_n815_));
  AND2_X1   g614(.A1(new_n815_), .A2(new_n497_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n809_), .B1(new_n816_), .B2(new_n808_), .ZN(G1340gat));
  INV_X1    g616(.A(G120gat), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n818_), .B1(new_n815_), .B2(new_n613_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n818_), .B1(new_n558_), .B2(KEYINPUT60), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n820_), .B1(KEYINPUT60), .B2(new_n818_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n806_), .A2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT120), .B1(new_n819_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT120), .ZN(new_n824_));
  INV_X1    g623(.A(new_n822_), .ZN(new_n825_));
  AOI211_X1 g624(.A(new_n558_), .B(new_n814_), .C1(new_n806_), .C2(KEYINPUT59), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n824_), .B(new_n825_), .C1(new_n826_), .C2(new_n818_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n823_), .A2(new_n827_), .ZN(G1341gat));
  AOI21_X1  g627(.A(G127gat), .B1(new_n807_), .B2(new_n578_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n327_), .B1(new_n578_), .B2(KEYINPUT121), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n830_), .B1(KEYINPUT121), .B2(new_n327_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n829_), .B1(new_n815_), .B2(new_n831_), .ZN(G1342gat));
  NAND3_X1  g631(.A1(new_n807_), .A2(new_n325_), .A3(new_n617_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n815_), .A2(new_n781_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n833_), .B1(new_n834_), .B2(new_n325_), .ZN(G1343gat));
  AND2_X1   g634(.A1(new_n796_), .A2(new_n803_), .ZN(new_n836_));
  NOR4_X1   g635(.A1(new_n637_), .A2(new_n623_), .A3(new_n256_), .A4(new_n444_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n497_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g639(.A1(new_n836_), .A2(new_n837_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n841_), .A2(new_n558_), .ZN(new_n842_));
  XOR2_X1   g641(.A(KEYINPUT122), .B(G148gat), .Z(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(G1345gat));
  NAND2_X1  g643(.A1(new_n838_), .A2(new_n578_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(KEYINPUT61), .B(G155gat), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n845_), .B(new_n846_), .ZN(G1346gat));
  AOI21_X1  g646(.A(G162gat), .B1(new_n838_), .B2(new_n617_), .ZN(new_n848_));
  INV_X1    g647(.A(G162gat), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n841_), .A2(new_n849_), .A3(new_n649_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n848_), .A2(new_n850_), .ZN(G1347gat));
  INV_X1    g650(.A(KEYINPUT62), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n804_), .A2(new_n375_), .A3(new_n443_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(new_n255_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n811_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n497_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n852_), .B1(new_n858_), .B2(G169gat), .ZN(new_n859_));
  AOI211_X1 g658(.A(KEYINPUT62), .B(new_n272_), .C1(new_n857_), .C2(new_n497_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n857_), .A2(new_n861_), .ZN(new_n862_));
  NOR3_X1   g661(.A1(new_n811_), .A2(KEYINPUT123), .A3(new_n856_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n497_), .A2(new_n287_), .ZN(new_n865_));
  OAI22_X1  g664(.A1(new_n859_), .A2(new_n860_), .B1(new_n864_), .B2(new_n865_), .ZN(G1348gat));
  AND2_X1   g665(.A1(new_n836_), .A2(new_n256_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n854_), .A2(new_n267_), .A3(new_n558_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n613_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n869_));
  AOI22_X1  g668(.A1(new_n867_), .A2(new_n868_), .B1(new_n869_), .B2(new_n286_), .ZN(G1349gat));
  NOR3_X1   g669(.A1(new_n864_), .A2(new_n395_), .A3(new_n577_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n867_), .A2(new_n578_), .A3(new_n853_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n871_), .B1(new_n295_), .B2(new_n872_), .ZN(G1350gat));
  OAI21_X1  g672(.A(G190gat), .B1(new_n864_), .B2(new_n607_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n617_), .A2(new_n394_), .ZN(new_n875_));
  XOR2_X1   g674(.A(new_n875_), .B(KEYINPUT124), .Z(new_n876_));
  OAI21_X1  g675(.A(new_n874_), .B1(new_n864_), .B2(new_n876_), .ZN(G1351gat));
  NOR4_X1   g676(.A1(new_n804_), .A2(new_n637_), .A3(new_n256_), .A4(new_n375_), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n796_), .A2(new_n803_), .A3(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n497_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n613_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g682(.A(KEYINPUT125), .ZN(new_n884_));
  XOR2_X1   g683(.A(KEYINPUT63), .B(G211gat), .Z(new_n885_));
  NAND4_X1  g684(.A1(new_n879_), .A2(new_n884_), .A3(new_n578_), .A4(new_n885_), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n796_), .A2(new_n803_), .A3(new_n578_), .A4(new_n878_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n885_), .ZN(new_n890_));
  OAI21_X1  g689(.A(KEYINPUT125), .B1(new_n887_), .B2(new_n890_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n886_), .A2(new_n889_), .A3(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT126), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n886_), .A2(new_n891_), .A3(KEYINPUT126), .A4(new_n889_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1354gat));
  NAND2_X1  g695(.A1(new_n879_), .A2(new_n617_), .ZN(new_n897_));
  XOR2_X1   g696(.A(KEYINPUT127), .B(G218gat), .Z(new_n898_));
  NOR2_X1   g697(.A1(new_n607_), .A2(new_n898_), .ZN(new_n899_));
  AOI22_X1  g698(.A1(new_n897_), .A2(new_n898_), .B1(new_n879_), .B2(new_n899_), .ZN(G1355gat));
endmodule


