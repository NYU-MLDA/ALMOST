//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 0 1 0 1 1 1 1 0 0 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n682_,
    new_n683_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n861_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n926_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT15), .ZN(new_n205_));
  OR2_X1    g004(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n206_));
  NAND2_X1  g005(.A1(KEYINPUT64), .A2(KEYINPUT9), .ZN(new_n207_));
  NAND4_X1  g006(.A1(new_n206_), .A2(G85gat), .A3(G92gat), .A4(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G85gat), .ZN(new_n209_));
  INV_X1    g008(.A(G92gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G85gat), .A2(G92gat), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n211_), .A2(KEYINPUT64), .A3(KEYINPUT9), .A4(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT6), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n216_), .A2(G99gat), .A3(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  OR2_X1    g017(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n219_));
  INV_X1    g018(.A(G106gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n208_), .A2(new_n213_), .A3(new_n218_), .A4(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n211_), .A2(new_n212_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NOR3_X1   g025(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  AOI211_X1 g027(.A(KEYINPUT8), .B(new_n224_), .C1(new_n228_), .C2(new_n218_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT8), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT7), .ZN(new_n231_));
  INV_X1    g030(.A(G99gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(new_n232_), .A3(new_n220_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n216_), .B1(G99gat), .B2(G106gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n225_), .B(new_n233_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n224_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n230_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n223_), .B1(new_n229_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n205_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT70), .ZN(new_n241_));
  INV_X1    g040(.A(new_n223_), .ZN(new_n242_));
  AND2_X1   g041(.A1(new_n215_), .A2(new_n217_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n233_), .A2(new_n225_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n237_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT8), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n236_), .A2(new_n230_), .A3(new_n237_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n242_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT35), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G232gat), .A2(G233gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT34), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  AOI22_X1  g051(.A1(new_n248_), .A2(new_n204_), .B1(new_n249_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n205_), .A2(new_n254_), .A3(new_n239_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n241_), .A2(new_n253_), .A3(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n252_), .A2(new_n249_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(KEYINPUT71), .A3(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(KEYINPUT71), .B1(new_n256_), .B2(new_n257_), .ZN(new_n260_));
  OR2_X1    g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT73), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G190gat), .B(G218gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G134gat), .B(G162gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n265_), .A2(KEYINPUT36), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n257_), .B(KEYINPUT72), .Z(new_n267_));
  NAND3_X1  g066(.A1(new_n253_), .A2(new_n240_), .A3(new_n267_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n261_), .A2(new_n262_), .A3(new_n266_), .A4(new_n268_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n266_), .B(new_n268_), .C1(new_n259_), .C2(new_n260_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT73), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n268_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n265_), .B(KEYINPUT36), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT74), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n269_), .A2(new_n271_), .A3(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT37), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(KEYINPUT75), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT37), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT75), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n272_), .A2(new_n280_), .A3(new_n274_), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n278_), .A2(new_n279_), .A3(new_n270_), .A4(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n277_), .A2(new_n282_), .ZN(new_n283_));
  XOR2_X1   g082(.A(G127gat), .B(G155gat), .Z(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT16), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G183gat), .B(G211gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT17), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n287_), .A2(new_n288_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G57gat), .B(G64gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT11), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT65), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT11), .ZN(new_n295_));
  INV_X1    g094(.A(G57gat), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n296_), .A2(G64gat), .ZN(new_n297_));
  INV_X1    g096(.A(G64gat), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n298_), .A2(G57gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n295_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(G71gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(G78gat), .ZN(new_n302_));
  INV_X1    g101(.A(G78gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(G71gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n294_), .B1(new_n300_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n298_), .A2(G57gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n296_), .A2(G64gat), .ZN(new_n308_));
  AOI21_X1  g107(.A(KEYINPUT11), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G71gat), .B(G78gat), .ZN(new_n310_));
  NOR3_X1   g109(.A1(new_n309_), .A2(KEYINPUT65), .A3(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n293_), .B1(new_n306_), .B2(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT65), .B1(new_n309_), .B2(new_n310_), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n305_), .B(new_n294_), .C1(new_n292_), .C2(KEYINPUT11), .ZN(new_n314_));
  INV_X1    g113(.A(new_n293_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n312_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G231gat), .A2(G233gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT76), .B(G15gat), .ZN(new_n320_));
  INV_X1    g119(.A(G22gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(KEYINPUT77), .B(G1gat), .Z(new_n323_));
  INV_X1    g122(.A(G8gat), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT14), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n322_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G1gat), .B(G8gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n319_), .B(new_n328_), .ZN(new_n329_));
  MUX2_X1   g128(.A(new_n291_), .B(new_n290_), .S(new_n329_), .Z(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT78), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n283_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT79), .ZN(new_n334_));
  XOR2_X1   g133(.A(G211gat), .B(G218gat), .Z(new_n335_));
  INV_X1    g134(.A(KEYINPUT21), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G197gat), .B(G204gat), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n335_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n337_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n340_), .A2(new_n335_), .A3(KEYINPUT21), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT87), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT86), .ZN(new_n347_));
  AND2_X1   g146(.A1(G141gat), .A2(G148gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT2), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT3), .ZN(new_n350_));
  OR2_X1    g149(.A1(new_n350_), .A2(KEYINPUT85), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(KEYINPUT85), .ZN(new_n352_));
  NOR2_X1   g151(.A1(G141gat), .A2(G148gat), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n345_), .A2(new_n347_), .A3(new_n349_), .A4(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G155gat), .A2(G162gat), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(G155gat), .A2(G162gat), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n355_), .A2(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n358_), .B1(KEYINPUT1), .B2(new_n356_), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n356_), .A2(KEYINPUT1), .ZN(new_n362_));
  AOI211_X1 g161(.A(new_n348_), .B(new_n353_), .C1(new_n361_), .C2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n360_), .A2(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n342_), .B1(new_n365_), .B2(KEYINPUT29), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G228gat), .A2(G233gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT88), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G78gat), .B(G106gat), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n368_), .A2(new_n369_), .A3(new_n371_), .ZN(new_n372_));
  OR3_X1    g171(.A1(new_n365_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT28), .B1(new_n365_), .B2(KEYINPUT29), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G22gat), .B(G50gat), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n373_), .A2(new_n374_), .A3(new_n376_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n370_), .B(KEYINPUT88), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n372_), .B(new_n380_), .C1(new_n368_), .C2(new_n381_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n371_), .A2(KEYINPUT89), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n368_), .A2(new_n383_), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n366_), .A2(new_n367_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n366_), .A2(new_n367_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n385_), .B(new_n386_), .C1(KEYINPUT89), .C2(new_n371_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n384_), .A2(new_n387_), .A3(new_n379_), .A4(new_n378_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n382_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT4), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G127gat), .B(G134gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(G113gat), .B(G120gat), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT84), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n392_), .B(new_n393_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT84), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n395_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n365_), .A2(new_n391_), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT92), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT92), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n365_), .A2(new_n401_), .A3(new_n391_), .A4(new_n398_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G225gat), .A2(G233gat), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n398_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n363_), .B1(new_n355_), .B2(new_n359_), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT91), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT91), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n365_), .A2(new_n409_), .A3(new_n398_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n407_), .A2(new_n396_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n408_), .A2(new_n410_), .A3(KEYINPUT4), .A4(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n403_), .A2(new_n405_), .A3(new_n412_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n408_), .A2(new_n410_), .A3(new_n404_), .A4(new_n411_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G1gat), .B(G29gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(G85gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT0), .B(G57gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n413_), .A2(new_n414_), .A3(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT93), .B(KEYINPUT33), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(KEYINPUT94), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n413_), .A2(KEYINPUT33), .A3(new_n414_), .A4(new_n419_), .ZN(new_n424_));
  INV_X1    g223(.A(G169gat), .ZN(new_n425_));
  INV_X1    g224(.A(G176gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G169gat), .A2(G176gat), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n427_), .A2(KEYINPUT24), .A3(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT81), .ZN(new_n430_));
  INV_X1    g229(.A(G183gat), .ZN(new_n431_));
  INV_X1    g230(.A(G190gat), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT23), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT82), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT82), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n435_), .B(KEYINPUT23), .C1(new_n431_), .C2(new_n432_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT23), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n438_), .A2(G183gat), .A3(G190gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n427_), .A2(KEYINPUT24), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT80), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT26), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n442_), .B1(new_n443_), .B2(G190gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT25), .B(G183gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT26), .B(G190gat), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n444_), .B(new_n445_), .C1(new_n446_), .C2(new_n442_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n430_), .A2(new_n440_), .A3(new_n441_), .A4(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(G169gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n433_), .A2(new_n439_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(G183gat), .A2(G190gat), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n450_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n448_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT83), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT83), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n448_), .A2(new_n457_), .A3(new_n454_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n339_), .A2(new_n341_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G226gat), .A2(G233gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT19), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n446_), .A2(new_n445_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n465_), .A2(new_n451_), .A3(new_n441_), .A4(new_n429_), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n466_), .A2(KEYINPUT90), .ZN(new_n467_));
  INV_X1    g266(.A(new_n439_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n468_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n450_), .B1(new_n469_), .B2(new_n453_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n466_), .A2(KEYINPUT90), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n467_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  OAI211_X1 g271(.A(KEYINPUT20), .B(new_n464_), .C1(new_n472_), .C2(new_n460_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n461_), .A2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G8gat), .B(G36gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT18), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G64gat), .B(G92gat), .ZN(new_n478_));
  XOR2_X1   g277(.A(new_n477_), .B(new_n478_), .Z(new_n479_));
  NAND3_X1  g278(.A1(new_n456_), .A2(new_n458_), .A3(new_n342_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT20), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n481_), .B1(new_n472_), .B2(new_n460_), .ZN(new_n482_));
  AND2_X1   g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n475_), .B(new_n479_), .C1(new_n483_), .C2(new_n464_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n403_), .A2(new_n404_), .A3(new_n412_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n408_), .A2(new_n410_), .A3(new_n405_), .A4(new_n411_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(new_n418_), .A3(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n479_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n464_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n473_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n488_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n424_), .A2(new_n484_), .A3(new_n487_), .A4(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT94), .B1(new_n420_), .B2(new_n421_), .ZN(new_n493_));
  NOR3_X1   g292(.A1(new_n423_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n413_), .A2(new_n414_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(new_n418_), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n496_), .A2(new_n420_), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n342_), .A2(new_n466_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n481_), .B1(new_n498_), .B2(new_n470_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n464_), .B1(new_n461_), .B2(new_n499_), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n480_), .A2(new_n464_), .A3(new_n482_), .ZN(new_n501_));
  OAI211_X1 g300(.A(KEYINPUT32), .B(new_n479_), .C1(new_n500_), .C2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n479_), .A2(KEYINPUT32), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n475_), .B(new_n503_), .C1(new_n483_), .C2(new_n464_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n497_), .A2(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n390_), .B1(new_n494_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n484_), .A2(new_n491_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT27), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n488_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n511_), .A2(KEYINPUT27), .A3(new_n484_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(new_n497_), .A3(new_n389_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n507_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G227gat), .A2(G233gat), .ZN(new_n517_));
  INV_X1    g316(.A(G15gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT30), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n459_), .B(new_n521_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n522_), .A2(new_n398_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n522_), .A2(new_n398_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G71gat), .B(G99gat), .ZN(new_n525_));
  INV_X1    g324(.A(G43gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT31), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  OR3_X1    g328(.A1(new_n523_), .A2(new_n524_), .A3(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n529_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n513_), .A2(new_n389_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n530_), .A2(new_n531_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(new_n497_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  AOI22_X1  g335(.A1(new_n516_), .A2(new_n532_), .B1(new_n533_), .B2(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n328_), .B(new_n204_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G229gat), .A2(G233gat), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n328_), .A2(new_n205_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n539_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n328_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n542_), .B1(new_n543_), .B2(new_n204_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n540_), .B1(new_n541_), .B2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G113gat), .B(G141gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G169gat), .B(G197gat), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n546_), .B(new_n547_), .Z(new_n548_));
  XNOR2_X1  g347(.A(new_n545_), .B(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n537_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G230gat), .A2(G233gat), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n552_), .B1(new_n317_), .B2(new_n239_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT68), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n246_), .A2(new_n247_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n555_), .A2(new_n316_), .A3(new_n312_), .A4(new_n223_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT68), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n556_), .A2(new_n557_), .A3(new_n552_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n554_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT67), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(KEYINPUT12), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n313_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n315_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n561_), .B1(new_n564_), .B2(new_n248_), .ZN(new_n565_));
  XOR2_X1   g364(.A(KEYINPUT67), .B(KEYINPUT12), .Z(new_n566_));
  NAND3_X1  g365(.A1(new_n317_), .A2(new_n239_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT66), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n570_), .B1(new_n317_), .B2(new_n239_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n564_), .A2(KEYINPUT66), .A3(new_n248_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n571_), .B(new_n572_), .C1(new_n564_), .C2(new_n248_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n552_), .ZN(new_n574_));
  AOI22_X1  g373(.A1(new_n559_), .A2(new_n569_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G120gat), .B(G148gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT5), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G176gat), .B(G204gat), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n577_), .B(new_n578_), .Z(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n575_), .B(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  AND2_X1   g381(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n583_));
  NOR2_X1   g382(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n582_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n581_), .B1(KEYINPUT69), .B2(KEYINPUT13), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n334_), .A2(new_n551_), .A3(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n496_), .A2(new_n420_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(new_n589_), .A3(new_n323_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n591_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n278_), .A2(new_n270_), .A3(new_n281_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT96), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n537_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n587_), .A2(new_n549_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n598_), .A2(new_n330_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(G1gat), .B1(new_n600_), .B2(new_n497_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n592_), .A2(new_n593_), .A3(new_n601_), .ZN(G1324gat));
  NAND3_X1  g401(.A1(new_n588_), .A2(new_n324_), .A3(new_n513_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT97), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(G8gat), .B1(new_n600_), .B2(new_n514_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT39), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT40), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(G1325gat));
  OAI21_X1  g409(.A(G15gat), .B1(new_n600_), .B2(new_n532_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT98), .Z(new_n612_));
  OR2_X1    g411(.A1(new_n612_), .A2(KEYINPUT41), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(KEYINPUT41), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n588_), .A2(new_n518_), .A3(new_n534_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n613_), .A2(new_n614_), .A3(new_n615_), .ZN(G1326gat));
  XOR2_X1   g415(.A(new_n389_), .B(KEYINPUT99), .Z(new_n617_));
  NAND3_X1  g416(.A1(new_n597_), .A2(new_n599_), .A3(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(G22gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT42), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n588_), .A2(new_n321_), .A3(new_n617_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(G1327gat));
  NAND2_X1  g421(.A1(new_n596_), .A2(new_n331_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n587_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n625_), .A2(new_n551_), .ZN(new_n626_));
  INV_X1    g425(.A(G29gat), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n626_), .A2(new_n627_), .A3(new_n589_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT101), .ZN(new_n629_));
  INV_X1    g428(.A(new_n283_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT43), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n534_), .B1(new_n507_), .B2(new_n515_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n535_), .A2(new_n389_), .A3(new_n513_), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n630_), .B(new_n631_), .C1(new_n632_), .C2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT100), .ZN(new_n635_));
  OAI21_X1  g434(.A(KEYINPUT43), .B1(new_n537_), .B2(new_n283_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n493_), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n484_), .A2(new_n487_), .A3(new_n491_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n637_), .A2(new_n638_), .A3(new_n422_), .A4(new_n424_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n505_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(new_n589_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n389_), .B1(new_n639_), .B2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n389_), .A2(new_n497_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n643_), .A2(new_n513_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n532_), .B1(new_n642_), .B2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n536_), .A2(new_n533_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n647_), .A2(new_n648_), .A3(new_n631_), .A4(new_n630_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n635_), .A2(new_n636_), .A3(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n598_), .A2(new_n332_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT44), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n650_), .A2(KEYINPUT44), .A3(new_n651_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(new_n589_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n629_), .B1(new_n657_), .B2(G29gat), .ZN(new_n658_));
  AOI211_X1 g457(.A(KEYINPUT101), .B(new_n627_), .C1(new_n656_), .C2(new_n589_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n628_), .B1(new_n658_), .B2(new_n659_), .ZN(G1328gat));
  INV_X1    g459(.A(G36gat), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n513_), .A2(KEYINPUT103), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n513_), .A2(KEYINPUT103), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n626_), .A2(new_n661_), .A3(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT45), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n654_), .A2(new_n513_), .A3(new_n655_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT102), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n667_), .A2(new_n668_), .A3(G36gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n667_), .B2(G36gat), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n666_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT46), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  OAI211_X1 g472(.A(KEYINPUT46), .B(new_n666_), .C1(new_n669_), .C2(new_n670_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1329gat));
  NAND3_X1  g474(.A1(new_n656_), .A2(G43gat), .A3(new_n534_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n626_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n526_), .B1(new_n677_), .B2(new_n532_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n679_), .B(new_n680_), .ZN(G1330gat));
  AOI21_X1  g480(.A(G50gat), .B1(new_n626_), .B2(new_n617_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n389_), .A2(G50gat), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n682_), .B1(new_n656_), .B2(new_n683_), .ZN(G1331gat));
  NOR2_X1   g483(.A1(new_n331_), .A2(new_n549_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n597_), .A2(new_n624_), .A3(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(G57gat), .B1(new_n686_), .B2(new_n497_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n647_), .A2(new_n550_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT105), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(new_n624_), .A3(new_n334_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT106), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n690_), .B(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n589_), .A2(new_n296_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n687_), .B1(new_n692_), .B2(new_n693_), .ZN(G1332gat));
  INV_X1    g493(.A(new_n664_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G64gat), .B1(new_n686_), .B2(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT48), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n664_), .A2(new_n298_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n697_), .B1(new_n692_), .B2(new_n698_), .ZN(G1333gat));
  OAI21_X1  g498(.A(G71gat), .B1(new_n686_), .B2(new_n532_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT49), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n534_), .A2(new_n301_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(new_n692_), .B2(new_n702_), .ZN(G1334gat));
  NAND4_X1  g502(.A1(new_n597_), .A2(new_n624_), .A3(new_n617_), .A4(new_n685_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(G78gat), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT50), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n617_), .A2(new_n303_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n706_), .B1(new_n692_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n708_), .B(new_n709_), .ZN(G1335gat));
  AND4_X1   g509(.A1(new_n624_), .A2(new_n689_), .A3(new_n331_), .A4(new_n596_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n711_), .A2(new_n209_), .A3(new_n589_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n650_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n332_), .A2(new_n549_), .A3(new_n587_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n713_), .A2(new_n497_), .A3(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n712_), .B1(new_n209_), .B2(new_n716_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT108), .Z(G1336gat));
  NAND3_X1  g517(.A1(new_n711_), .A2(new_n210_), .A3(new_n513_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n713_), .A2(new_n695_), .A3(new_n715_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n210_), .B2(new_n720_), .ZN(G1337gat));
  NAND4_X1  g520(.A1(new_n711_), .A2(new_n534_), .A3(new_n219_), .A4(new_n221_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n650_), .A2(new_n534_), .A3(new_n714_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n723_), .A2(new_n724_), .A3(G99gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n723_), .B2(G99gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n722_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g527(.A1(new_n711_), .A2(new_n220_), .A3(new_n389_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n650_), .A2(new_n389_), .A3(new_n714_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT52), .ZN(new_n731_));
  AND4_X1   g530(.A1(KEYINPUT110), .A2(new_n730_), .A3(new_n731_), .A4(G106gat), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n220_), .B1(new_n733_), .B2(KEYINPUT52), .ZN(new_n734_));
  AOI22_X1  g533(.A1(new_n730_), .A2(new_n734_), .B1(KEYINPUT110), .B2(new_n731_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n729_), .B1(new_n732_), .B2(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g536(.A1(new_n685_), .A2(new_n283_), .A3(new_n587_), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT54), .Z(new_n739_));
  NAND2_X1  g538(.A1(new_n575_), .A2(new_n580_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n550_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT55), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n559_), .A2(new_n569_), .A3(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n559_), .B2(new_n569_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n565_), .A2(new_n571_), .A3(new_n572_), .A4(new_n567_), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n746_), .A2(KEYINPUT111), .A3(new_n574_), .ZN(new_n747_));
  AOI21_X1  g546(.A(KEYINPUT111), .B1(new_n746_), .B2(new_n574_), .ZN(new_n748_));
  OAI22_X1  g547(.A1(new_n744_), .A2(new_n745_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT112), .ZN(new_n750_));
  AOI211_X1 g549(.A(KEYINPUT68), .B(new_n574_), .C1(new_n564_), .C2(new_n248_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n557_), .B1(new_n556_), .B2(new_n552_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT55), .B1(new_n753_), .B2(new_n568_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n559_), .A2(new_n569_), .A3(new_n743_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n746_), .A2(new_n574_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT111), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n746_), .A2(KEYINPUT111), .A3(new_n574_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT112), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n756_), .A2(new_n761_), .A3(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n580_), .B1(new_n750_), .B2(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(KEYINPUT113), .B1(new_n764_), .B2(KEYINPUT56), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n756_), .A2(new_n761_), .A3(new_n762_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n762_), .B1(new_n756_), .B2(new_n761_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n579_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT56), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n768_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n765_), .A2(new_n771_), .ZN(new_n772_));
  OAI211_X1 g571(.A(KEYINPUT56), .B(new_n579_), .C1(new_n766_), .C2(new_n767_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n764_), .A2(KEYINPUT114), .A3(KEYINPUT56), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n742_), .B1(new_n772_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n543_), .A2(new_n204_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(new_n542_), .A3(new_n541_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n548_), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n780_), .B(new_n781_), .C1(new_n538_), .C2(new_n542_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n545_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n782_), .B1(new_n783_), .B2(new_n781_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n784_), .A2(new_n582_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n596_), .B1(new_n778_), .B2(new_n786_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n784_), .A2(new_n741_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n764_), .A2(KEYINPUT56), .ZN(new_n789_));
  INV_X1    g588(.A(new_n773_), .ZN(new_n790_));
  OAI211_X1 g589(.A(KEYINPUT58), .B(new_n788_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT117), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n768_), .A2(new_n770_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n773_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT117), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n794_), .A2(new_n795_), .A3(KEYINPUT58), .A4(new_n788_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n792_), .A2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT58), .B1(new_n794_), .B2(new_n788_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n798_), .A2(new_n283_), .ZN(new_n799_));
  AOI22_X1  g598(.A1(new_n787_), .A2(KEYINPUT57), .B1(new_n797_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n801_));
  XNOR2_X1  g600(.A(KEYINPUT115), .B(KEYINPUT57), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n787_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n802_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n765_), .A2(new_n771_), .A3(new_n775_), .A4(new_n776_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n785_), .B1(new_n805_), .B2(new_n742_), .ZN(new_n806_));
  OAI211_X1 g605(.A(KEYINPUT116), .B(new_n804_), .C1(new_n806_), .C2(new_n596_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n800_), .A2(new_n803_), .A3(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n739_), .B1(new_n808_), .B2(new_n330_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n532_), .A2(new_n497_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n533_), .ZN(new_n811_));
  OAI21_X1  g610(.A(KEYINPUT59), .B1(new_n809_), .B2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n804_), .B1(new_n806_), .B2(new_n596_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n800_), .A2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n739_), .B1(new_n814_), .B2(new_n331_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT59), .ZN(new_n817_));
  INV_X1    g616(.A(new_n811_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n817_), .B1(new_n818_), .B2(KEYINPUT118), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n819_), .B1(KEYINPUT118), .B2(new_n818_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n816_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(G113gat), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n550_), .A2(new_n822_), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n812_), .A2(new_n821_), .A3(new_n823_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n809_), .A2(new_n811_), .ZN(new_n825_));
  AOI21_X1  g624(.A(G113gat), .B1(new_n825_), .B2(new_n549_), .ZN(new_n826_));
  OAI21_X1  g625(.A(KEYINPUT119), .B1(new_n824_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n808_), .A2(new_n330_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n739_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n818_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n822_), .B1(new_n831_), .B2(new_n550_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n812_), .A2(new_n821_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n823_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n832_), .B(new_n833_), .C1(new_n834_), .C2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n827_), .A2(new_n836_), .ZN(G1340gat));
  OAI21_X1  g636(.A(G120gat), .B1(new_n834_), .B2(new_n587_), .ZN(new_n838_));
  INV_X1    g637(.A(G120gat), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n839_), .B1(new_n587_), .B2(KEYINPUT60), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(KEYINPUT60), .B2(new_n839_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n838_), .B1(new_n831_), .B2(new_n841_), .ZN(G1341gat));
  AOI21_X1  g641(.A(G127gat), .B1(new_n825_), .B2(new_n332_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n834_), .ZN(new_n844_));
  INV_X1    g643(.A(G127gat), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT120), .ZN(new_n846_));
  OR2_X1    g645(.A1(new_n845_), .A2(KEYINPUT120), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n330_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n843_), .B1(new_n844_), .B2(new_n848_), .ZN(G1342gat));
  OAI21_X1  g648(.A(G134gat), .B1(new_n834_), .B2(new_n283_), .ZN(new_n850_));
  INV_X1    g649(.A(G134gat), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n825_), .A2(new_n851_), .A3(new_n596_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(G1343gat));
  NOR3_X1   g652(.A1(new_n664_), .A2(new_n497_), .A3(new_n390_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n809_), .A2(new_n534_), .A3(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n549_), .ZN(new_n857_));
  XOR2_X1   g656(.A(KEYINPUT121), .B(G141gat), .Z(new_n858_));
  XNOR2_X1  g657(.A(new_n857_), .B(new_n858_), .ZN(G1344gat));
  NAND2_X1  g658(.A1(new_n856_), .A2(new_n624_), .ZN(new_n860_));
  XOR2_X1   g659(.A(KEYINPUT122), .B(G148gat), .Z(new_n861_));
  XNOR2_X1  g660(.A(new_n860_), .B(new_n861_), .ZN(G1345gat));
  XNOR2_X1  g661(.A(KEYINPUT61), .B(G155gat), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n830_), .A2(new_n532_), .A3(new_n332_), .A4(new_n854_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n865_), .A2(KEYINPUT123), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT123), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n867_), .B1(new_n856_), .B2(new_n332_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n864_), .B1(new_n866_), .B2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n865_), .A2(KEYINPUT123), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n856_), .A2(new_n867_), .A3(new_n332_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n870_), .A2(new_n871_), .A3(new_n863_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n869_), .A2(new_n872_), .ZN(G1346gat));
  INV_X1    g672(.A(new_n856_), .ZN(new_n874_));
  OAI21_X1  g673(.A(G162gat), .B1(new_n874_), .B2(new_n283_), .ZN(new_n875_));
  INV_X1    g674(.A(G162gat), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n856_), .A2(new_n876_), .A3(new_n596_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(G1347gat));
  INV_X1    g677(.A(KEYINPUT62), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n695_), .A2(new_n535_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  NOR4_X1   g680(.A1(new_n815_), .A2(new_n550_), .A3(new_n617_), .A4(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT22), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n879_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(G169gat), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n425_), .B1(new_n882_), .B2(new_n879_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n884_), .B2(new_n886_), .ZN(G1348gat));
  NOR3_X1   g686(.A1(new_n815_), .A2(new_n617_), .A3(new_n881_), .ZN(new_n888_));
  AOI21_X1  g687(.A(G176gat), .B1(new_n888_), .B2(new_n624_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n809_), .A2(new_n389_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n881_), .A2(new_n587_), .A3(new_n426_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n889_), .B1(new_n890_), .B2(new_n891_), .ZN(G1349gat));
  NOR2_X1   g691(.A1(new_n881_), .A2(new_n617_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n330_), .A2(new_n445_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n816_), .A2(new_n893_), .A3(new_n894_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(KEYINPUT124), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n881_), .A2(new_n331_), .ZN(new_n897_));
  AOI21_X1  g696(.A(G183gat), .B1(new_n890_), .B2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n896_), .A2(new_n898_), .ZN(G1350gat));
  NAND3_X1  g698(.A1(new_n888_), .A2(new_n446_), .A3(new_n596_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n888_), .A2(new_n630_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n432_), .ZN(G1351gat));
  NOR2_X1   g701(.A1(new_n695_), .A2(new_n643_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n830_), .A2(new_n532_), .A3(new_n549_), .A4(new_n903_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(KEYINPUT125), .A2(G197gat), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT125), .B(G197gat), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n904_), .B2(new_n907_), .ZN(G1352gat));
  NAND2_X1  g707(.A1(new_n830_), .A2(new_n532_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n903_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n909_), .A2(new_n587_), .A3(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(G204gat), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n911_), .B(new_n912_), .ZN(G1353gat));
  NOR2_X1   g712(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(KEYINPUT126), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n909_), .A2(new_n910_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n330_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n915_), .B1(new_n916_), .B2(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n915_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n917_), .ZN(new_n920_));
  NOR4_X1   g719(.A1(new_n909_), .A2(new_n910_), .A3(new_n919_), .A4(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n918_), .A2(new_n921_), .ZN(G1354gat));
  NAND2_X1  g721(.A1(new_n916_), .A2(new_n596_), .ZN(new_n923_));
  INV_X1    g722(.A(G218gat), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n283_), .A2(new_n924_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(KEYINPUT127), .ZN(new_n926_));
  AOI22_X1  g725(.A1(new_n923_), .A2(new_n924_), .B1(new_n916_), .B2(new_n926_), .ZN(G1355gat));
endmodule


