//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 0 1 1 0 1 0 0 0 1 1 0 0 0 1 1 0 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 1 0 1 1 0 1 0 0 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n841_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n877_, new_n878_, new_n879_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G71gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G78gat), .ZN(new_n211_));
  INV_X1    g010(.A(G78gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(G71gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G57gat), .B(G64gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n214_), .B1(new_n215_), .B2(KEYINPUT11), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT68), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n217_), .B1(new_n215_), .B2(KEYINPUT11), .ZN(new_n218_));
  INV_X1    g017(.A(G64gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(G57gat), .ZN(new_n220_));
  INV_X1    g019(.A(G57gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(G64gat), .ZN(new_n222_));
  AND4_X1   g021(.A1(new_n217_), .A2(new_n220_), .A3(new_n222_), .A4(KEYINPUT11), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n216_), .B1(new_n218_), .B2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n220_), .A2(new_n222_), .A3(KEYINPUT11), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT68), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n220_), .A2(new_n222_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT11), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n220_), .A2(new_n222_), .A3(new_n217_), .A4(KEYINPUT11), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n226_), .A2(new_n229_), .A3(new_n214_), .A4(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n224_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n209_), .B(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G231gat), .A2(G233gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT77), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(G183gat), .B(G211gat), .Z(new_n238_));
  XNOR2_X1  g037(.A(G127gat), .B(G155gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n237_), .B(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n242_));
  OR2_X1    g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n242_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT17), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n235_), .A2(new_n246_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n243_), .A2(new_n244_), .A3(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT37), .ZN(new_n251_));
  XOR2_X1   g050(.A(KEYINPUT71), .B(KEYINPUT35), .Z(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G232gat), .A2(G233gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT34), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n253_), .A2(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n253_), .A2(new_n255_), .ZN(new_n257_));
  INV_X1    g056(.A(G85gat), .ZN(new_n258_));
  INV_X1    g057(.A(G92gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G85gat), .A2(G92gat), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G99gat), .A2(G106gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT6), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT6), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(G99gat), .A3(G106gat), .ZN(new_n266_));
  AND2_X1   g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT7), .ZN(new_n268_));
  INV_X1    g067(.A(G99gat), .ZN(new_n269_));
  INV_X1    g068(.A(G106gat), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n268_), .A2(new_n269_), .A3(new_n270_), .A4(KEYINPUT67), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT67), .ZN(new_n272_));
  OAI22_X1  g071(.A1(new_n272_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n262_), .B1(new_n267_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT8), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  OAI211_X1 g076(.A(KEYINPUT8), .B(new_n262_), .C1(new_n267_), .C2(new_n274_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT10), .B(G99gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT65), .B1(new_n279_), .B2(G106gat), .ZN(new_n280_));
  AND2_X1   g079(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n281_));
  NOR2_X1   g080(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT65), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n283_), .A2(new_n284_), .A3(new_n270_), .ZN(new_n285_));
  OR2_X1    g084(.A1(KEYINPUT66), .A2(KEYINPUT9), .ZN(new_n286_));
  NAND2_X1  g085(.A1(KEYINPUT66), .A2(KEYINPUT9), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n286_), .A2(new_n260_), .A3(new_n261_), .A4(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n261_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT9), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n264_), .A2(new_n266_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n280_), .A2(new_n285_), .A3(new_n288_), .A4(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n277_), .A2(new_n278_), .A3(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G43gat), .B(G50gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(G36gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(G29gat), .ZN(new_n298_));
  INV_X1    g097(.A(G29gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(G36gat), .ZN(new_n300_));
  AND3_X1   g099(.A1(new_n298_), .A2(new_n300_), .A3(KEYINPUT72), .ZN(new_n301_));
  AOI21_X1  g100(.A(KEYINPUT72), .B1(new_n298_), .B2(new_n300_), .ZN(new_n302_));
  NOR3_X1   g101(.A1(new_n301_), .A2(new_n302_), .A3(KEYINPUT73), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT73), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT72), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n299_), .A2(G36gat), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n297_), .A2(G29gat), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n305_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n298_), .A2(new_n300_), .A3(KEYINPUT72), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n304_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n296_), .B1(new_n303_), .B2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT73), .B1(new_n301_), .B2(new_n302_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n308_), .A2(new_n304_), .A3(new_n309_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n312_), .A2(new_n313_), .A3(new_n295_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n311_), .A2(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n257_), .B1(new_n294_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT74), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n256_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT15), .ZN(new_n319_));
  AND3_X1   g118(.A1(new_n312_), .A2(new_n295_), .A3(new_n313_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n295_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n319_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n311_), .A2(KEYINPUT15), .A3(new_n314_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n322_), .A2(new_n323_), .A3(new_n293_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n316_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n318_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT75), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n316_), .B(new_n324_), .C1(new_n317_), .C2(new_n256_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT36), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G190gat), .B(G218gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G134gat), .B(G162gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n329_), .A2(new_n330_), .A3(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n326_), .A2(new_n333_), .A3(new_n328_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n330_), .B1(new_n329_), .B2(new_n334_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n251_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n338_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n340_), .A2(KEYINPUT37), .A3(new_n336_), .A4(new_n335_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n250_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT78), .ZN(new_n344_));
  NOR3_X1   g143(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(KEYINPUT25), .B(G183gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT26), .B(G190gat), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n345_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G183gat), .A2(G190gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT23), .ZN(new_n350_));
  INV_X1    g149(.A(G169gat), .ZN(new_n351_));
  INV_X1    g150(.A(G176gat), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n348_), .B(new_n350_), .C1(new_n353_), .C2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n350_), .B1(G183gat), .B2(G190gat), .ZN(new_n356_));
  NOR2_X1   g155(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(G169gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n355_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G71gat), .B(G99gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(G43gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n360_), .B(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G127gat), .B(G134gat), .Z(new_n364_));
  XOR2_X1   g163(.A(G113gat), .B(G120gat), .Z(new_n365_));
  XOR2_X1   g164(.A(new_n364_), .B(new_n365_), .Z(new_n366_));
  XNOR2_X1  g165(.A(new_n363_), .B(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G227gat), .A2(G233gat), .ZN(new_n368_));
  INV_X1    g167(.A(G15gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT30), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT31), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n367_), .B(new_n372_), .Z(new_n373_));
  XOR2_X1   g172(.A(G1gat), .B(G29gat), .Z(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G57gat), .B(G85gat), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n376_), .B(new_n377_), .Z(new_n378_));
  NAND2_X1  g177(.A1(G225gat), .A2(G233gat), .ZN(new_n379_));
  NOR2_X1   g178(.A1(G155gat), .A2(G162gat), .ZN(new_n380_));
  XOR2_X1   g179(.A(new_n380_), .B(KEYINPUT83), .Z(new_n381_));
  NAND2_X1  g180(.A1(G155gat), .A2(G162gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT84), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(G141gat), .A2(G148gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT3), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G141gat), .A2(G148gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT2), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT85), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n386_), .A2(KEYINPUT85), .A3(new_n388_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n384_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n383_), .A2(KEYINPUT1), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT84), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n382_), .B(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT1), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n395_), .A2(new_n399_), .A3(new_n381_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n385_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n400_), .A2(new_n401_), .A3(new_n387_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n366_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n394_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n400_), .A2(new_n401_), .A3(new_n387_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n366_), .B1(new_n405_), .B2(new_n393_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n404_), .A2(new_n406_), .A3(KEYINPUT4), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n394_), .A2(new_n402_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT4), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(new_n409_), .A3(new_n366_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n379_), .B1(new_n407_), .B2(new_n410_), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n404_), .A2(new_n406_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n379_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n378_), .B1(new_n411_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT95), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT33), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT33), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n415_), .A2(new_n416_), .A3(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G8gat), .B(G36gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G64gat), .B(G92gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT20), .ZN(new_n427_));
  XOR2_X1   g226(.A(G211gat), .B(G218gat), .Z(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT88), .B(G197gat), .ZN(new_n429_));
  INV_X1    g228(.A(G204gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT21), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n432_), .B1(G197gat), .B2(G204gat), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n428_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(G197gat), .A2(G204gat), .ZN(new_n435_));
  XOR2_X1   g234(.A(KEYINPUT88), .B(G197gat), .Z(new_n436_));
  AOI21_X1  g235(.A(new_n435_), .B1(new_n436_), .B2(G204gat), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n434_), .B1(KEYINPUT21), .B2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(KEYINPUT21), .A3(new_n428_), .ZN(new_n439_));
  AND2_X1   g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n360_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n427_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n438_), .A2(new_n439_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n360_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G226gat), .A2(G233gat), .ZN(new_n445_));
  XOR2_X1   g244(.A(new_n445_), .B(KEYINPUT19), .Z(new_n446_));
  AND3_X1   g245(.A1(new_n442_), .A2(new_n444_), .A3(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n446_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n426_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n442_), .A2(new_n444_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n446_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n442_), .A2(new_n444_), .A3(new_n446_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n452_), .A2(new_n425_), .A3(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n449_), .A2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n378_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n407_), .A2(new_n410_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n456_), .B1(new_n413_), .B2(new_n457_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n418_), .A2(new_n420_), .A3(new_n455_), .A4(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n413_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n378_), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n460_), .B(new_n461_), .C1(new_n413_), .C2(new_n412_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT96), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(new_n463_), .A3(new_n415_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n452_), .A2(new_n453_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n426_), .A2(KEYINPUT32), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  OAI211_X1 g266(.A(KEYINPUT96), .B(new_n378_), .C1(new_n411_), .C2(new_n414_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n464_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n459_), .A2(new_n469_), .ZN(new_n470_));
  AND2_X1   g269(.A1(KEYINPUT86), .A2(G233gat), .ZN(new_n471_));
  NOR2_X1   g270(.A1(KEYINPUT86), .A2(G233gat), .ZN(new_n472_));
  OAI21_X1  g271(.A(G228gat), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT87), .ZN(new_n474_));
  XOR2_X1   g273(.A(new_n474_), .B(KEYINPUT89), .Z(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT29), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n477_), .B1(new_n394_), .B2(new_n402_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n476_), .B1(new_n478_), .B2(new_n440_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G78gat), .B(G106gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT90), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n474_), .A2(KEYINPUT89), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n405_), .A2(new_n393_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n443_), .B(new_n483_), .C1(new_n484_), .C2(new_n477_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n479_), .A2(new_n481_), .A3(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT91), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G22gat), .B(G50gat), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NOR3_X1   g289(.A1(new_n408_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT28), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n492_), .B1(new_n484_), .B2(new_n477_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n490_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT28), .B1(new_n408_), .B2(KEYINPUT29), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n484_), .A2(new_n492_), .A3(new_n477_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(new_n496_), .A3(new_n489_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n494_), .A2(new_n497_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n479_), .A2(KEYINPUT91), .A3(new_n485_), .A4(new_n481_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n479_), .A2(new_n485_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n481_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n488_), .A2(new_n498_), .A3(new_n499_), .A4(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n486_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n480_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n505_), .B1(new_n479_), .B2(new_n485_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n497_), .B(new_n494_), .C1(new_n504_), .C2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT92), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n503_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n508_), .B1(new_n503_), .B2(new_n507_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n470_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n503_), .A2(new_n507_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT92), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(new_n509_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n464_), .A2(new_n468_), .ZN(new_n517_));
  XOR2_X1   g316(.A(KEYINPUT98), .B(KEYINPUT27), .Z(new_n518_));
  NOR2_X1   g317(.A1(new_n455_), .A2(new_n518_), .ZN(new_n519_));
  NOR3_X1   g318(.A1(new_n447_), .A2(new_n448_), .A3(new_n426_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n425_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n521_));
  OAI21_X1  g320(.A(KEYINPUT27), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT97), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT97), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n455_), .A2(new_n524_), .A3(KEYINPUT27), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n519_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n516_), .A2(new_n517_), .A3(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n373_), .B1(new_n513_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n464_), .A2(new_n468_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n373_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT99), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n523_), .A2(new_n525_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n519_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n533_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  AOI211_X1 g335(.A(KEYINPUT99), .B(new_n519_), .C1(new_n523_), .C2(new_n525_), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n532_), .B(new_n512_), .C1(new_n536_), .C2(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n538_), .A2(KEYINPUT100), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT100), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n524_), .B1(new_n455_), .B2(KEYINPUT27), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT27), .ZN(new_n542_));
  AOI211_X1 g341(.A(KEYINPUT97), .B(new_n542_), .C1(new_n449_), .C2(new_n454_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n535_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT99), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n534_), .A2(new_n533_), .A3(new_n535_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n516_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n540_), .B1(new_n547_), .B2(new_n532_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n529_), .B1(new_n539_), .B2(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n209_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n311_), .A2(new_n208_), .A3(new_n314_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(KEYINPUT79), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G229gat), .A2(G233gat), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT79), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n311_), .A2(new_n555_), .A3(new_n208_), .A4(new_n314_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n552_), .A2(new_n554_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT80), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n552_), .A2(new_n556_), .A3(KEYINPUT80), .A4(new_n554_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n322_), .A2(new_n208_), .A3(new_n323_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n562_), .A2(new_n553_), .A3(new_n550_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT81), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n562_), .A2(KEYINPUT81), .A3(new_n553_), .A4(new_n550_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n561_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G113gat), .B(G141gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT82), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G169gat), .B(G197gat), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n570_), .B(new_n571_), .Z(new_n572_));
  NAND2_X1  g371(.A1(new_n568_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n572_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n561_), .A2(new_n567_), .A3(new_n574_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n549_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT13), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G120gat), .B(G148gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT5), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G176gat), .B(G204gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n224_), .A2(new_n231_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n284_), .B1(new_n283_), .B2(new_n270_), .ZN(new_n586_));
  NOR4_X1   g385(.A1(new_n281_), .A2(new_n282_), .A3(KEYINPUT65), .A4(G106gat), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n291_), .A2(new_n288_), .ZN(new_n589_));
  AOI22_X1  g388(.A1(new_n588_), .A2(new_n589_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n585_), .A2(new_n590_), .A3(new_n278_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n293_), .A2(new_n232_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G230gat), .A2(G233gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT64), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT69), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n593_), .A2(KEYINPUT69), .A3(new_n595_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n591_), .A2(new_n592_), .A3(KEYINPUT12), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT12), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n293_), .A2(new_n602_), .A3(new_n232_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n595_), .B1(new_n601_), .B2(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n584_), .B1(new_n600_), .B2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n601_), .A2(new_n603_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n595_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n608_), .A2(new_n598_), .A3(new_n599_), .A4(new_n583_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n605_), .A2(new_n609_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n610_), .A2(KEYINPUT70), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(KEYINPUT70), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n579_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n611_), .A2(new_n612_), .A3(new_n579_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NOR3_X1   g416(.A1(new_n344_), .A2(new_n578_), .A3(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n618_), .A2(new_n203_), .A3(new_n530_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n620_), .A2(KEYINPUT38), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT102), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n538_), .A2(KEYINPUT100), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n547_), .A2(new_n540_), .A3(new_n532_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n528_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n337_), .A2(new_n338_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n615_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n629_), .A2(new_n577_), .A3(new_n613_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT101), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n628_), .A2(new_n250_), .A3(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n203_), .B1(new_n632_), .B2(new_n530_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n633_), .B1(new_n620_), .B2(KEYINPUT38), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n622_), .A2(new_n634_), .ZN(G1324gat));
  NAND2_X1  g434(.A1(new_n545_), .A2(new_n546_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n618_), .A2(new_n204_), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n632_), .A2(new_n637_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(KEYINPUT103), .B(KEYINPUT39), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n639_), .A2(G8gat), .A3(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n640_), .B1(new_n639_), .B2(G8gat), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n638_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT40), .Z(G1325gat));
  AOI21_X1  g443(.A(new_n369_), .B1(new_n632_), .B2(new_n373_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT41), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n618_), .A2(new_n369_), .A3(new_n373_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(G1326gat));
  INV_X1    g447(.A(G22gat), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n618_), .A2(new_n649_), .A3(new_n516_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n632_), .B2(new_n516_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n651_), .A2(new_n652_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n650_), .B1(new_n653_), .B2(new_n654_), .ZN(G1327gat));
  NAND3_X1  g454(.A1(new_n247_), .A2(new_n627_), .A3(new_n249_), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n578_), .A2(new_n617_), .A3(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(new_n299_), .A3(new_n530_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n342_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n549_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT43), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n250_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n549_), .A2(KEYINPUT43), .A3(new_n659_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n662_), .A2(KEYINPUT44), .A3(new_n631_), .A4(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n661_), .B1(new_n625_), .B2(new_n342_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n247_), .A2(new_n249_), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n663_), .A2(new_n665_), .A3(new_n666_), .A4(new_n631_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n664_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(new_n530_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n671_), .A2(KEYINPUT105), .ZN(new_n672_));
  OAI21_X1  g471(.A(G29gat), .B1(new_n671_), .B2(KEYINPUT105), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n658_), .B1(new_n672_), .B2(new_n673_), .ZN(G1328gat));
  INV_X1    g473(.A(KEYINPUT106), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n675_), .A2(KEYINPUT46), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n664_), .A2(new_n669_), .A3(new_n637_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G36gat), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n617_), .A2(new_n656_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n636_), .A2(G36gat), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n549_), .A2(new_n679_), .A3(new_n577_), .A4(new_n680_), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT45), .Z(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n678_), .A2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT107), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT107), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n678_), .A2(new_n686_), .A3(new_n683_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n676_), .B1(new_n685_), .B2(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n686_), .B1(new_n678_), .B2(new_n683_), .ZN(new_n689_));
  AOI211_X1 g488(.A(KEYINPUT107), .B(new_n682_), .C1(new_n677_), .C2(G36gat), .ZN(new_n690_));
  INV_X1    g489(.A(new_n676_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n689_), .A2(new_n690_), .A3(new_n691_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n688_), .A2(new_n692_), .ZN(G1329gat));
  NAND3_X1  g492(.A1(new_n664_), .A2(new_n669_), .A3(new_n373_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(G43gat), .ZN(new_n695_));
  INV_X1    g494(.A(G43gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n657_), .A2(new_n696_), .A3(new_n373_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g498(.A(G50gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n657_), .A2(new_n700_), .A3(new_n516_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n670_), .A2(KEYINPUT108), .A3(new_n516_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(G50gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT108), .B1(new_n670_), .B2(new_n516_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n701_), .B1(new_n703_), .B2(new_n704_), .ZN(G1331gat));
  NOR2_X1   g504(.A1(new_n344_), .A2(new_n616_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT109), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n625_), .A2(new_n577_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT110), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n710_), .A2(new_n221_), .A3(new_n530_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n666_), .A2(new_n577_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n628_), .A2(new_n617_), .A3(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(G57gat), .B1(new_n713_), .B2(new_n517_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n711_), .A2(new_n714_), .ZN(G1332gat));
  NOR2_X1   g514(.A1(new_n636_), .A2(G64gat), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT111), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n710_), .A2(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(G64gat), .B1(new_n713_), .B2(new_n636_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT48), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1333gat));
  NAND3_X1  g520(.A1(new_n710_), .A2(new_n210_), .A3(new_n373_), .ZN(new_n722_));
  OAI21_X1  g521(.A(G71gat), .B1(new_n713_), .B2(new_n531_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT49), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(G1334gat));
  NAND3_X1  g524(.A1(new_n710_), .A2(new_n212_), .A3(new_n516_), .ZN(new_n726_));
  OAI21_X1  g525(.A(G78gat), .B1(new_n713_), .B2(new_n512_), .ZN(new_n727_));
  XOR2_X1   g526(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n728_));
  XNOR2_X1  g527(.A(new_n727_), .B(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n726_), .A2(new_n729_), .ZN(G1335gat));
  NOR2_X1   g529(.A1(new_n616_), .A2(new_n577_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n662_), .A2(new_n663_), .A3(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(G85gat), .B1(new_n732_), .B2(new_n517_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n709_), .A2(new_n617_), .A3(new_n627_), .A4(new_n666_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n530_), .A2(new_n258_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n733_), .B1(new_n734_), .B2(new_n735_), .ZN(G1336gat));
  OAI21_X1  g535(.A(G92gat), .B1(new_n732_), .B2(new_n636_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n637_), .A2(new_n259_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n737_), .B1(new_n734_), .B2(new_n738_), .ZN(G1337gat));
  INV_X1    g538(.A(KEYINPUT113), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT51), .ZN(new_n741_));
  OAI21_X1  g540(.A(KEYINPUT114), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(G99gat), .B1(new_n732_), .B2(new_n531_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n373_), .A2(new_n283_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(new_n734_), .B2(new_n744_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n741_), .A2(KEYINPUT114), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n742_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n747_), .B1(new_n742_), .B2(new_n745_), .ZN(G1338gat));
  OAI21_X1  g547(.A(G106gat), .B1(new_n732_), .B2(new_n512_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n749_), .A2(KEYINPUT52), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n751_), .B(G106gat), .C1(new_n732_), .C2(new_n512_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n516_), .A2(new_n270_), .ZN(new_n754_));
  OAI22_X1  g553(.A1(new_n750_), .A2(new_n753_), .B1(new_n734_), .B2(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g555(.A(KEYINPUT54), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n712_), .A2(new_n757_), .A3(new_n616_), .A4(new_n342_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n616_), .A2(new_n576_), .A3(new_n250_), .ZN(new_n759_));
  OAI21_X1  g558(.A(KEYINPUT54), .B1(new_n759_), .B2(new_n659_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n758_), .A2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n552_), .A2(new_n553_), .A3(new_n556_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n562_), .A2(new_n554_), .A3(new_n550_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n762_), .A2(new_n763_), .A3(new_n572_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n575_), .A2(KEYINPUT116), .A3(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(KEYINPUT116), .B1(new_n575_), .B2(new_n764_), .ZN(new_n767_));
  OAI22_X1  g566(.A1(new_n611_), .A2(new_n612_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n601_), .A2(new_n595_), .A3(new_n603_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n769_), .A2(new_n604_), .A3(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n606_), .A2(new_n770_), .A3(new_n607_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(new_n584_), .ZN(new_n773_));
  OAI21_X1  g572(.A(KEYINPUT56), .B1(new_n771_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT56), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n583_), .B1(new_n604_), .B2(new_n770_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n608_), .A2(KEYINPUT55), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n775_), .B(new_n776_), .C1(new_n777_), .C2(new_n769_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n774_), .A2(new_n609_), .A3(new_n778_), .ZN(new_n779_));
  OR3_X1    g578(.A1(new_n576_), .A2(new_n779_), .A3(KEYINPUT115), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT115), .B1(new_n576_), .B2(new_n779_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n768_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n626_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT57), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT58), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n575_), .A2(new_n764_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT116), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n779_), .B1(new_n789_), .B2(new_n765_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n786_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n774_), .A2(new_n609_), .A3(new_n778_), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n793_), .B(new_n791_), .C1(new_n766_), .C2(new_n767_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  OAI211_X1 g594(.A(KEYINPUT118), .B(new_n659_), .C1(new_n792_), .C2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n790_), .A2(KEYINPUT58), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n793_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT117), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n800_), .A2(new_n786_), .A3(new_n794_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT118), .B1(new_n801_), .B2(new_n659_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n785_), .B1(new_n798_), .B2(new_n802_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n783_), .A2(new_n784_), .ZN(new_n804_));
  OR2_X1    g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n761_), .B1(new_n805_), .B2(new_n666_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n547_), .A2(new_n530_), .A3(new_n373_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(G113gat), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(new_n809_), .A3(new_n577_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT59), .B1(new_n806_), .B2(new_n807_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n804_), .B1(new_n803_), .B2(KEYINPUT120), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT120), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n785_), .B(new_n813_), .C1(new_n798_), .C2(new_n802_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n666_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n761_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT59), .B1(new_n807_), .B2(KEYINPUT119), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n820_), .B1(KEYINPUT119), .B2(new_n807_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n811_), .B(new_n577_), .C1(new_n819_), .C2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n810_), .B1(new_n823_), .B2(new_n809_), .ZN(G1340gat));
  INV_X1    g623(.A(G120gat), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n825_), .B1(new_n616_), .B2(KEYINPUT60), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n808_), .B(new_n826_), .C1(KEYINPUT60), .C2(new_n825_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n811_), .B(new_n617_), .C1(new_n819_), .C2(new_n821_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n827_), .B1(new_n829_), .B2(new_n825_), .ZN(G1341gat));
  INV_X1    g629(.A(G127gat), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n808_), .A2(new_n831_), .A3(new_n250_), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n811_), .B(new_n250_), .C1(new_n819_), .C2(new_n821_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n832_), .B1(new_n834_), .B2(new_n831_), .ZN(G1342gat));
  INV_X1    g634(.A(G134gat), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n808_), .A2(new_n836_), .A3(new_n627_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n811_), .B(new_n659_), .C1(new_n819_), .C2(new_n821_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n837_), .B1(new_n839_), .B2(new_n836_), .ZN(G1343gat));
  NAND2_X1  g639(.A1(new_n805_), .A2(new_n666_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n373_), .B1(new_n841_), .B2(new_n817_), .ZN(new_n842_));
  AND4_X1   g641(.A1(new_n516_), .A2(new_n842_), .A3(new_n530_), .A4(new_n636_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n577_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n617_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g646(.A1(new_n843_), .A2(new_n250_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT61), .B(G155gat), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n848_), .B(new_n849_), .ZN(G1346gat));
  AOI21_X1  g649(.A(G162gat), .B1(new_n843_), .B2(new_n627_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n659_), .A2(G162gat), .ZN(new_n852_));
  XOR2_X1   g651(.A(new_n852_), .B(KEYINPUT121), .Z(new_n853_));
  AOI21_X1  g652(.A(new_n851_), .B1(new_n843_), .B2(new_n853_), .ZN(G1347gat));
  NAND2_X1  g653(.A1(new_n637_), .A2(new_n532_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n855_), .A2(new_n516_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n250_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n577_), .B(new_n856_), .C1(new_n857_), .C2(new_n761_), .ZN(new_n858_));
  OAI21_X1  g657(.A(KEYINPUT62), .B1(new_n858_), .B2(KEYINPUT22), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT62), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n818_), .A2(new_n860_), .A3(new_n577_), .A4(new_n856_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n859_), .A2(G169gat), .A3(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT122), .ZN(new_n863_));
  OAI211_X1 g662(.A(KEYINPUT62), .B(new_n351_), .C1(new_n858_), .C2(KEYINPUT22), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n862_), .A2(new_n863_), .A3(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n863_), .B1(new_n862_), .B2(new_n864_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n865_), .A2(new_n866_), .ZN(G1348gat));
  AND2_X1   g666(.A1(new_n818_), .A2(new_n856_), .ZN(new_n868_));
  AOI21_X1  g667(.A(G176gat), .B1(new_n868_), .B2(new_n617_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n806_), .A2(new_n516_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n855_), .A2(new_n616_), .A3(new_n352_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n869_), .B1(new_n870_), .B2(new_n871_), .ZN(G1349gat));
  NOR2_X1   g671(.A1(new_n666_), .A2(new_n855_), .ZN(new_n873_));
  AOI21_X1  g672(.A(G183gat), .B1(new_n870_), .B2(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n666_), .A2(new_n346_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n868_), .B2(new_n875_), .ZN(G1350gat));
  NAND2_X1  g675(.A1(new_n868_), .A2(new_n659_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(G190gat), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n868_), .A2(new_n347_), .A3(new_n627_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1351gat));
  NAND2_X1  g679(.A1(new_n516_), .A2(new_n517_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n636_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n806_), .A2(new_n373_), .A3(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n577_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT123), .B(G197gat), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n885_), .B(new_n886_), .ZN(G1352gat));
  NAND2_X1  g686(.A1(new_n884_), .A2(new_n617_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g688(.A(new_n666_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n884_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT124), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n891_), .A2(KEYINPUT124), .ZN(new_n894_));
  OAI22_X1  g693(.A1(new_n893_), .A2(new_n894_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n895_));
  INV_X1    g694(.A(new_n894_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n896_), .A2(new_n897_), .A3(new_n892_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n895_), .A2(new_n898_), .ZN(G1354gat));
  NAND3_X1  g698(.A1(new_n884_), .A2(G218gat), .A3(new_n659_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT125), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n842_), .A2(new_n901_), .A3(new_n627_), .A4(new_n882_), .ZN(new_n902_));
  INV_X1    g701(.A(G218gat), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n901_), .B1(new_n884_), .B2(new_n627_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n900_), .B1(new_n904_), .B2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(KEYINPUT126), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT126), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n908_), .B(new_n900_), .C1(new_n904_), .C2(new_n905_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n907_), .A2(new_n909_), .ZN(G1355gat));
endmodule


