//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 1 1 0 0 0 1 1 1 0 0 1 1 1 1 0 0 0 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 1 1 0 1 1 1 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n803_, new_n804_, new_n805_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n881_, new_n882_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n203_));
  XOR2_X1   g002(.A(G71gat), .B(G78gat), .Z(new_n204_));
  OR2_X1    g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n204_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n205_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT66), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT7), .ZN(new_n210_));
  OAI211_X1 g009(.A(new_n209_), .B(new_n210_), .C1(G99gat), .C2(G106gat), .ZN(new_n211_));
  INV_X1    g010(.A(G99gat), .ZN(new_n212_));
  INV_X1    g011(.A(G106gat), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n212_), .B(new_n213_), .C1(KEYINPUT66), .C2(KEYINPUT7), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT6), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT6), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(G99gat), .A3(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n215_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT8), .ZN(new_n222_));
  INV_X1    g021(.A(G85gat), .ZN(new_n223_));
  INV_X1    g022(.A(G92gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G85gat), .A2(G92gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n221_), .A2(new_n222_), .A3(new_n228_), .ZN(new_n229_));
  AOI22_X1  g028(.A1(new_n220_), .A2(KEYINPUT67), .B1(new_n211_), .B2(new_n214_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT67), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n217_), .A2(new_n219_), .A3(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n227_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n229_), .B1(new_n233_), .B2(new_n222_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT10), .B(G99gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT64), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(new_n213_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT9), .ZN(new_n238_));
  INV_X1    g037(.A(new_n226_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n238_), .B(new_n225_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n225_), .A2(KEYINPUT65), .A3(KEYINPUT9), .A4(new_n226_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n241_), .A2(new_n220_), .A3(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n237_), .A2(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n208_), .B1(new_n234_), .B2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT70), .B(KEYINPUT12), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT71), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT71), .ZN(new_n249_));
  INV_X1    g048(.A(new_n247_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n243_), .B1(new_n236_), .B2(new_n213_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n218_), .B1(G99gat), .B2(G106gat), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n216_), .A2(KEYINPUT6), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT67), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n254_), .A2(new_n232_), .A3(new_n215_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(new_n228_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT8), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n251_), .B1(new_n257_), .B2(new_n229_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n249_), .B(new_n250_), .C1(new_n258_), .C2(new_n208_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n248_), .A2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n222_), .B1(new_n255_), .B2(new_n228_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n229_), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT69), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n264_), .B(new_n229_), .C1(new_n233_), .C2(new_n222_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(new_n245_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n205_), .B(KEYINPUT12), .C1(new_n207_), .C2(new_n206_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G230gat), .A2(G233gat), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n272_), .B1(new_n258_), .B2(new_n208_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n260_), .A2(new_n270_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT72), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  AOI22_X1  g075(.A1(new_n248_), .A2(new_n259_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n277_), .A2(KEYINPUT72), .A3(new_n273_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n271_), .B1(new_n246_), .B2(KEYINPUT68), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n258_), .A2(new_n208_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT68), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n279_), .B1(new_n282_), .B2(new_n246_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n276_), .A2(new_n278_), .A3(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G120gat), .B(G148gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT5), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G176gat), .B(G204gat), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n286_), .B(new_n287_), .Z(new_n288_));
  NAND2_X1  g087(.A1(new_n284_), .A2(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n288_), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n276_), .A2(new_n278_), .A3(new_n283_), .A4(new_n290_), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n289_), .A2(KEYINPUT13), .A3(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(KEYINPUT13), .B1(new_n289_), .B2(new_n291_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G229gat), .A2(G233gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G15gat), .B(G22gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT79), .ZN(new_n298_));
  INV_X1    g097(.A(G1gat), .ZN(new_n299_));
  INV_X1    g098(.A(G8gat), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT14), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT80), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n298_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G1gat), .B(G8gat), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n304_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G29gat), .B(G36gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G43gat), .B(G50gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n305_), .A2(new_n306_), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n309_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n296_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  XOR2_X1   g112(.A(KEYINPUT73), .B(KEYINPUT15), .Z(new_n314_));
  XNOR2_X1  g113(.A(new_n309_), .B(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n306_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n303_), .A2(new_n304_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n315_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(new_n310_), .A3(new_n295_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n313_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G113gat), .B(G141gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G169gat), .B(G197gat), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n321_), .B(new_n322_), .Z(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT81), .ZN(new_n325_));
  XOR2_X1   g124(.A(new_n320_), .B(new_n325_), .Z(new_n326_));
  NAND2_X1  g125(.A1(new_n294_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G127gat), .B(G134gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G113gat), .B(G120gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT83), .B(KEYINPUT84), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n330_), .A2(new_n331_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n333_), .A2(KEYINPUT85), .A3(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT85), .ZN(new_n336_));
  INV_X1    g135(.A(new_n334_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n336_), .B1(new_n337_), .B2(new_n332_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G71gat), .B(G99gat), .ZN(new_n339_));
  INV_X1    g138(.A(G43gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT30), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G227gat), .A2(G233gat), .ZN(new_n343_));
  INV_X1    g142(.A(G15gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n342_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G183gat), .A2(G190gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT23), .ZN(new_n348_));
  NOR2_X1   g147(.A1(G169gat), .A2(G176gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT24), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n348_), .A2(new_n351_), .ZN(new_n352_));
  AND2_X1   g151(.A1(G169gat), .A2(G176gat), .ZN(new_n353_));
  NOR3_X1   g152(.A1(new_n353_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT25), .B(G183gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT82), .B(G190gat), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n357_), .A2(KEYINPUT26), .ZN(new_n358_));
  NOR2_X1   g157(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n356_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n355_), .A2(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n348_), .B1(G183gat), .B2(new_n357_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(G169gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n361_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n342_), .A2(new_n345_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n346_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT87), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n367_), .B1(new_n346_), .B2(new_n368_), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n335_), .B(new_n338_), .C1(new_n370_), .C2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n371_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n338_), .A2(new_n335_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n373_), .A2(KEYINPUT87), .A3(new_n374_), .A4(new_n369_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n372_), .A2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT86), .B(KEYINPUT31), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n372_), .A2(new_n377_), .A3(new_n375_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(G155gat), .ZN(new_n382_));
  INV_X1    g181(.A(G162gat), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT88), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT88), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(G155gat), .A3(G162gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  AOI22_X1  g186(.A1(new_n387_), .A2(KEYINPUT1), .B1(new_n382_), .B2(new_n383_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n388_), .B1(KEYINPUT1), .B2(new_n387_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G141gat), .A2(G148gat), .ZN(new_n390_));
  INV_X1    g189(.A(G141gat), .ZN(new_n391_));
  INV_X1    g190(.A(G148gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n389_), .A2(new_n390_), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT89), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n390_), .A2(new_n395_), .ZN(new_n396_));
  OR2_X1    g195(.A1(new_n396_), .A2(KEYINPUT2), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n393_), .A2(KEYINPUT3), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(KEYINPUT2), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n393_), .A2(KEYINPUT3), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .A4(new_n400_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n401_), .B(new_n387_), .C1(G155gat), .C2(G162gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n394_), .A2(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT28), .B1(new_n403_), .B2(KEYINPUT29), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT28), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT29), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n394_), .A2(new_n405_), .A3(new_n406_), .A4(new_n402_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n403_), .A2(KEYINPUT29), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT90), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G211gat), .B(G218gat), .ZN(new_n410_));
  OR2_X1    g209(.A1(new_n410_), .A2(KEYINPUT92), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(KEYINPUT92), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(G204gat), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n414_), .A2(G197gat), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n414_), .A2(G197gat), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT21), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n416_), .B1(new_n415_), .B2(KEYINPUT91), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n418_), .B1(KEYINPUT91), .B2(new_n415_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n413_), .B(new_n417_), .C1(new_n419_), .C2(KEYINPUT21), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n419_), .A2(KEYINPUT21), .A3(new_n412_), .A4(new_n411_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n408_), .A2(new_n409_), .A3(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n409_), .B1(new_n408_), .B2(new_n422_), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n404_), .B(new_n407_), .C1(new_n423_), .C2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n424_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n404_), .A2(new_n407_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n408_), .A2(new_n409_), .A3(new_n422_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n426_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G228gat), .A2(G233gat), .ZN(new_n430_));
  INV_X1    g229(.A(G78gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(new_n213_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G22gat), .B(G50gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n425_), .A2(new_n429_), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n435_), .B1(new_n425_), .B2(new_n429_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n338_), .A2(new_n335_), .A3(new_n403_), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n394_), .B(new_n402_), .C1(new_n337_), .C2(new_n332_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(KEYINPUT4), .A3(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G225gat), .A2(G233gat), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT4), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n338_), .A2(new_n335_), .A3(new_n403_), .A4(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n441_), .A2(new_n443_), .A3(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G1gat), .B(G29gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(G85gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(KEYINPUT0), .B(G57gat), .ZN(new_n449_));
  XOR2_X1   g248(.A(new_n448_), .B(new_n449_), .Z(new_n450_));
  NAND3_X1  g249(.A1(new_n439_), .A2(new_n440_), .A3(new_n442_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n446_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT33), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n439_), .A2(new_n440_), .A3(new_n443_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n450_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT96), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n441_), .A2(new_n442_), .A3(new_n445_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n455_), .A2(KEYINPUT96), .A3(new_n456_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n446_), .A2(KEYINPUT33), .A3(new_n450_), .A4(new_n451_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G226gat), .A2(G233gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT19), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT20), .B1(new_n422_), .B2(new_n366_), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n352_), .A2(KEYINPUT93), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n352_), .A2(KEYINPUT93), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT26), .B(G190gat), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n354_), .B1(new_n356_), .B2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n467_), .A2(new_n468_), .A3(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n348_), .B1(G183gat), .B2(G190gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(new_n364_), .ZN(new_n473_));
  AOI22_X1  g272(.A1(new_n471_), .A2(new_n473_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n465_), .B1(new_n466_), .B2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G64gat), .B(G92gat), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT95), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  XOR2_X1   g277(.A(G8gat), .B(G36gat), .Z(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT20), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n483_), .B1(new_n422_), .B2(new_n366_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n465_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n471_), .A2(new_n420_), .A3(new_n421_), .A4(new_n473_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n484_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n475_), .A2(new_n482_), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n482_), .B1(new_n475_), .B2(new_n487_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n454_), .A2(new_n462_), .A3(new_n463_), .A4(new_n491_), .ZN(new_n492_));
  NOR3_X1   g291(.A1(new_n466_), .A2(new_n474_), .A3(new_n465_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n485_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n475_), .A2(new_n487_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n482_), .A2(KEYINPUT32), .ZN(new_n497_));
  MUX2_X1   g296(.A(new_n495_), .B(new_n496_), .S(new_n497_), .Z(new_n498_));
  INV_X1    g297(.A(new_n452_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n450_), .B1(new_n446_), .B2(new_n451_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n498_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n438_), .B1(new_n492_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n435_), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n426_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n427_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n503_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n500_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n425_), .A2(new_n429_), .A3(new_n435_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n506_), .A2(new_n507_), .A3(new_n508_), .A4(new_n452_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n482_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n510_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n511_), .A2(KEYINPUT27), .A3(new_n488_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT97), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT97), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n511_), .A2(new_n514_), .A3(KEYINPUT27), .A4(new_n488_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT27), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n516_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n513_), .A2(new_n515_), .A3(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n509_), .A2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n381_), .B1(new_n502_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n507_), .A2(new_n452_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n381_), .A2(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n518_), .A2(new_n438_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n327_), .B1(new_n520_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n305_), .A2(new_n306_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(new_n208_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G231gat), .A2(G233gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n527_), .B(new_n528_), .Z(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT17), .ZN(new_n531_));
  XOR2_X1   g330(.A(G127gat), .B(G155gat), .Z(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT16), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G183gat), .B(G211gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  OR3_X1    g334(.A1(new_n530_), .A2(new_n531_), .A3(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(KEYINPUT17), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n530_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G232gat), .A2(G233gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT34), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT35), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n315_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n545_), .B1(new_n266_), .B2(new_n245_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n234_), .A2(new_n245_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n309_), .ZN(new_n548_));
  OAI22_X1  g347(.A1(new_n547_), .A2(new_n548_), .B1(KEYINPUT35), .B2(new_n541_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n544_), .B1(new_n546_), .B2(new_n549_), .ZN(new_n550_));
  AOI22_X1  g349(.A1(new_n258_), .A2(new_n309_), .B1(new_n543_), .B2(new_n542_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n544_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n251_), .B1(new_n263_), .B2(new_n265_), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n551_), .B(new_n552_), .C1(new_n545_), .C2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G190gat), .B(G218gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G134gat), .B(G162gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n557_), .A2(KEYINPUT36), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n550_), .A2(new_n554_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n557_), .B(KEYINPUT36), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n561_), .B1(new_n550_), .B2(new_n554_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n560_), .B1(new_n563_), .B2(KEYINPUT76), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT77), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT37), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT76), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n562_), .A2(new_n567_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n564_), .A2(new_n565_), .A3(new_n566_), .A4(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n563_), .A2(KEYINPUT76), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n570_), .A2(new_n566_), .A3(new_n568_), .A4(new_n559_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(KEYINPUT77), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT74), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n559_), .B(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n550_), .A2(new_n554_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n561_), .ZN(new_n576_));
  AOI21_X1  g375(.A(KEYINPUT75), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT75), .ZN(new_n578_));
  AOI211_X1 g377(.A(new_n578_), .B(new_n561_), .C1(new_n550_), .C2(new_n554_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n566_), .B1(new_n574_), .B2(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n569_), .B1(new_n572_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT78), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT78), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n584_), .B(new_n569_), .C1(new_n572_), .C2(new_n581_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n539_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n525_), .A2(new_n586_), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n587_), .A2(KEYINPUT98), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(KEYINPUT98), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n590_), .A2(new_n299_), .A3(new_n521_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT100), .ZN(new_n592_));
  XOR2_X1   g391(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n593_));
  OR3_X1    g392(.A1(new_n591_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n564_), .A2(new_n568_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT101), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n596_), .B1(new_n520_), .B2(new_n524_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n539_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n327_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n597_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n299_), .B1(new_n601_), .B2(new_n521_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n591_), .B1(new_n593_), .B2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n592_), .B1(new_n591_), .B2(new_n593_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n594_), .A2(new_n603_), .A3(new_n604_), .ZN(G1324gat));
  INV_X1    g404(.A(new_n518_), .ZN(new_n606_));
  OAI21_X1  g405(.A(G8gat), .B1(new_n600_), .B2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT39), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n588_), .A2(new_n300_), .A3(new_n518_), .A4(new_n589_), .ZN(new_n609_));
  AOI21_X1  g408(.A(KEYINPUT102), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n608_), .A2(KEYINPUT102), .A3(new_n609_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n611_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n613_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(G1325gat));
  INV_X1    g415(.A(new_n381_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n590_), .A2(new_n344_), .A3(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(G15gat), .B1(new_n600_), .B2(new_n381_), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n619_), .B(KEYINPUT41), .Z(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(G1326gat));
  INV_X1    g420(.A(new_n438_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n622_), .A2(G22gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT104), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n590_), .A2(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(G22gat), .B1(new_n600_), .B2(new_n622_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT42), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT105), .Z(G1327gat));
  INV_X1    g428(.A(new_n596_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n630_), .A2(new_n598_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n525_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT107), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT107), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n525_), .A2(new_n634_), .A3(new_n631_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(G29gat), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(new_n637_), .A3(new_n521_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n520_), .A2(new_n524_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n639_), .A2(new_n583_), .A3(new_n585_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(KEYINPUT43), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT43), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n639_), .A2(new_n583_), .A3(new_n642_), .A4(new_n585_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n327_), .A2(new_n598_), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT44), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT44), .ZN(new_n647_));
  INV_X1    g446(.A(new_n645_), .ZN(new_n648_));
  AOI211_X1 g447(.A(new_n647_), .B(new_n648_), .C1(new_n641_), .C2(new_n643_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n646_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT106), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n650_), .A2(new_n651_), .A3(new_n521_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(G29gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n651_), .B1(new_n650_), .B2(new_n521_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n638_), .B1(new_n653_), .B2(new_n654_), .ZN(G1328gat));
  NOR2_X1   g454(.A1(new_n606_), .A2(G36gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n633_), .A2(new_n635_), .A3(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT45), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n644_), .A2(new_n645_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(new_n647_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT108), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n644_), .A2(KEYINPUT44), .A3(new_n645_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n660_), .A2(new_n661_), .A3(new_n518_), .A4(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(G36gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n661_), .B1(new_n650_), .B2(new_n518_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n658_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT46), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  OAI211_X1 g467(.A(KEYINPUT46), .B(new_n658_), .C1(new_n664_), .C2(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1329gat));
  NAND3_X1  g469(.A1(new_n650_), .A2(G43gat), .A3(new_n617_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n636_), .A2(new_n617_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(G43gat), .B2(new_n672_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g473(.A(G50gat), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n636_), .A2(new_n675_), .A3(new_n438_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n650_), .A2(KEYINPUT109), .A3(new_n438_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G50gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(KEYINPUT109), .B1(new_n650_), .B2(new_n438_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n676_), .B1(new_n678_), .B2(new_n679_), .ZN(G1331gat));
  NOR2_X1   g479(.A1(new_n294_), .A2(new_n326_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n597_), .A2(new_n598_), .A3(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n521_), .ZN(new_n683_));
  OAI21_X1  g482(.A(G57gat), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n639_), .A2(new_n681_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(new_n586_), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n683_), .A2(G57gat), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n684_), .B1(new_n686_), .B2(new_n687_), .ZN(G1332gat));
  OAI21_X1  g487(.A(G64gat), .B1(new_n682_), .B2(new_n606_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT110), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n691_), .A2(KEYINPUT48), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(KEYINPUT48), .ZN(new_n693_));
  OR3_X1    g492(.A1(new_n686_), .A2(G64gat), .A3(new_n606_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n692_), .A2(new_n693_), .A3(new_n694_), .ZN(G1333gat));
  OAI21_X1  g494(.A(G71gat), .B1(new_n682_), .B2(new_n381_), .ZN(new_n696_));
  XOR2_X1   g495(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n697_));
  XNOR2_X1  g496(.A(new_n696_), .B(new_n697_), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n381_), .A2(G71gat), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n698_), .B1(new_n686_), .B2(new_n699_), .ZN(G1334gat));
  OAI21_X1  g499(.A(G78gat), .B1(new_n682_), .B2(new_n622_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT50), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n438_), .A2(new_n431_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n686_), .B2(new_n703_), .ZN(G1335gat));
  NAND2_X1  g503(.A1(new_n685_), .A2(new_n631_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G85gat), .B1(new_n706_), .B2(new_n521_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n641_), .A2(KEYINPUT112), .A3(new_n643_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n681_), .A2(new_n539_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(KEYINPUT112), .B1(new_n641_), .B2(new_n643_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT113), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n521_), .A2(G85gat), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT114), .Z(new_n716_));
  AOI21_X1  g515(.A(new_n707_), .B1(new_n714_), .B2(new_n716_), .ZN(G1336gat));
  NAND3_X1  g516(.A1(new_n706_), .A2(new_n224_), .A3(new_n518_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n714_), .A2(new_n518_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n719_), .B2(new_n224_), .ZN(G1337gat));
  NAND3_X1  g519(.A1(new_n706_), .A2(new_n236_), .A3(new_n617_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n711_), .A2(new_n381_), .A3(new_n712_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n722_), .B2(new_n212_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g523(.A1(new_n706_), .A2(new_n213_), .A3(new_n438_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n709_), .A2(new_n622_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n213_), .B1(new_n644_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT52), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n727_), .A2(new_n728_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n725_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g531(.A1(new_n326_), .A2(new_n291_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT55), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n276_), .A2(new_n734_), .A3(new_n278_), .ZN(new_n735_));
  NAND4_X1  g534(.A1(new_n260_), .A2(KEYINPUT55), .A3(new_n270_), .A4(new_n273_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT116), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n277_), .A2(KEYINPUT116), .A3(KEYINPUT55), .A4(new_n273_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n735_), .A2(new_n738_), .A3(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(KEYINPUT115), .B1(new_n277_), .B2(new_n280_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n277_), .A2(KEYINPUT115), .A3(new_n280_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n271_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n288_), .B1(new_n740_), .B2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT56), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n738_), .A2(new_n739_), .ZN(new_n748_));
  AND4_X1   g547(.A1(KEYINPUT115), .A2(new_n260_), .A3(new_n270_), .A4(new_n280_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n272_), .B1(new_n749_), .B2(new_n741_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n748_), .A2(new_n750_), .A3(new_n735_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n751_), .A2(KEYINPUT56), .A3(new_n288_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n733_), .B1(new_n747_), .B2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n289_), .A2(new_n291_), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n313_), .A2(new_n323_), .A3(new_n319_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT117), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n318_), .A2(new_n310_), .A3(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n318_), .B2(new_n310_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n296_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  OR3_X1    g558(.A1(new_n311_), .A2(new_n296_), .A3(new_n312_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n755_), .B1(new_n761_), .B2(new_n324_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n754_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  OAI211_X1 g563(.A(KEYINPUT57), .B(new_n630_), .C1(new_n753_), .C2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n733_), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n751_), .A2(KEYINPUT56), .A3(new_n288_), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT56), .B1(new_n751_), .B2(new_n288_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n766_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n596_), .B1(new_n769_), .B2(new_n763_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n291_), .A2(new_n762_), .A3(KEYINPUT119), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT119), .B1(new_n291_), .B2(new_n762_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n774_), .B1(new_n747_), .B2(new_n752_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n583_), .B(new_n585_), .C1(new_n775_), .C2(KEYINPUT58), .ZN(new_n776_));
  INV_X1    g575(.A(new_n774_), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n777_), .B(KEYINPUT58), .C1(new_n767_), .C2(new_n768_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  OAI221_X1 g578(.A(new_n765_), .B1(new_n770_), .B2(new_n771_), .C1(new_n776_), .C2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n294_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n781_), .A2(new_n326_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n586_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT54), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n586_), .A2(new_n785_), .A3(new_n782_), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n780_), .A2(new_n539_), .B1(new_n784_), .B2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n523_), .A2(new_n521_), .A3(new_n617_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(G113gat), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n790_), .A3(new_n326_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n326_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n789_), .A2(KEYINPUT59), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT59), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n794_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n792_), .B1(new_n793_), .B2(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n791_), .B1(new_n796_), .B2(new_n790_), .ZN(G1340gat));
  INV_X1    g596(.A(G120gat), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n798_), .B1(new_n294_), .B2(KEYINPUT60), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n789_), .B(new_n799_), .C1(KEYINPUT60), .C2(new_n798_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n294_), .B1(new_n793_), .B2(new_n795_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n800_), .B1(new_n801_), .B2(new_n798_), .ZN(G1341gat));
  INV_X1    g601(.A(G127gat), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n789_), .A2(new_n803_), .A3(new_n598_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n539_), .B1(new_n793_), .B2(new_n795_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(new_n803_), .ZN(G1342gat));
  INV_X1    g605(.A(G134gat), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n789_), .A2(new_n807_), .A3(new_n596_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n583_), .A2(new_n585_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n809_), .B1(new_n793_), .B2(new_n795_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n808_), .B1(new_n810_), .B2(new_n807_), .ZN(G1343gat));
  OAI21_X1  g610(.A(new_n765_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n776_), .A2(new_n779_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n539_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n784_), .A2(new_n786_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n617_), .A2(new_n683_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n817_), .A2(new_n438_), .A3(new_n606_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n816_), .A2(new_n819_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n820_), .A2(new_n792_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(new_n391_), .ZN(G1344gat));
  NOR2_X1   g621(.A1(new_n820_), .A2(new_n294_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(new_n392_), .ZN(G1345gat));
  NOR2_X1   g623(.A1(new_n787_), .A2(new_n818_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n598_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(KEYINPUT61), .B(G155gat), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n826_), .B(new_n827_), .ZN(G1346gat));
  NAND4_X1  g627(.A1(new_n816_), .A2(new_n383_), .A3(new_n596_), .A4(new_n819_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n820_), .A2(new_n809_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(new_n383_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT120), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n829_), .B(KEYINPUT120), .C1(new_n830_), .C2(new_n383_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(G1347gat));
  NAND2_X1  g634(.A1(new_n522_), .A2(new_n622_), .ZN(new_n836_));
  NOR3_X1   g635(.A1(new_n836_), .A2(new_n792_), .A3(new_n606_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n838_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(KEYINPUT22), .B(G169gat), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT62), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT121), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n769_), .A2(new_n763_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n771_), .B1(new_n845_), .B2(new_n630_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847_));
  AOI211_X1 g646(.A(new_n847_), .B(new_n596_), .C1(new_n769_), .C2(new_n763_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  OR2_X1    g648(.A1(new_n775_), .A2(KEYINPUT58), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n850_), .A2(new_n583_), .A3(new_n585_), .A4(new_n778_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n598_), .B1(new_n849_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n786_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n785_), .B1(new_n586_), .B2(new_n782_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n837_), .B1(new_n852_), .B2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(G169gat), .B1(new_n842_), .B2(KEYINPUT121), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n844_), .B1(new_n856_), .B2(new_n858_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n839_), .A2(new_n857_), .A3(new_n843_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n841_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(KEYINPUT122), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT122), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n863_), .B(new_n841_), .C1(new_n859_), .C2(new_n860_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(G1348gat));
  NAND2_X1  g664(.A1(new_n816_), .A2(new_n518_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n836_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n781_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(G176gat), .ZN(G1349gat));
  AOI21_X1  g668(.A(new_n606_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n356_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n836_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n870_), .A2(new_n598_), .A3(new_n871_), .A4(new_n872_), .ZN(new_n873_));
  NOR4_X1   g672(.A1(new_n787_), .A2(new_n539_), .A3(new_n606_), .A4(new_n836_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n874_), .B2(G183gat), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT123), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT123), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n877_), .B(new_n873_), .C1(new_n874_), .C2(G183gat), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(G1350gat));
  NAND3_X1  g678(.A1(new_n867_), .A2(new_n469_), .A3(new_n596_), .ZN(new_n880_));
  INV_X1    g679(.A(G190gat), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n866_), .A2(new_n809_), .A3(new_n836_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n880_), .B1(new_n881_), .B2(new_n882_), .ZN(G1351gat));
  NOR2_X1   g682(.A1(new_n617_), .A2(new_n509_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n870_), .A2(new_n326_), .A3(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(KEYINPUT124), .A2(G197gat), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(KEYINPUT124), .B(G197gat), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n885_), .B2(new_n888_), .ZN(G1352gat));
  AND2_X1   g688(.A1(new_n870_), .A2(new_n884_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n781_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g691(.A(KEYINPUT63), .ZN(new_n893_));
  INV_X1    g692(.A(G211gat), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n598_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(KEYINPUT125), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n890_), .A2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n893_), .A2(new_n894_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n897_), .B(new_n898_), .ZN(G1354gat));
  NAND2_X1  g698(.A1(new_n890_), .A2(new_n596_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(KEYINPUT126), .B(G218gat), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n809_), .A2(new_n901_), .ZN(new_n902_));
  AOI22_X1  g701(.A1(new_n900_), .A2(new_n901_), .B1(new_n890_), .B2(new_n902_), .ZN(G1355gat));
endmodule


