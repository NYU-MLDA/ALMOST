//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 1 0 0 0 0 0 0 0 1 0 1 1 1 1 1 1 0 1 1 0 1 1 0 1 0 1 0 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n904_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_;
  XOR2_X1   g000(.A(G85gat), .B(G92gat), .Z(new_n202_));
  NOR2_X1   g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT7), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT67), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT67), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n203_), .A2(new_n207_), .A3(new_n204_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT66), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  INV_X1    g011(.A(G99gat), .ZN(new_n213_));
  INV_X1    g012(.A(G106gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n212_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT66), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n216_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n211_), .A2(new_n215_), .A3(new_n217_), .A4(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n202_), .B1(new_n209_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT68), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT8), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  NOR4_X1   g022(.A1(KEYINPUT67), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n207_), .B1(new_n203_), .B2(new_n204_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n211_), .A2(new_n217_), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n215_), .A2(new_n218_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n221_), .A2(new_n222_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(KEYINPUT68), .A2(KEYINPUT8), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n229_), .A2(new_n202_), .A3(new_n230_), .A4(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT9), .ZN(new_n233_));
  INV_X1    g032(.A(G85gat), .ZN(new_n234_));
  INV_X1    g033(.A(G92gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n233_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  OAI211_X1 g035(.A(KEYINPUT65), .B(new_n236_), .C1(new_n202_), .C2(new_n233_), .ZN(new_n237_));
  XOR2_X1   g036(.A(KEYINPUT10), .B(G99gat), .Z(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(new_n214_), .ZN(new_n239_));
  OR4_X1    g038(.A1(KEYINPUT65), .A2(new_n233_), .A3(new_n234_), .A4(new_n235_), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n237_), .A2(new_n239_), .A3(new_n228_), .A4(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n223_), .A2(new_n232_), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT69), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n223_), .A2(new_n232_), .A3(new_n244_), .A4(new_n241_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G57gat), .B(G64gat), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n247_), .A2(KEYINPUT11), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(KEYINPUT11), .ZN(new_n249_));
  XOR2_X1   g048(.A(G71gat), .B(G78gat), .Z(new_n250_));
  NAND3_X1  g049(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n249_), .A2(new_n250_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n246_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n253_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n243_), .A2(new_n255_), .A3(new_n245_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G230gat), .A2(G233gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT64), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT12), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n256_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n259_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n253_), .B(KEYINPUT70), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n264_), .A2(KEYINPUT12), .A3(new_n242_), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n262_), .A2(new_n254_), .A3(new_n263_), .A4(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n260_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G120gat), .B(G148gat), .ZN(new_n268_));
  INV_X1    g067(.A(G204gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT5), .ZN(new_n271_));
  INV_X1    g070(.A(G176gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n267_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n260_), .A2(new_n266_), .A3(new_n273_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  AND2_X1   g076(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n278_));
  NOR2_X1   g077(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n277_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n280_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT2), .ZN(new_n283_));
  INV_X1    g082(.A(G141gat), .ZN(new_n284_));
  INV_X1    g083(.A(G148gat), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n283_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT3), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n287_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n288_));
  OAI21_X1  g087(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n289_));
  NAND3_X1  g088(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n290_));
  NAND4_X1  g089(.A1(new_n286_), .A2(new_n288_), .A3(new_n289_), .A4(new_n290_), .ZN(new_n291_));
  AND2_X1   g090(.A1(G155gat), .A2(G162gat), .ZN(new_n292_));
  NOR2_X1   g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n291_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT88), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT1), .ZN(new_n298_));
  AOI22_X1  g097(.A1(new_n294_), .A2(new_n298_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n299_));
  AOI22_X1  g098(.A1(new_n292_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n297_), .A2(new_n301_), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n302_), .A2(KEYINPUT29), .ZN(new_n303_));
  XOR2_X1   g102(.A(G78gat), .B(G106gat), .Z(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n302_), .A2(KEYINPUT29), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G211gat), .B(G218gat), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n308_), .A2(KEYINPUT21), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(KEYINPUT21), .ZN(new_n310_));
  XOR2_X1   g109(.A(G197gat), .B(G204gat), .Z(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n310_), .A2(new_n311_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n307_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(G233gat), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT89), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n317_), .A2(G228gat), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(G228gat), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n316_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n315_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G22gat), .B(G50gat), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n323_), .B(KEYINPUT28), .Z(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n314_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n326_), .B1(new_n302_), .B2(KEYINPUT29), .ZN(new_n327_));
  INV_X1    g126(.A(new_n321_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n322_), .A2(new_n325_), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n325_), .B1(new_n322_), .B2(new_n329_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n306_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n332_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n334_), .A2(new_n330_), .A3(new_n305_), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT87), .B(KEYINPUT31), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G15gat), .B(G43gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(G71gat), .B(G99gat), .Z(new_n340_));
  XOR2_X1   g139(.A(new_n339_), .B(new_n340_), .Z(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT86), .B(KEYINPUT30), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT26), .B(G190gat), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT82), .ZN(new_n345_));
  INV_X1    g144(.A(G183gat), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n345_), .B1(new_n346_), .B2(KEYINPUT25), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT25), .B(G183gat), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n344_), .B(new_n347_), .C1(new_n348_), .C2(new_n345_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT24), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n350_), .B1(G169gat), .B2(G176gat), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n351_), .B1(G169gat), .B2(G176gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n349_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT83), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G183gat), .A2(G190gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT23), .ZN(new_n357_));
  NOR2_X1   g156(.A1(G169gat), .A2(G176gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(new_n350_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n349_), .A2(KEYINPUT83), .A3(new_n352_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n355_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n357_), .B1(G183gat), .B2(G190gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G169gat), .A2(G176gat), .ZN(new_n364_));
  INV_X1    g163(.A(G169gat), .ZN(new_n365_));
  OAI21_X1  g164(.A(KEYINPUT22), .B1(new_n365_), .B2(KEYINPUT84), .ZN(new_n366_));
  OR2_X1    g165(.A1(new_n365_), .A2(KEYINPUT22), .ZN(new_n367_));
  OAI211_X1 g166(.A(new_n272_), .B(new_n366_), .C1(new_n367_), .C2(KEYINPUT84), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n363_), .A2(new_n364_), .A3(new_n368_), .ZN(new_n369_));
  AND3_X1   g168(.A1(new_n362_), .A2(KEYINPUT85), .A3(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(KEYINPUT85), .B1(new_n362_), .B2(new_n369_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n343_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n362_), .A2(new_n369_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT85), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n362_), .A2(new_n369_), .A3(KEYINPUT85), .ZN(new_n376_));
  INV_X1    g175(.A(new_n343_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n372_), .A2(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G127gat), .B(G134gat), .ZN(new_n380_));
  INV_X1    g179(.A(G113gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(G120gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n379_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G227gat), .A2(G233gat), .ZN(new_n385_));
  INV_X1    g184(.A(G120gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n382_), .B(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n372_), .A2(new_n378_), .A3(new_n387_), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n384_), .A2(new_n385_), .A3(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n385_), .B1(new_n384_), .B2(new_n388_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n342_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n372_), .A2(new_n378_), .A3(new_n387_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n387_), .B1(new_n372_), .B2(new_n378_), .ZN(new_n393_));
  OAI211_X1 g192(.A(G227gat), .B(G233gat), .C1(new_n392_), .C2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n384_), .A2(new_n385_), .A3(new_n388_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n394_), .A2(new_n395_), .A3(new_n341_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n391_), .A2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n326_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G226gat), .A2(G233gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT19), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n344_), .A2(new_n348_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT90), .ZN(new_n403_));
  AND3_X1   g202(.A1(new_n364_), .A2(new_n403_), .A3(KEYINPUT24), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n403_), .B1(new_n364_), .B2(KEYINPUT24), .ZN(new_n405_));
  OR2_X1    g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  OAI211_X1 g205(.A(KEYINPUT91), .B(new_n402_), .C1(new_n406_), .C2(new_n358_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT91), .ZN(new_n408_));
  INV_X1    g207(.A(new_n402_), .ZN(new_n409_));
  NOR3_X1   g208(.A1(new_n404_), .A2(new_n405_), .A3(new_n358_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n408_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n407_), .A2(new_n411_), .A3(new_n360_), .ZN(new_n412_));
  XOR2_X1   g211(.A(KEYINPUT22), .B(G169gat), .Z(new_n413_));
  OAI211_X1 g212(.A(new_n363_), .B(new_n364_), .C1(G176gat), .C2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  OAI211_X1 g214(.A(KEYINPUT20), .B(new_n401_), .C1(new_n415_), .C2(new_n314_), .ZN(new_n416_));
  OR2_X1    g215(.A1(new_n398_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n375_), .A2(new_n376_), .A3(new_n326_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n415_), .A2(new_n314_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT92), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n415_), .A2(KEYINPUT92), .A3(new_n314_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n418_), .A2(new_n421_), .A3(KEYINPUT20), .A4(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT93), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n423_), .A2(new_n424_), .A3(new_n400_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n424_), .B1(new_n423_), .B2(new_n400_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n417_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT18), .B(G64gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(G92gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G8gat), .B(G36gat), .ZN(new_n430_));
  XOR2_X1   g229(.A(new_n429_), .B(new_n430_), .Z(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n427_), .A2(new_n432_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n417_), .B(new_n431_), .C1(new_n425_), .C2(new_n426_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n302_), .A2(new_n383_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n387_), .A2(new_n301_), .A3(new_n297_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G225gat), .A2(G233gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT94), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(KEYINPUT0), .B(G57gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(G85gat), .ZN(new_n442_));
  XOR2_X1   g241(.A(G1gat), .B(G29gat), .Z(new_n443_));
  XOR2_X1   g242(.A(new_n442_), .B(new_n443_), .Z(new_n444_));
  NAND3_X1  g243(.A1(new_n440_), .A2(KEYINPUT95), .A3(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n438_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n435_), .A2(KEYINPUT4), .A3(new_n436_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n447_), .B1(KEYINPUT4), .B2(new_n435_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n445_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(KEYINPUT95), .B1(new_n440_), .B2(new_n444_), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n447_), .B(new_n439_), .C1(KEYINPUT4), .C2(new_n435_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n437_), .A2(new_n438_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n444_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT33), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n433_), .A2(new_n434_), .A3(new_n451_), .A4(new_n456_), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n431_), .A2(KEYINPUT32), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT96), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n415_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n412_), .A2(KEYINPUT96), .A3(new_n414_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n460_), .A2(new_n326_), .A3(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT20), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT97), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n398_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n462_), .A2(KEYINPUT97), .A3(KEYINPUT20), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n401_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n423_), .A2(new_n400_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n458_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n452_), .A2(new_n453_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n444_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n455_), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n469_), .B(new_n472_), .C1(new_n427_), .C2(new_n458_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n397_), .B1(new_n457_), .B2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT27), .B1(new_n433_), .B2(new_n434_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n432_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n476_), .A2(KEYINPUT27), .A3(new_n434_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT98), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n472_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n471_), .A2(KEYINPUT98), .A3(new_n455_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n394_), .A2(new_n395_), .A3(new_n341_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n341_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n336_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n333_), .A2(new_n335_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n391_), .A2(new_n396_), .A3(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n482_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n336_), .A2(new_n474_), .B1(new_n478_), .B2(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(G1gat), .A2(G8gat), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT73), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G1gat), .A2(G8gat), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  AND2_X1   g293(.A1(G1gat), .A2(G8gat), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT73), .B1(new_n495_), .B2(new_n490_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n493_), .A2(KEYINPUT14), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT72), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  OR2_X1    g299(.A1(G15gat), .A2(G22gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G15gat), .A2(G22gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n493_), .A2(KEYINPUT72), .A3(KEYINPUT14), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n500_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n497_), .A2(new_n505_), .ZN(new_n506_));
  AOI22_X1  g305(.A1(new_n499_), .A2(new_n498_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n507_));
  AOI22_X1  g306(.A1(new_n507_), .A2(new_n504_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  AND2_X1   g308(.A1(G29gat), .A2(G36gat), .ZN(new_n510_));
  NOR2_X1   g309(.A1(G29gat), .A2(G36gat), .ZN(new_n511_));
  OAI21_X1  g310(.A(G43gat), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(G29gat), .ZN(new_n513_));
  INV_X1    g312(.A(G36gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(G43gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G29gat), .A2(G36gat), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n515_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n512_), .A2(new_n518_), .A3(G50gat), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(G50gat), .B1(new_n512_), .B2(new_n518_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT15), .ZN(new_n522_));
  NOR3_X1   g321(.A1(new_n520_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n512_), .A2(new_n518_), .ZN(new_n524_));
  INV_X1    g323(.A(G50gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(KEYINPUT15), .B1(new_n526_), .B2(new_n519_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n509_), .B1(new_n523_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT77), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G229gat), .A2(G233gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n497_), .B(new_n505_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n520_), .A2(new_n521_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT77), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n509_), .B(new_n534_), .C1(new_n523_), .C2(new_n527_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n529_), .A2(new_n530_), .A3(new_n533_), .A4(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n531_), .B(new_n532_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n530_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n536_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT78), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G113gat), .B(G141gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(new_n365_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(G197gat), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n545_), .B(KEYINPUT79), .Z(new_n546_));
  NAND3_X1  g345(.A1(new_n536_), .A2(new_n539_), .A3(KEYINPUT78), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n542_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT80), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n536_), .A2(new_n539_), .A3(new_n545_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n542_), .A2(KEYINPUT80), .A3(new_n546_), .A4(new_n547_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n550_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT81), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT81), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n550_), .A2(new_n555_), .A3(new_n551_), .A4(new_n552_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT99), .B1(new_n489_), .B2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n457_), .A2(new_n473_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n397_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n560_), .A2(new_n561_), .A3(new_n336_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n485_), .A2(new_n487_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n482_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT27), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n423_), .A2(new_n400_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(KEYINPUT93), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n423_), .A2(new_n424_), .A3(new_n400_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n431_), .B1(new_n569_), .B2(new_n417_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n434_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n565_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n476_), .A2(KEYINPUT27), .A3(new_n434_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n563_), .A2(new_n564_), .A3(new_n572_), .A4(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n562_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT99), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n575_), .A2(new_n576_), .A3(new_n557_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n282_), .B1(new_n559_), .B2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n246_), .A2(new_n532_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n242_), .B1(new_n523_), .B2(new_n527_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G232gat), .A2(G233gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT34), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n579_), .B(new_n580_), .C1(KEYINPUT35), .C2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(KEYINPUT35), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n583_), .A2(new_n584_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(G134gat), .ZN(new_n589_));
  INV_X1    g388(.A(G162gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  OAI22_X1  g391(.A1(new_n586_), .A2(new_n587_), .B1(KEYINPUT36), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n587_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n591_), .B(KEYINPUT36), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n594_), .A2(new_n596_), .A3(new_n585_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT37), .ZN(new_n598_));
  AND3_X1   g397(.A1(new_n593_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n598_), .B1(new_n593_), .B2(new_n597_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n509_), .B(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(new_n264_), .ZN(new_n603_));
  XOR2_X1   g402(.A(KEYINPUT75), .B(KEYINPUT17), .Z(new_n604_));
  XOR2_X1   g403(.A(G127gat), .B(G155gat), .Z(new_n605_));
  XNOR2_X1  g404(.A(G183gat), .B(G211gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n603_), .A2(new_n604_), .A3(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n602_), .B(new_n253_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n609_), .B(KEYINPUT17), .Z(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n610_), .A2(new_n613_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n599_), .A2(new_n600_), .A3(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT76), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n578_), .A2(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT100), .ZN(new_n618_));
  INV_X1    g417(.A(G1gat), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n618_), .A2(new_n619_), .A3(new_n482_), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n620_), .A2(KEYINPUT38), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n593_), .A2(new_n597_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n575_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT101), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n614_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n282_), .A2(new_n558_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n626_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G1gat), .B1(new_n630_), .B2(new_n564_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n620_), .A2(KEYINPUT38), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n621_), .A2(new_n631_), .A3(new_n632_), .ZN(G1324gat));
  INV_X1    g432(.A(G8gat), .ZN(new_n634_));
  INV_X1    g433(.A(new_n478_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n618_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT39), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n629_), .A2(new_n635_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n638_), .B2(G8gat), .ZN(new_n639_));
  AOI211_X1 g438(.A(KEYINPUT39), .B(new_n634_), .C1(new_n629_), .C2(new_n635_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n636_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT40), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n636_), .B(KEYINPUT40), .C1(new_n639_), .C2(new_n640_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(G1325gat));
  OR3_X1    g444(.A1(new_n617_), .A2(G15gat), .A3(new_n561_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n629_), .A2(new_n397_), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n647_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n648_));
  AOI21_X1  g447(.A(KEYINPUT41), .B1(new_n647_), .B2(G15gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n646_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  OAI211_X1 g451(.A(KEYINPUT102), .B(new_n646_), .C1(new_n648_), .C2(new_n649_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1326gat));
  XNOR2_X1  g453(.A(new_n486_), .B(KEYINPUT103), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G22gat), .B1(new_n630_), .B2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT42), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n656_), .A2(G22gat), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n658_), .B1(new_n617_), .B2(new_n659_), .ZN(G1327gat));
  INV_X1    g459(.A(KEYINPUT43), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n599_), .A2(new_n600_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n661_), .B1(new_n575_), .B2(new_n663_), .ZN(new_n664_));
  AOI211_X1 g463(.A(KEYINPUT43), .B(new_n662_), .C1(new_n562_), .C2(new_n574_), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n614_), .B(new_n628_), .C1(new_n664_), .C2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(KEYINPUT43), .B1(new_n489_), .B2(new_n662_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n575_), .A2(new_n661_), .A3(new_n663_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n671_), .A2(KEYINPUT44), .A3(new_n614_), .A4(new_n628_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n668_), .A2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n673_), .A2(G29gat), .A3(new_n482_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n623_), .A2(new_n627_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n578_), .A2(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n513_), .B1(new_n676_), .B2(new_n564_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n674_), .A2(new_n677_), .ZN(G1328gat));
  NAND3_X1  g477(.A1(new_n668_), .A2(new_n635_), .A3(new_n672_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(G36gat), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT104), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n578_), .A2(new_n514_), .A3(new_n635_), .A4(new_n675_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT45), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n679_), .A2(KEYINPUT104), .A3(G36gat), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n682_), .A2(new_n684_), .A3(new_n685_), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n686_), .A2(KEYINPUT105), .A3(KEYINPUT46), .ZN(new_n687_));
  AOI21_X1  g486(.A(KEYINPUT46), .B1(new_n686_), .B2(KEYINPUT105), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1329gat));
  NAND3_X1  g488(.A1(new_n673_), .A2(G43gat), .A3(new_n397_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n516_), .B1(new_n676_), .B2(new_n561_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g492(.A1(new_n673_), .A2(KEYINPUT106), .A3(new_n486_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n668_), .A2(new_n486_), .A3(new_n672_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n694_), .A2(G50gat), .A3(new_n697_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n698_), .A2(KEYINPUT107), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n698_), .A2(KEYINPUT107), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n655_), .A2(new_n525_), .ZN(new_n701_));
  OAI22_X1  g500(.A1(new_n699_), .A2(new_n700_), .B1(new_n676_), .B2(new_n701_), .ZN(G1331gat));
  NAND2_X1  g501(.A1(new_n282_), .A2(new_n558_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n489_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(new_n616_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G57gat), .B1(new_n706_), .B2(new_n482_), .ZN(new_n707_));
  AND4_X1   g506(.A1(new_n627_), .A2(new_n626_), .A3(new_n558_), .A4(new_n282_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n708_), .A2(new_n482_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n707_), .B1(new_n709_), .B2(G57gat), .ZN(G1332gat));
  INV_X1    g509(.A(G64gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n711_), .B1(new_n708_), .B2(new_n635_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT48), .Z(new_n713_));
  NAND3_X1  g512(.A1(new_n706_), .A2(new_n711_), .A3(new_n635_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1333gat));
  INV_X1    g514(.A(G71gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n708_), .B2(new_n397_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT49), .Z(new_n718_));
  NAND3_X1  g517(.A1(new_n706_), .A2(new_n716_), .A3(new_n397_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1334gat));
  INV_X1    g519(.A(G78gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n721_), .B1(new_n708_), .B2(new_n655_), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT50), .Z(new_n723_));
  NAND3_X1  g522(.A1(new_n706_), .A2(new_n721_), .A3(new_n655_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1335gat));
  NAND2_X1  g524(.A1(new_n704_), .A2(new_n675_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n726_), .A2(G85gat), .A3(new_n564_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n703_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n614_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(new_n482_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n727_), .B1(new_n731_), .B2(G85gat), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT108), .Z(G1336gat));
  INV_X1    g532(.A(new_n726_), .ZN(new_n734_));
  AOI21_X1  g533(.A(G92gat), .B1(new_n734_), .B2(new_n635_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n729_), .A2(new_n478_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n736_), .B2(G92gat), .ZN(G1337gat));
  NAND2_X1  g536(.A1(new_n730_), .A2(new_n397_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n397_), .A2(new_n238_), .ZN(new_n739_));
  AOI22_X1  g538(.A1(new_n738_), .A2(G99gat), .B1(new_n734_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n741_), .A2(KEYINPUT109), .A3(KEYINPUT51), .ZN(new_n742_));
  AOI21_X1  g541(.A(KEYINPUT109), .B1(new_n741_), .B2(KEYINPUT51), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n741_), .A2(KEYINPUT110), .A3(KEYINPUT51), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT51), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n740_), .B2(new_n746_), .ZN(new_n747_));
  OAI22_X1  g546(.A1(new_n742_), .A2(new_n743_), .B1(new_n744_), .B2(new_n747_), .ZN(G1338gat));
  INV_X1    g547(.A(KEYINPUT111), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n749_), .B1(new_n729_), .B2(new_n336_), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n728_), .A2(KEYINPUT111), .A3(new_n614_), .A4(new_n486_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(G106gat), .A3(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT52), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n750_), .A2(new_n754_), .A3(G106gat), .A4(new_n751_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n734_), .A2(new_n214_), .A3(new_n486_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT53), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT53), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n756_), .A2(new_n760_), .A3(new_n757_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1339gat));
  NAND2_X1  g561(.A1(new_n281_), .A2(new_n558_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n600_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n593_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n764_), .A2(new_n627_), .A3(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(KEYINPUT54), .B1(new_n763_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT54), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n615_), .A2(new_n281_), .A3(new_n768_), .A4(new_n558_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n276_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n545_), .B1(new_n537_), .B2(new_n530_), .ZN(new_n772_));
  OR2_X1    g571(.A1(new_n772_), .A2(KEYINPUT112), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n529_), .A2(new_n538_), .A3(new_n533_), .A4(new_n535_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(KEYINPUT112), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n773_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n551_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT113), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n776_), .A2(KEYINPUT113), .A3(new_n551_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n771_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n255_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n782_), .B1(new_n261_), .B2(new_n256_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n263_), .B1(new_n783_), .B2(new_n265_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n266_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n262_), .A2(new_n254_), .A3(new_n265_), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n787_), .A2(new_n785_), .A3(new_n259_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n786_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT56), .B1(new_n790_), .B2(new_n274_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT56), .ZN(new_n792_));
  AOI211_X1 g591(.A(new_n792_), .B(new_n273_), .C1(new_n786_), .C2(new_n789_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n781_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT58), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n662_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  OAI211_X1 g595(.A(KEYINPUT58), .B(new_n781_), .C1(new_n791_), .C2(new_n793_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  AND4_X1   g598(.A1(new_n263_), .A2(new_n262_), .A3(new_n254_), .A4(new_n265_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n787_), .A2(new_n259_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(KEYINPUT55), .B2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n274_), .B1(new_n802_), .B2(new_n788_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n792_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n790_), .A2(KEYINPUT56), .A3(new_n274_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n806_), .A2(KEYINPUT114), .A3(KEYINPUT58), .A4(new_n781_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n796_), .A2(new_n799_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n779_), .A2(new_n780_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n277_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n791_), .A2(new_n793_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n557_), .A2(new_n276_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n810_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n813_), .A2(KEYINPUT57), .A3(new_n623_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n815_));
  INV_X1    g614(.A(new_n810_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n771_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n816_), .B1(new_n806_), .B2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n815_), .B1(new_n818_), .B2(new_n622_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n808_), .A2(new_n814_), .A3(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n770_), .B1(new_n820_), .B2(new_n614_), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n635_), .A2(new_n564_), .A3(new_n485_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n821_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n381_), .B1(new_n825_), .B2(new_n558_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n826_), .A2(KEYINPUT115), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n826_), .A2(KEYINPUT115), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n823_), .A2(KEYINPUT116), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT116), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT59), .B1(new_n822_), .B2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT57), .B1(new_n813_), .B2(new_n623_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n818_), .A2(new_n815_), .A3(new_n622_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n627_), .B1(new_n834_), .B2(new_n808_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n829_), .B(new_n831_), .C1(new_n835_), .C2(new_n770_), .ZN(new_n836_));
  OAI21_X1  g635(.A(KEYINPUT59), .B1(new_n821_), .B2(new_n823_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n558_), .A2(new_n381_), .ZN(new_n839_));
  AOI211_X1 g638(.A(new_n827_), .B(new_n828_), .C1(new_n838_), .C2(new_n839_), .ZN(G1340gat));
  NAND3_X1  g639(.A1(new_n836_), .A2(new_n282_), .A3(new_n837_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT117), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n836_), .A2(new_n837_), .A3(new_n843_), .A4(new_n282_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n842_), .A2(G120gat), .A3(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n386_), .B1(new_n281_), .B2(KEYINPUT60), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n824_), .B(new_n846_), .C1(KEYINPUT60), .C2(new_n386_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(KEYINPUT118), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n845_), .A2(new_n850_), .A3(new_n847_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n851_), .ZN(G1341gat));
  OAI21_X1  g651(.A(G127gat), .B1(new_n614_), .B2(KEYINPUT119), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n838_), .B(new_n853_), .C1(KEYINPUT119), .C2(G127gat), .ZN(new_n854_));
  INV_X1    g653(.A(G127gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n825_), .B2(new_n614_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n854_), .A2(new_n856_), .ZN(G1342gat));
  AOI21_X1  g656(.A(G134gat), .B1(new_n824_), .B2(new_n622_), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n838_), .A2(new_n663_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n858_), .B1(new_n859_), .B2(G134gat), .ZN(G1343gat));
  NOR2_X1   g659(.A1(new_n821_), .A2(new_n487_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n635_), .A2(new_n564_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(new_n558_), .ZN(new_n864_));
  XOR2_X1   g663(.A(KEYINPUT120), .B(G141gat), .Z(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1344gat));
  NOR2_X1   g665(.A1(new_n863_), .A2(new_n281_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(new_n285_), .ZN(G1345gat));
  NOR2_X1   g667(.A1(new_n863_), .A2(new_n614_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(KEYINPUT61), .B(G155gat), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(KEYINPUT121), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n869_), .B(new_n871_), .ZN(G1346gat));
  NOR3_X1   g671(.A1(new_n863_), .A2(new_n590_), .A3(new_n662_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n861_), .A2(new_n622_), .A3(new_n862_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n873_), .B1(new_n590_), .B2(new_n874_), .ZN(G1347gat));
  NOR2_X1   g674(.A1(new_n478_), .A2(new_n482_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n397_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(new_n558_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(KEYINPUT122), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n879_), .A2(new_n656_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n821_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n365_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT62), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(KEYINPUT123), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT123), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n882_), .A2(new_n886_), .A3(new_n883_), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n885_), .B(new_n887_), .C1(new_n883_), .C2(new_n882_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n821_), .A2(new_n655_), .A3(new_n877_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n558_), .A2(new_n413_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(KEYINPUT124), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n888_), .A2(new_n892_), .ZN(G1348gat));
  NOR2_X1   g692(.A1(new_n821_), .A2(new_n486_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n877_), .ZN(new_n895_));
  AND4_X1   g694(.A1(G176gat), .A2(new_n894_), .A3(new_n282_), .A4(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(G176gat), .B1(new_n889_), .B2(new_n282_), .ZN(new_n897_));
  OR2_X1    g696(.A1(new_n897_), .A2(KEYINPUT125), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(KEYINPUT125), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n896_), .B1(new_n898_), .B2(new_n899_), .ZN(G1349gat));
  NAND3_X1  g699(.A1(new_n894_), .A2(new_n627_), .A3(new_n895_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n614_), .A2(new_n348_), .ZN(new_n902_));
  AOI22_X1  g701(.A1(new_n901_), .A2(new_n346_), .B1(new_n889_), .B2(new_n902_), .ZN(G1350gat));
  NAND3_X1  g702(.A1(new_n889_), .A2(new_n622_), .A3(new_n344_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n889_), .A2(new_n663_), .ZN(new_n905_));
  INV_X1    g704(.A(G190gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n904_), .B1(new_n905_), .B2(new_n906_), .ZN(G1351gat));
  NAND2_X1  g706(.A1(new_n861_), .A2(new_n876_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n908_), .A2(new_n558_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(KEYINPUT126), .B(G197gat), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n909_), .B2(new_n912_), .ZN(G1352gat));
  NOR2_X1   g712(.A1(new_n908_), .A2(new_n281_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(new_n269_), .ZN(G1353gat));
  INV_X1    g714(.A(new_n908_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n627_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n918_));
  AND2_X1   g717(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n917_), .A2(new_n918_), .A3(new_n919_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n920_), .B1(new_n917_), .B2(new_n918_), .ZN(G1354gat));
  AOI21_X1  g720(.A(G218gat), .B1(new_n916_), .B2(new_n622_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n663_), .A2(G218gat), .ZN(new_n923_));
  XOR2_X1   g722(.A(new_n923_), .B(KEYINPUT127), .Z(new_n924_));
  AOI21_X1  g723(.A(new_n922_), .B1(new_n916_), .B2(new_n924_), .ZN(G1355gat));
endmodule


