//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 1 0 0 1 0 1 1 0 0 1 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1 0 0 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0 1 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n927_, new_n928_, new_n929_,
    new_n931_, new_n932_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n940_, new_n941_, new_n943_, new_n944_, new_n945_,
    new_n947_, new_n948_;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n203_));
  XOR2_X1   g002(.A(KEYINPUT65), .B(G92gat), .Z(new_n204_));
  INV_X1    g003(.A(G85gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(new_n203_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(G85gat), .A2(G92gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT9), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G85gat), .A2(G92gat), .ZN(new_n209_));
  OAI211_X1 g008(.A(new_n206_), .B(new_n207_), .C1(new_n208_), .C2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT6), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G99gat), .A3(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(KEYINPUT10), .B(G99gat), .Z(new_n216_));
  INV_X1    g015(.A(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n210_), .A2(new_n215_), .A3(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT8), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT67), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n213_), .B1(G99gat), .B2(G106gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n211_), .A2(KEYINPUT6), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n222_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n212_), .A2(new_n214_), .A3(KEYINPUT67), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT7), .ZN(new_n227_));
  INV_X1    g026(.A(G99gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n228_), .A3(new_n217_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n230_));
  AND3_X1   g029(.A1(new_n229_), .A2(KEYINPUT68), .A3(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(KEYINPUT68), .B1(new_n229_), .B2(new_n230_), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n225_), .B(new_n226_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n207_), .A2(new_n209_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n221_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n215_), .A2(new_n230_), .A3(new_n229_), .ZN(new_n237_));
  XOR2_X1   g036(.A(KEYINPUT66), .B(KEYINPUT8), .Z(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(new_n235_), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT69), .B1(new_n236_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n212_), .A2(new_n214_), .A3(KEYINPUT67), .ZN(new_n243_));
  AOI21_X1  g042(.A(KEYINPUT67), .B1(new_n212_), .B2(new_n214_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n246_));
  INV_X1    g045(.A(new_n230_), .ZN(new_n247_));
  NOR3_X1   g046(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n246_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n229_), .A2(KEYINPUT68), .A3(new_n230_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n234_), .B1(new_n245_), .B2(new_n251_), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n242_), .B(new_n239_), .C1(new_n252_), .C2(new_n221_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n220_), .B1(new_n241_), .B2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G57gat), .B(G64gat), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n255_), .A2(KEYINPUT11), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(KEYINPUT11), .ZN(new_n257_));
  XOR2_X1   g056(.A(G71gat), .B(G78gat), .Z(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n257_), .A2(new_n258_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT12), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n239_), .B1(new_n252_), .B2(new_n221_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n261_), .B1(new_n264_), .B2(new_n219_), .ZN(new_n265_));
  OAI22_X1  g064(.A1(new_n254_), .A2(new_n263_), .B1(KEYINPUT12), .B2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n264_), .A2(new_n261_), .A3(new_n219_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G230gat), .A2(G233gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n202_), .B1(new_n266_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n241_), .A2(new_n253_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n219_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n263_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n219_), .B1(new_n236_), .B2(new_n240_), .ZN(new_n275_));
  AOI21_X1  g074(.A(KEYINPUT12), .B1(new_n275_), .B2(new_n262_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n269_), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n274_), .A2(KEYINPUT70), .A3(new_n277_), .A4(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n270_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n265_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n268_), .B1(new_n281_), .B2(new_n267_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G120gat), .B(G148gat), .ZN(new_n285_));
  INV_X1    g084(.A(G204gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT5), .ZN(new_n288_));
  INV_X1    g087(.A(G176gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n284_), .A2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n280_), .A2(new_n283_), .A3(new_n290_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n294_), .A2(KEYINPUT13), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(KEYINPUT13), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT71), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n295_), .A2(new_n296_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT71), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G190gat), .B(G218gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(G134gat), .ZN(new_n304_));
  XOR2_X1   g103(.A(new_n304_), .B(G162gat), .Z(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G29gat), .B(G36gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(G43gat), .ZN(new_n308_));
  INV_X1    g107(.A(G50gat), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(G43gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n307_), .B(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n312_), .A2(G50gat), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n310_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n264_), .A2(new_n314_), .A3(new_n219_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G232gat), .A2(G233gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT34), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n312_), .A2(G50gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n308_), .A2(new_n309_), .ZN(new_n319_));
  AND3_X1   g118(.A1(new_n318_), .A2(new_n319_), .A3(KEYINPUT15), .ZN(new_n320_));
  AOI21_X1  g119(.A(KEYINPUT15), .B1(new_n318_), .B2(new_n319_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  OAI221_X1 g121(.A(new_n315_), .B1(KEYINPUT35), .B2(new_n317_), .C1(new_n254_), .C2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT72), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n315_), .A2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n325_), .A2(KEYINPUT35), .A3(new_n317_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n323_), .B(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT74), .B(KEYINPUT36), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n306_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n330_));
  NAND2_X1  g129(.A1(new_n327_), .A2(new_n330_), .ZN(new_n331_));
  AND3_X1   g130(.A1(new_n325_), .A2(KEYINPUT35), .A3(new_n317_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n323_), .B(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n328_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n333_), .A2(new_n334_), .A3(new_n305_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n329_), .A2(new_n331_), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT37), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT37), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n329_), .A2(new_n335_), .A3(new_n338_), .A4(new_n331_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G15gat), .B(G22gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G1gat), .A2(G8gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT14), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G1gat), .B(G8gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G231gat), .A2(G233gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(new_n262_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT17), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT16), .B(G183gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(G211gat), .ZN(new_n353_));
  XOR2_X1   g152(.A(G127gat), .B(G155gat), .Z(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  NOR3_X1   g154(.A1(new_n350_), .A2(new_n351_), .A3(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(new_n356_), .B(KEYINPUT75), .Z(new_n357_));
  XNOR2_X1  g156(.A(new_n355_), .B(new_n351_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT76), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n350_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n340_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G127gat), .B(G134gat), .ZN(new_n363_));
  INV_X1    g162(.A(G113gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(G120gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT83), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT25), .B(G183gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT26), .B(G190gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(G169gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(new_n289_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G169gat), .A2(G176gat), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(KEYINPUT24), .A3(new_n374_), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n371_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G183gat), .A2(G190gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT23), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n376_), .B(new_n378_), .C1(KEYINPUT24), .C2(new_n373_), .ZN(new_n379_));
  OR3_X1    g178(.A1(new_n377_), .A2(KEYINPUT80), .A3(KEYINPUT23), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT80), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n380_), .B1(new_n378_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(G183gat), .ZN(new_n383_));
  INV_X1    g182(.A(G190gat), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n382_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT79), .ZN(new_n386_));
  OR3_X1    g185(.A1(new_n386_), .A2(new_n372_), .A3(KEYINPUT22), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT22), .B1(new_n386_), .B2(new_n372_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n387_), .A2(new_n289_), .A3(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n374_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n379_), .B1(new_n385_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT81), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n379_), .B(KEYINPUT81), .C1(new_n385_), .C2(new_n390_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  OR2_X1    g194(.A1(new_n395_), .A2(KEYINPUT30), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(KEYINPUT30), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n368_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G15gat), .B(G43gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT82), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G71gat), .B(G99gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G227gat), .A2(G233gat), .ZN(new_n403_));
  XOR2_X1   g202(.A(new_n402_), .B(new_n403_), .Z(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT31), .B1(new_n398_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NOR3_X1   g205(.A1(new_n398_), .A2(KEYINPUT31), .A3(new_n404_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n367_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n407_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n367_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n409_), .A2(new_n410_), .A3(new_n405_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n408_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n396_), .A2(new_n397_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n413_), .A2(KEYINPUT83), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n412_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n408_), .A2(new_n411_), .A3(new_n414_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(G141gat), .ZN(new_n420_));
  INV_X1    g219(.A(G148gat), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(new_n421_), .A3(KEYINPUT85), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT85), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n423_), .B1(G141gat), .B2(G148gat), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT3), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n422_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT86), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT84), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n429_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT2), .ZN(new_n431_));
  NAND3_X1  g230(.A1(KEYINPUT84), .A2(G141gat), .A3(G148gat), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n420_), .A2(new_n421_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT3), .ZN(new_n435_));
  NAND3_X1  g234(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n433_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT87), .B1(new_n428_), .B2(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(G155gat), .B(G162gat), .Z(new_n439_));
  XNOR2_X1  g238(.A(new_n426_), .B(KEYINPUT86), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT87), .ZN(new_n441_));
  INV_X1    g240(.A(new_n437_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n438_), .A2(new_n439_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT1), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n439_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n448_), .A2(new_n434_), .A3(new_n430_), .A4(new_n432_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n444_), .A2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(KEYINPUT90), .B1(new_n450_), .B2(KEYINPUT29), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G197gat), .A2(G204gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT91), .B(G197gat), .ZN(new_n453_));
  OAI211_X1 g252(.A(KEYINPUT21), .B(new_n452_), .C1(new_n453_), .C2(G204gat), .ZN(new_n454_));
  XOR2_X1   g253(.A(G211gat), .B(G218gat), .Z(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n286_), .A2(G197gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n457_), .B1(new_n453_), .B2(new_n286_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n454_), .B(new_n456_), .C1(new_n458_), .C2(KEYINPUT21), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(KEYINPUT21), .A3(new_n455_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n451_), .A2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G78gat), .B(G106gat), .ZN(new_n463_));
  XOR2_X1   g262(.A(new_n462_), .B(new_n463_), .Z(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(G233gat), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT88), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n467_), .A2(G228gat), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(G228gat), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n466_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT28), .B1(new_n450_), .B2(KEYINPUT29), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT89), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT28), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT29), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n444_), .A2(new_n475_), .A3(new_n476_), .A4(new_n449_), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n473_), .A2(new_n474_), .A3(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n474_), .B1(new_n473_), .B2(new_n477_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n472_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n473_), .A2(new_n477_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT89), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n473_), .A2(new_n474_), .A3(new_n477_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n482_), .A2(new_n471_), .A3(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G22gat), .B(G50gat), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  AND3_X1   g285(.A1(new_n480_), .A2(new_n484_), .A3(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n486_), .B1(new_n480_), .B2(new_n484_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n465_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NOR3_X1   g288(.A1(new_n478_), .A2(new_n479_), .A3(new_n472_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n471_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n485_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n480_), .A2(new_n484_), .A3(new_n486_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n492_), .A2(new_n464_), .A3(new_n493_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n489_), .A2(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n378_), .B1(G183gat), .B2(G190gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT22), .B(G169gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(new_n289_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n496_), .A2(new_n374_), .A3(new_n498_), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n499_), .A2(KEYINPUT94), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(KEYINPUT94), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n373_), .A2(KEYINPUT24), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT92), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n502_), .B1(new_n376_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n371_), .A2(new_n375_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n382_), .B1(KEYINPUT92), .B2(new_n505_), .ZN(new_n506_));
  AND3_X1   g305(.A1(new_n504_), .A2(new_n506_), .A3(KEYINPUT93), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT93), .B1(new_n504_), .B2(new_n506_), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n500_), .B(new_n501_), .C1(new_n507_), .C2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n461_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G226gat), .A2(G233gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT19), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n461_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n393_), .A2(new_n394_), .A3(new_n514_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n510_), .A2(KEYINPUT20), .A3(new_n513_), .A4(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT98), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT20), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n519_), .B1(new_n395_), .B2(new_n461_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n504_), .A2(new_n506_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n521_), .A2(new_n514_), .A3(new_n499_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n512_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n519_), .B1(new_n509_), .B2(new_n461_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n525_), .A2(KEYINPUT98), .A3(new_n513_), .A4(new_n515_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n518_), .A2(new_n524_), .A3(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT18), .B(G64gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(G92gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G8gat), .B(G36gat), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n529_), .B(new_n530_), .Z(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n527_), .A2(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n513_), .B1(new_n525_), .B2(new_n515_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n509_), .A2(new_n461_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n536_), .A2(new_n513_), .A3(new_n520_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n535_), .A2(new_n537_), .A3(new_n531_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n533_), .A2(KEYINPUT27), .A3(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT27), .ZN(new_n540_));
  INV_X1    g339(.A(new_n537_), .ZN(new_n541_));
  NOR3_X1   g340(.A1(new_n541_), .A2(new_n534_), .A3(new_n532_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n531_), .B1(new_n535_), .B2(new_n537_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n540_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n539_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT95), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n444_), .A2(new_n546_), .A3(new_n449_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n410_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n444_), .A2(new_n546_), .A3(new_n449_), .A4(new_n367_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n548_), .A2(KEYINPUT4), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT4), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n450_), .A2(new_n551_), .A3(new_n410_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G225gat), .A2(G233gat), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT0), .B(G57gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(G85gat), .ZN(new_n558_));
  XOR2_X1   g357(.A(G1gat), .B(G29gat), .Z(new_n559_));
  XOR2_X1   g358(.A(new_n558_), .B(new_n559_), .Z(new_n560_));
  AOI21_X1  g359(.A(new_n555_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n556_), .A2(new_n560_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n560_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n554_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n564_), .B1(new_n565_), .B2(new_n561_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n495_), .A2(KEYINPUT100), .A3(new_n545_), .A4(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT100), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n489_), .A2(new_n494_), .A3(new_n544_), .A4(new_n539_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n570_), .B1(new_n571_), .B2(new_n567_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n572_), .ZN(new_n573_));
  OR3_X1    g372(.A1(new_n565_), .A2(KEYINPUT33), .A3(new_n561_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n532_), .B1(new_n541_), .B2(new_n534_), .ZN(new_n575_));
  OAI211_X1 g374(.A(KEYINPUT33), .B(new_n564_), .C1(new_n565_), .C2(new_n561_), .ZN(new_n576_));
  AND4_X1   g375(.A1(new_n574_), .A2(new_n575_), .A3(new_n538_), .A4(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(KEYINPUT96), .B1(new_n553_), .B2(new_n555_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n548_), .A2(new_n555_), .A3(new_n549_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT96), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n550_), .A2(new_n580_), .A3(new_n554_), .A4(new_n552_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n578_), .A2(new_n579_), .A3(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT33), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n560_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT97), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n577_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n564_), .B1(new_n582_), .B2(KEYINPUT33), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n574_), .A2(new_n575_), .A3(new_n538_), .A4(new_n576_), .ZN(new_n588_));
  OAI21_X1  g387(.A(KEYINPUT97), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n586_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n531_), .A2(KEYINPUT32), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n535_), .A2(new_n537_), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n591_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n527_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n567_), .A2(new_n592_), .A3(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n595_), .A2(KEYINPUT99), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT99), .ZN(new_n597_));
  AOI22_X1  g396(.A1(new_n563_), .A2(new_n566_), .B1(new_n527_), .B2(new_n593_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n597_), .B1(new_n598_), .B2(new_n592_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n596_), .A2(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n495_), .B1(new_n590_), .B2(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n419_), .B1(new_n573_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n545_), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n603_), .A2(new_n495_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n418_), .A2(new_n568_), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n602_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n346_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n314_), .A2(new_n608_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n310_), .A2(new_n313_), .A3(new_n346_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G229gat), .A2(G233gat), .ZN(new_n612_));
  OAI21_X1  g411(.A(KEYINPUT77), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n346_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n610_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n614_), .A2(new_n612_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT77), .ZN(new_n617_));
  INV_X1    g416(.A(new_n612_), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n617_), .B(new_n618_), .C1(new_n609_), .C2(new_n610_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G113gat), .B(G141gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(new_n372_), .ZN(new_n621_));
  INV_X1    g420(.A(G197gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n613_), .A2(new_n616_), .A3(new_n619_), .A4(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT78), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n613_), .A2(new_n616_), .A3(new_n619_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n623_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n626_), .B(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(KEYINPUT101), .B1(new_n607_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT101), .ZN(new_n631_));
  INV_X1    g430(.A(new_n629_), .ZN(new_n632_));
  AOI211_X1 g431(.A(new_n631_), .B(new_n632_), .C1(new_n602_), .C2(new_n606_), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n302_), .B(new_n362_), .C1(new_n630_), .C2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT102), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n604_), .A2(new_n605_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n595_), .A2(KEYINPUT99), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n598_), .A2(new_n597_), .A3(new_n592_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n639_), .B1(new_n589_), .B2(new_n586_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n572_), .B(new_n569_), .C1(new_n640_), .C2(new_n495_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n636_), .B1(new_n641_), .B2(new_n419_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n631_), .B1(new_n642_), .B2(new_n632_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n607_), .A2(KEYINPUT101), .A3(new_n629_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT102), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n645_), .A2(new_n646_), .A3(new_n302_), .A4(new_n362_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n635_), .A2(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n568_), .A2(G1gat), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT38), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n302_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n653_), .A2(new_n632_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n361_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n336_), .B(KEYINPUT103), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT104), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n607_), .A2(new_n654_), .A3(new_n655_), .A4(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G1gat), .B1(new_n658_), .B2(new_n568_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n648_), .A2(KEYINPUT38), .A3(new_n649_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n652_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT105), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n652_), .A2(new_n660_), .A3(KEYINPUT105), .A4(new_n659_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1324gat));
  NOR2_X1   g464(.A1(new_n545_), .A2(G8gat), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n648_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT106), .ZN(new_n668_));
  OAI21_X1  g467(.A(G8gat), .B1(new_n658_), .B2(new_n545_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT39), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n667_), .A2(new_n668_), .A3(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n666_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n672_), .B1(new_n635_), .B2(new_n647_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT39), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n669_), .B(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(KEYINPUT106), .B1(new_n673_), .B2(new_n675_), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n671_), .A2(KEYINPUT40), .A3(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT40), .B1(new_n671_), .B2(new_n676_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1325gat));
  OAI21_X1  g478(.A(G15gat), .B1(new_n658_), .B2(new_n419_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT41), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n634_), .A2(G15gat), .A3(new_n419_), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1326gat));
  XOR2_X1   g482(.A(new_n495_), .B(KEYINPUT107), .Z(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G22gat), .B1(new_n658_), .B2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT42), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n685_), .A2(G22gat), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n687_), .B1(new_n634_), .B2(new_n688_), .ZN(G1327gat));
  AOI21_X1  g488(.A(new_n653_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n656_), .A2(new_n655_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(G29gat), .B1(new_n693_), .B2(new_n567_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n695_), .B1(new_n607_), .B2(new_n340_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n340_), .ZN(new_n697_));
  AOI211_X1 g496(.A(KEYINPUT43), .B(new_n697_), .C1(new_n602_), .C2(new_n606_), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n361_), .B(new_n654_), .C1(new_n696_), .C2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700_));
  OAI21_X1  g499(.A(KEYINPUT108), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n654_), .ZN(new_n702_));
  OAI21_X1  g501(.A(KEYINPUT43), .B1(new_n642_), .B2(new_n697_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n607_), .A2(new_n695_), .A3(new_n340_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n702_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT108), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n705_), .A2(new_n706_), .A3(KEYINPUT44), .A4(new_n361_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n568_), .B1(new_n701_), .B2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n699_), .A2(new_n700_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n709_), .A2(G29gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n694_), .B1(new_n708_), .B2(new_n710_), .ZN(G1328gat));
  INV_X1    g510(.A(G36gat), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n701_), .A2(new_n707_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n545_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n712_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n545_), .A2(G36gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n693_), .A2(KEYINPUT45), .A3(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT45), .ZN(new_n718_));
  INV_X1    g517(.A(new_n716_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n692_), .B2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n717_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT46), .ZN(new_n722_));
  OR3_X1    g521(.A1(new_n715_), .A2(new_n721_), .A3(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(new_n715_), .B2(new_n721_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1329gat));
  NAND4_X1  g524(.A1(new_n713_), .A2(G43gat), .A3(new_n418_), .A4(new_n709_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n311_), .B1(new_n692_), .B2(new_n419_), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n726_), .A2(new_n727_), .A3(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n727_), .B1(new_n726_), .B2(new_n728_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1330gat));
  NAND4_X1  g530(.A1(new_n713_), .A2(G50gat), .A3(new_n495_), .A4(new_n709_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n309_), .B1(new_n692_), .B2(new_n685_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n732_), .A2(KEYINPUT110), .A3(new_n733_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(G1331gat));
  NAND2_X1  g537(.A1(new_n653_), .A2(new_n362_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT111), .Z(new_n740_));
  NOR3_X1   g539(.A1(new_n740_), .A2(new_n642_), .A3(new_n629_), .ZN(new_n741_));
  AOI21_X1  g540(.A(G57gat), .B1(new_n741_), .B2(new_n567_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n653_), .A2(new_n632_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n657_), .ZN(new_n744_));
  NOR4_X1   g543(.A1(new_n642_), .A2(new_n743_), .A3(new_n361_), .A4(new_n744_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n745_), .A2(new_n567_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n742_), .B1(G57gat), .B2(new_n746_), .ZN(G1332gat));
  INV_X1    g546(.A(G64gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n745_), .B2(new_n603_), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT48), .Z(new_n750_));
  NAND3_X1  g549(.A1(new_n741_), .A2(new_n748_), .A3(new_n603_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1333gat));
  INV_X1    g551(.A(G71gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n745_), .B2(new_n418_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT49), .Z(new_n755_));
  NAND3_X1  g554(.A1(new_n741_), .A2(new_n753_), .A3(new_n418_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT112), .ZN(G1334gat));
  INV_X1    g557(.A(G78gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n745_), .B2(new_n684_), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT50), .Z(new_n761_));
  NAND3_X1  g560(.A1(new_n741_), .A2(new_n759_), .A3(new_n684_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(G1335gat));
  NAND3_X1  g562(.A1(new_n653_), .A2(new_n361_), .A3(new_n632_), .ZN(new_n764_));
  NOR3_X1   g563(.A1(new_n642_), .A2(new_n764_), .A3(new_n656_), .ZN(new_n765_));
  AOI21_X1  g564(.A(G85gat), .B1(new_n765_), .B2(new_n567_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n764_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(new_n567_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n766_), .B1(new_n769_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g569(.A(G92gat), .B1(new_n765_), .B2(new_n603_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n545_), .A2(new_n204_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n767_), .B2(new_n772_), .ZN(G1337gat));
  AOI21_X1  g572(.A(new_n228_), .B1(new_n767_), .B2(new_n418_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n418_), .A2(new_n216_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n765_), .B2(new_n775_), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n776_), .B(KEYINPUT51), .Z(G1338gat));
  AOI21_X1  g576(.A(new_n217_), .B1(new_n767_), .B2(new_n495_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779_));
  OAI21_X1  g578(.A(KEYINPUT114), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n778_), .A2(KEYINPUT113), .A3(new_n779_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT113), .ZN(new_n782_));
  INV_X1    g581(.A(new_n764_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n495_), .B(new_n783_), .C1(new_n696_), .C2(new_n698_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(G106gat), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n782_), .B1(new_n785_), .B2(KEYINPUT52), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n785_), .A2(new_n787_), .A3(KEYINPUT52), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n780_), .A2(new_n781_), .A3(new_n786_), .A4(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n765_), .A2(new_n217_), .A3(new_n495_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT53), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n789_), .A2(new_n793_), .A3(new_n790_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(G1339gat));
  INV_X1    g594(.A(KEYINPUT122), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n604_), .A2(new_n419_), .A3(new_n568_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT57), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT118), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n276_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT70), .B1(new_n802_), .B2(new_n278_), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n266_), .A2(new_n202_), .A3(new_n269_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n801_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n268_), .B1(new_n802_), .B2(new_n267_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n266_), .A2(new_n801_), .A3(new_n269_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n805_), .A2(new_n806_), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT55), .B1(new_n270_), .B2(new_n279_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n802_), .A2(KEYINPUT55), .A3(new_n278_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n268_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n267_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n813_), .B1(new_n266_), .B2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n812_), .A2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(KEYINPUT117), .B1(new_n811_), .B2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n810_), .A2(new_n817_), .A3(new_n291_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT56), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n810_), .A2(new_n817_), .A3(KEYINPUT56), .A4(new_n291_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n629_), .A2(new_n293_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n800_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n825_));
  AOI211_X1 g624(.A(KEYINPUT118), .B(new_n823_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n614_), .A2(new_n618_), .A3(new_n615_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n618_), .B2(new_n611_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n625_), .B1(new_n624_), .B2(new_n828_), .ZN(new_n829_));
  XOR2_X1   g628(.A(new_n829_), .B(KEYINPUT119), .Z(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n294_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n825_), .A2(new_n826_), .A3(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n656_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n799_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n822_), .A2(new_n824_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT118), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n822_), .A2(new_n800_), .A3(new_n824_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(new_n831_), .A3(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(KEYINPUT57), .A3(new_n656_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT58), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n822_), .A2(KEYINPUT120), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n830_), .B(new_n293_), .C1(new_n821_), .C2(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n841_), .B1(new_n842_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n844_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n846_), .B(KEYINPUT58), .C1(KEYINPUT120), .C2(new_n822_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n845_), .A2(new_n340_), .A3(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n835_), .A2(new_n840_), .A3(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(new_n361_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n337_), .A2(new_n655_), .A3(new_n632_), .A4(new_n339_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n297_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(KEYINPUT115), .A3(new_n853_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n362_), .A2(new_n853_), .A3(new_n632_), .A4(new_n299_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT116), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n859_));
  OAI211_X1 g658(.A(KEYINPUT116), .B(KEYINPUT54), .C1(new_n297_), .C2(new_n851_), .ZN(new_n860_));
  AND4_X1   g659(.A1(new_n854_), .A2(new_n857_), .A3(new_n859_), .A4(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n798_), .B1(new_n850_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT59), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n796_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n861_), .B1(new_n849_), .B2(new_n361_), .ZN(new_n866_));
  NOR4_X1   g665(.A1(new_n866_), .A2(KEYINPUT122), .A3(KEYINPUT59), .A4(new_n798_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n865_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n870_));
  OAI211_X1 g669(.A(KEYINPUT121), .B(KEYINPUT59), .C1(new_n866_), .C2(new_n798_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n868_), .A2(new_n872_), .A3(G113gat), .A4(new_n629_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n863_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n364_), .B1(new_n874_), .B2(new_n632_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n873_), .A2(new_n875_), .ZN(G1340gat));
  OAI21_X1  g675(.A(new_n366_), .B1(new_n302_), .B2(KEYINPUT60), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n863_), .B(new_n877_), .C1(KEYINPUT60), .C2(new_n366_), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n868_), .A2(new_n653_), .A3(new_n872_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n879_), .B2(new_n366_), .ZN(G1341gat));
  NAND2_X1  g679(.A1(new_n655_), .A2(G127gat), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n868_), .A2(new_n872_), .A3(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(G127gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(new_n874_), .B2(new_n361_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT123), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n883_), .A2(KEYINPUT123), .A3(new_n885_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(G1342gat));
  AOI21_X1  g689(.A(G134gat), .B1(new_n863_), .B2(new_n744_), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n868_), .A2(new_n340_), .A3(new_n872_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(G134gat), .ZN(G1343gat));
  NAND2_X1  g692(.A1(new_n850_), .A2(new_n862_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n571_), .A2(new_n568_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n894_), .A2(new_n419_), .A3(new_n895_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(KEYINPUT124), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n629_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n653_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(KEYINPUT125), .B(G148gat), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n900_), .B(new_n902_), .ZN(G1345gat));
  NAND2_X1  g702(.A1(new_n897_), .A2(new_n655_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(KEYINPUT61), .B(G155gat), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n904_), .B(new_n905_), .ZN(G1346gat));
  AOI21_X1  g705(.A(G162gat), .B1(new_n897_), .B2(new_n744_), .ZN(new_n907_));
  AND2_X1   g706(.A1(new_n897_), .A2(new_n340_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(G162gat), .B2(new_n908_), .ZN(G1347gat));
  INV_X1    g708(.A(KEYINPUT126), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n605_), .A2(new_n545_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n866_), .A2(new_n684_), .A3(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n629_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n910_), .B1(new_n915_), .B2(new_n372_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n914_), .A2(KEYINPUT126), .A3(G169gat), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n916_), .A2(KEYINPUT62), .A3(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n915_), .A2(new_n497_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n920_));
  OAI211_X1 g719(.A(new_n910_), .B(new_n920_), .C1(new_n915_), .C2(new_n372_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n918_), .A2(new_n919_), .A3(new_n921_), .ZN(G1348gat));
  AOI21_X1  g721(.A(G176gat), .B1(new_n913_), .B2(new_n653_), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n866_), .A2(new_n495_), .A3(new_n912_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n302_), .A2(new_n289_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n923_), .B1(new_n924_), .B2(new_n925_), .ZN(G1349gat));
  AOI21_X1  g725(.A(G183gat), .B1(new_n924_), .B2(new_n655_), .ZN(new_n927_));
  OR2_X1    g726(.A1(new_n361_), .A2(new_n369_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n927_), .B1(new_n913_), .B2(new_n929_), .ZN(G1350gat));
  NAND3_X1  g729(.A1(new_n913_), .A2(new_n744_), .A3(new_n370_), .ZN(new_n931_));
  AND2_X1   g730(.A1(new_n913_), .A2(new_n340_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n932_), .B2(new_n384_), .ZN(G1351gat));
  NAND2_X1  g732(.A1(new_n894_), .A2(new_n419_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n603_), .A2(new_n568_), .A3(new_n495_), .ZN(new_n935_));
  NOR3_X1   g734(.A1(new_n934_), .A2(new_n632_), .A3(new_n935_), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n936_), .A2(KEYINPUT127), .A3(new_n622_), .ZN(new_n937_));
  XOR2_X1   g736(.A(KEYINPUT127), .B(G197gat), .Z(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n936_), .B2(new_n938_), .ZN(G1352gat));
  NOR2_X1   g738(.A1(new_n934_), .A2(new_n935_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(new_n653_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(G204gat), .ZN(G1353gat));
  NOR3_X1   g741(.A1(new_n934_), .A2(new_n361_), .A3(new_n935_), .ZN(new_n943_));
  NOR3_X1   g742(.A1(new_n943_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n944_));
  XOR2_X1   g743(.A(KEYINPUT63), .B(G211gat), .Z(new_n945_));
  AOI21_X1  g744(.A(new_n944_), .B1(new_n943_), .B2(new_n945_), .ZN(G1354gat));
  NOR3_X1   g745(.A1(new_n934_), .A2(new_n657_), .A3(new_n935_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n940_), .A2(new_n340_), .ZN(new_n948_));
  MUX2_X1   g747(.A(new_n947_), .B(new_n948_), .S(G218gat), .Z(G1355gat));
endmodule


