//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 1 0 0 0 1 1 0 1 1 0 0 0 1 0 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n777_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n910_, new_n912_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n946_, new_n947_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n959_, new_n960_, new_n962_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n969_, new_n970_,
    new_n971_;
  NOR2_X1   g000(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G169gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT23), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND3_X1  g005(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n207_));
  OAI211_X1 g006(.A(new_n206_), .B(new_n207_), .C1(G183gat), .C2(G190gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n203_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT26), .B(G190gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT25), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G183gat), .ZN(new_n212_));
  OR2_X1    g011(.A1(new_n211_), .A2(G183gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n210_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  AND2_X1   g013(.A1(new_n206_), .A2(new_n207_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT24), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n214_), .A2(new_n215_), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT24), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n221_), .A2(KEYINPUT91), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT91), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n223_), .B1(new_n220_), .B2(KEYINPUT24), .ZN(new_n224_));
  NOR3_X1   g023(.A1(new_n222_), .A2(new_n224_), .A3(new_n216_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n209_), .B1(new_n219_), .B2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G197gat), .B(G204gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT88), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G211gat), .B(G218gat), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  OR2_X1    g030(.A1(G197gat), .A2(G204gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G197gat), .A2(G204gat), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(KEYINPUT88), .A3(new_n233_), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n229_), .A2(new_n231_), .A3(KEYINPUT21), .A4(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n227_), .A2(KEYINPUT21), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT21), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n232_), .A2(new_n237_), .A3(new_n233_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n231_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n235_), .B1(new_n239_), .B2(KEYINPUT87), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT87), .ZN(new_n241_));
  AOI211_X1 g040(.A(new_n241_), .B(new_n231_), .C1(new_n236_), .C2(new_n238_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n226_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT77), .B(G183gat), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n245_), .A2(KEYINPUT78), .A3(KEYINPUT25), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n210_), .A2(new_n212_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT78), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n248_), .B1(new_n244_), .B2(new_n211_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n246_), .A2(new_n247_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n215_), .A2(new_n218_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n221_), .A2(new_n216_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n250_), .A2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n215_), .B1(G190gat), .B2(new_n244_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(new_n203_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n238_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n237_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n230_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(new_n241_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n239_), .A2(KEYINPUT87), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n261_), .A2(new_n262_), .A3(new_n235_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n243_), .B(KEYINPUT20), .C1(new_n257_), .C2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G226gat), .A2(G233gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT19), .ZN(new_n266_));
  OR2_X1    g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n257_), .A2(new_n263_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n240_), .A2(new_n242_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n226_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n268_), .A2(new_n271_), .A3(KEYINPUT20), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n266_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n267_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G64gat), .B(G92gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n275_), .B(KEYINPUT94), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT95), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n276_), .B(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G8gat), .B(G36gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n274_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT27), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n264_), .A2(new_n266_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n266_), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n268_), .A2(new_n271_), .A3(KEYINPUT20), .A4(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n285_), .A2(KEYINPUT92), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT92), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n264_), .A2(new_n289_), .A3(new_n266_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n282_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT103), .B1(new_n284_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n291_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT103), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n293_), .A2(new_n294_), .A3(KEYINPUT27), .A4(new_n283_), .ZN(new_n295_));
  AND3_X1   g094(.A1(new_n288_), .A2(new_n282_), .A3(new_n290_), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n296_), .A2(new_n291_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT27), .ZN(new_n298_));
  AOI22_X1  g097(.A1(new_n292_), .A2(new_n295_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G155gat), .B(G162gat), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n300_), .A2(KEYINPUT1), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G141gat), .A2(G148gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT83), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT83), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n304_), .A2(G141gat), .A3(G148gat), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(G141gat), .A2(G148gat), .ZN(new_n307_));
  AND2_X1   g106(.A1(G155gat), .A2(G162gat), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n307_), .B1(new_n308_), .B2(KEYINPUT1), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n301_), .A2(new_n306_), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT3), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n307_), .A2(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n312_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT2), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n303_), .A2(new_n305_), .A3(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n300_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n310_), .B1(new_n318_), .B2(KEYINPUT84), .ZN(new_n319_));
  INV_X1    g118(.A(new_n300_), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n303_), .A2(new_n305_), .A3(new_n316_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n312_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n320_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT84), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n319_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT29), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT28), .B(G22gat), .ZN(new_n328_));
  INV_X1    g127(.A(G50gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n326_), .A2(new_n327_), .A3(new_n331_), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n306_), .A2(new_n309_), .ZN(new_n333_));
  AOI22_X1  g132(.A1(new_n323_), .A2(new_n324_), .B1(new_n333_), .B2(new_n301_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n318_), .A2(KEYINPUT84), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n334_), .A2(new_n327_), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n330_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n332_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT85), .B(KEYINPUT86), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G228gat), .A2(G233gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n327_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n343_), .B1(new_n344_), .B2(new_n269_), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n263_), .B(new_n342_), .C1(new_n326_), .C2(new_n327_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G78gat), .B(G106gat), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n345_), .A2(new_n346_), .A3(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n332_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n341_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  AOI211_X1 g150(.A(KEYINPUT90), .B(new_n348_), .C1(new_n345_), .C2(new_n346_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n348_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT90), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n341_), .A2(new_n350_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n349_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n357_), .B1(new_n358_), .B2(new_n354_), .ZN(new_n359_));
  AOI22_X1  g158(.A1(new_n353_), .A2(new_n356_), .B1(new_n359_), .B2(KEYINPUT89), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n359_), .A2(KEYINPUT89), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G127gat), .B(G134gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G113gat), .B(G120gat), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n365_), .A2(KEYINPUT81), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n363_), .B(new_n364_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n366_), .B1(new_n367_), .B2(KEYINPUT81), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n368_), .B1(new_n319_), .B2(new_n325_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n334_), .A2(new_n367_), .A3(new_n335_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n369_), .A2(new_n370_), .A3(KEYINPUT4), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT96), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n369_), .A2(new_n370_), .A3(KEYINPUT96), .A4(KEYINPUT4), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT98), .B(KEYINPUT4), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n368_), .B(new_n376_), .C1(new_n319_), .C2(new_n325_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G225gat), .A2(G233gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT97), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n375_), .A2(new_n380_), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n369_), .A2(new_n370_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n382_), .A2(KEYINPUT100), .A3(new_n378_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n369_), .A2(new_n370_), .A3(new_n378_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT100), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n383_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n381_), .A2(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(G1gat), .B(G29gat), .Z(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT99), .B(G85gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT0), .B(G57gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n388_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n381_), .A2(new_n393_), .A3(new_n387_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G227gat), .A2(G233gat), .ZN(new_n399_));
  XOR2_X1   g198(.A(new_n399_), .B(KEYINPUT80), .Z(new_n400_));
  XOR2_X1   g199(.A(new_n400_), .B(KEYINPUT30), .Z(new_n401_));
  XNOR2_X1  g200(.A(new_n257_), .B(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G15gat), .B(G43gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT79), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(G71gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n402_), .B(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n368_), .B(KEYINPUT31), .ZN(new_n407_));
  XOR2_X1   g206(.A(new_n407_), .B(G99gat), .Z(new_n408_));
  OR2_X1    g207(.A1(new_n406_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n406_), .A2(new_n408_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n299_), .A2(new_n362_), .A3(new_n398_), .A4(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n281_), .A2(KEYINPUT32), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n413_), .B1(new_n273_), .B2(new_n267_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n288_), .A2(new_n290_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n414_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n397_), .A2(new_n416_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n296_), .A2(new_n291_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT33), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n396_), .A2(new_n419_), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n377_), .A2(new_n378_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n375_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT102), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT102), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n375_), .A2(new_n424_), .A3(new_n421_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n393_), .B1(new_n382_), .B2(new_n379_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n423_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n418_), .A2(new_n420_), .A3(new_n427_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n381_), .A2(new_n387_), .A3(KEYINPUT33), .A4(new_n393_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT101), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n375_), .A2(new_n380_), .B1(new_n383_), .B2(new_n386_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT101), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n431_), .A2(new_n432_), .A3(KEYINPUT33), .A4(new_n393_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n430_), .A2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n417_), .B1(new_n428_), .B2(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n397_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n435_), .A2(new_n362_), .B1(new_n299_), .B2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n411_), .B(KEYINPUT82), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n412_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G1gat), .B(G8gat), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT75), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(G15gat), .ZN(new_n444_));
  INV_X1    g243(.A(G22gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G15gat), .A2(G22gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G1gat), .A2(G8gat), .ZN(new_n448_));
  AOI22_X1  g247(.A1(new_n446_), .A2(new_n447_), .B1(KEYINPUT14), .B2(new_n448_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n443_), .A2(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n443_), .A2(new_n449_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G43gat), .B(G50gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G29gat), .B(G36gat), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n454_), .A2(KEYINPUT73), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(KEYINPUT73), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n453_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n455_), .A2(new_n456_), .A3(new_n453_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n452_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n443_), .B(new_n449_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n459_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n463_), .A2(new_n457_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n461_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G229gat), .A2(G233gat), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT15), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n470_), .B1(new_n463_), .B2(new_n457_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n458_), .A2(KEYINPUT15), .A3(new_n459_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(new_n472_), .A3(new_n462_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(new_n461_), .A3(new_n467_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n469_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G113gat), .B(G141gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G169gat), .B(G197gat), .ZN(new_n478_));
  XOR2_X1   g277(.A(new_n477_), .B(new_n478_), .Z(new_n479_));
  NAND2_X1  g278(.A1(new_n476_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n479_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n475_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n440_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT11), .ZN(new_n485_));
  INV_X1    g284(.A(G57gat), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n486_), .A2(G64gat), .ZN(new_n487_));
  INV_X1    g286(.A(G64gat), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n488_), .A2(G57gat), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n485_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(G57gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n486_), .A2(G64gat), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(new_n492_), .A3(KEYINPUT11), .ZN(new_n493_));
  INV_X1    g292(.A(G78gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(G71gat), .ZN(new_n495_));
  INV_X1    g294(.A(G71gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(G78gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n490_), .A2(new_n493_), .A3(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G57gat), .B(G64gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G71gat), .B(G78gat), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(new_n501_), .A3(KEYINPUT11), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n499_), .A2(KEYINPUT12), .A3(new_n502_), .ZN(new_n503_));
  OR2_X1    g302(.A1(G85gat), .A2(G92gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G85gat), .A2(G92gat), .ZN(new_n505_));
  AOI21_X1  g304(.A(KEYINPUT8), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  OR2_X1    g305(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT65), .ZN(new_n508_));
  INV_X1    g307(.A(G106gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(KEYINPUT65), .A2(G106gat), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n507_), .A2(new_n510_), .A3(new_n511_), .A4(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(G92gat), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n514_), .A2(KEYINPUT9), .ZN(new_n515_));
  AND2_X1   g314(.A1(KEYINPUT66), .A2(G85gat), .ZN(new_n516_));
  NOR2_X1   g315(.A1(KEYINPUT66), .A2(G85gat), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n515_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n504_), .A2(KEYINPUT9), .A3(new_n505_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n513_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  OR3_X1    g319(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT8), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n521_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n520_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT6), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n526_), .B1(G99gat), .B2(G106gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G99gat), .A2(G106gat), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n528_), .A2(KEYINPUT6), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT67), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(KEYINPUT6), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n526_), .A2(G99gat), .A3(G106gat), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT67), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n530_), .A2(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n506_), .B1(new_n525_), .B2(new_n535_), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT68), .B1(new_n527_), .B2(new_n529_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT68), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n531_), .A2(new_n532_), .A3(new_n538_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n537_), .A2(new_n539_), .A3(new_n521_), .A4(new_n523_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n504_), .A2(KEYINPUT8), .A3(new_n505_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n503_), .B1(new_n536_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n525_), .A2(new_n535_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n506_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(new_n542_), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT69), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n493_), .A2(new_n498_), .ZN(new_n548_));
  AOI21_X1  g347(.A(KEYINPUT11), .B1(new_n491_), .B2(new_n492_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n547_), .B(new_n502_), .C1(new_n548_), .C2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n547_), .B1(new_n499_), .B2(new_n502_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n546_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT12), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n543_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G230gat), .A2(G233gat), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n557_), .B(KEYINPUT64), .Z(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n546_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n553_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n559_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n556_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT70), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n546_), .A2(new_n553_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(new_n554_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(new_n559_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT70), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n556_), .A2(new_n569_), .A3(new_n562_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n564_), .A2(new_n568_), .A3(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G120gat), .B(G148gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT5), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G176gat), .B(G204gat), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n573_), .B(new_n574_), .Z(new_n575_));
  NAND2_X1  g374(.A1(new_n571_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n575_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n564_), .A2(new_n568_), .A3(new_n570_), .A4(new_n577_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n576_), .A2(KEYINPUT13), .A3(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(KEYINPUT13), .B1(new_n576_), .B2(new_n578_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT71), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT71), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n583_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n584_));
  AOI21_X1  g383(.A(KEYINPUT72), .B1(new_n582_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n582_), .A2(new_n584_), .A3(KEYINPUT72), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n452_), .B(KEYINPUT76), .ZN(new_n589_));
  AND2_X1   g388(.A1(G231gat), .A2(G233gat), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n590_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n499_), .A2(new_n502_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(G127gat), .B(G155gat), .Z(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT16), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G183gat), .B(G211gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT17), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n591_), .A2(new_n502_), .A3(new_n499_), .A4(new_n592_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n595_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n593_), .A2(new_n553_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n591_), .A2(new_n592_), .A3(new_n561_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n599_), .B(KEYINPUT17), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n604_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n603_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n471_), .A2(new_n546_), .A3(new_n472_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G232gat), .A2(G233gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT34), .ZN(new_n612_));
  OAI22_X1  g411(.A1(new_n546_), .A2(new_n464_), .B1(KEYINPUT35), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n612_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT35), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  OR3_X1    g415(.A1(new_n610_), .A2(new_n613_), .A3(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n616_), .B1(new_n610_), .B2(new_n613_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G190gat), .B(G218gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G134gat), .B(G162gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT36), .Z(new_n623_));
  NAND2_X1  g422(.A1(new_n619_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n622_), .A2(KEYINPUT36), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n617_), .A2(new_n618_), .A3(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n624_), .A2(KEYINPUT37), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT74), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n624_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n619_), .A2(KEYINPUT74), .A3(new_n623_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n630_), .A2(new_n626_), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT37), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n628_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n484_), .A2(new_n588_), .A3(new_n609_), .A4(new_n634_), .ZN(new_n635_));
  OR3_X1    g434(.A1(new_n635_), .A2(G1gat), .A3(new_n398_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT38), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n440_), .A2(new_n632_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n582_), .A2(new_n584_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(new_n483_), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n639_), .A2(new_n608_), .A3(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G1gat), .B1(new_n644_), .B2(new_n398_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n636_), .A2(new_n637_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n638_), .A2(new_n645_), .A3(new_n646_), .ZN(G1324gat));
  XNOR2_X1  g446(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n642_), .A2(new_n608_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n299_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n649_), .A2(new_n650_), .A3(new_n440_), .A4(new_n632_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(G8gat), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT39), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n651_), .A2(KEYINPUT39), .A3(G8gat), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT104), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n299_), .A2(G8gat), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n657_), .B1(new_n635_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n588_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n634_), .A2(new_n609_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n663_), .A2(KEYINPUT104), .A3(new_n484_), .A4(new_n658_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n660_), .A2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n648_), .B1(new_n656_), .B2(new_n665_), .ZN(new_n666_));
  AND4_X1   g465(.A1(new_n665_), .A2(new_n655_), .A3(new_n654_), .A4(new_n648_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1325gat));
  INV_X1    g467(.A(new_n635_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n444_), .A3(new_n439_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n643_), .A2(new_n439_), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n671_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT41), .B1(new_n671_), .B2(G15gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n670_), .B1(new_n672_), .B2(new_n673_), .ZN(G1326gat));
  INV_X1    g473(.A(new_n362_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n669_), .A2(new_n445_), .A3(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n643_), .A2(new_n675_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n677_), .A2(G22gat), .A3(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n678_), .B1(new_n677_), .B2(G22gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n676_), .B1(new_n679_), .B2(new_n680_), .ZN(G1327gat));
  NAND3_X1  g480(.A1(new_n641_), .A2(new_n483_), .A3(new_n608_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT43), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n630_), .A2(new_n626_), .A3(new_n631_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n627_), .B1(new_n685_), .B2(KEYINPUT37), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n440_), .A2(new_n684_), .A3(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n684_), .B1(new_n440_), .B2(new_n686_), .ZN(new_n688_));
  OAI211_X1 g487(.A(KEYINPUT44), .B(new_n683_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n440_), .A2(new_n686_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT43), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n440_), .A2(new_n684_), .A3(new_n686_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n682_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  XOR2_X1   g492(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n694_));
  OAI21_X1  g493(.A(new_n689_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n397_), .A2(G29gat), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(G29gat), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n685_), .A2(new_n608_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n640_), .A2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n484_), .A2(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n698_), .B1(new_n701_), .B2(new_n398_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n697_), .A2(new_n702_), .ZN(G1328gat));
  OAI211_X1 g502(.A(new_n689_), .B(new_n650_), .C1(new_n693_), .C2(new_n694_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(G36gat), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n299_), .A2(G36gat), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n484_), .A2(new_n700_), .A3(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT45), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n705_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT46), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n705_), .A2(KEYINPUT46), .A3(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1329gat));
  XOR2_X1   g512(.A(KEYINPUT108), .B(G43gat), .Z(new_n714_));
  OAI21_X1  g513(.A(new_n714_), .B1(new_n701_), .B2(new_n438_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n411_), .A2(G43gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n715_), .B1(new_n695_), .B2(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI211_X1 g517(.A(new_n689_), .B(new_n675_), .C1(new_n693_), .C2(new_n694_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT109), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n719_), .A2(new_n720_), .A3(G50gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n719_), .B2(G50gat), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n362_), .A2(G50gat), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT110), .ZN(new_n724_));
  OAI22_X1  g523(.A1(new_n721_), .A2(new_n722_), .B1(new_n701_), .B2(new_n724_), .ZN(G1331gat));
  INV_X1    g524(.A(new_n483_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n440_), .A2(new_n726_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n727_), .A2(new_n641_), .A3(new_n662_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n728_), .A2(new_n486_), .A3(new_n397_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n608_), .A2(new_n483_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n586_), .A2(new_n587_), .A3(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(KEYINPUT111), .B1(new_n639_), .B2(new_n731_), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n582_), .A2(new_n584_), .A3(KEYINPUT72), .ZN(new_n733_));
  INV_X1    g532(.A(new_n730_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n733_), .A2(new_n585_), .A3(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT111), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n735_), .A2(new_n736_), .A3(new_n440_), .A4(new_n632_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n732_), .A2(new_n737_), .A3(new_n397_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n729_), .B1(new_n738_), .B2(new_n486_), .ZN(G1332gat));
  NAND3_X1  g538(.A1(new_n728_), .A2(new_n488_), .A3(new_n650_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n732_), .A2(new_n737_), .A3(new_n650_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT48), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n741_), .A2(new_n742_), .A3(G64gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n741_), .B2(G64gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(KEYINPUT112), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT112), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n747_), .B(new_n740_), .C1(new_n743_), .C2(new_n744_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(G1333gat));
  NAND3_X1  g548(.A1(new_n728_), .A2(new_n496_), .A3(new_n439_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n732_), .A2(new_n737_), .A3(new_n439_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT49), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n751_), .A2(new_n752_), .A3(G71gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n751_), .B2(G71gat), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n750_), .B1(new_n753_), .B2(new_n754_), .ZN(G1334gat));
  NAND3_X1  g554(.A1(new_n728_), .A2(new_n494_), .A3(new_n675_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n732_), .A2(new_n737_), .A3(new_n675_), .ZN(new_n757_));
  XOR2_X1   g556(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n758_));
  AND3_X1   g557(.A1(new_n757_), .A2(G78gat), .A3(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n757_), .B2(G78gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n756_), .B1(new_n759_), .B2(new_n760_), .ZN(G1335gat));
  NOR3_X1   g560(.A1(new_n727_), .A2(new_n588_), .A3(new_n699_), .ZN(new_n762_));
  AOI21_X1  g561(.A(G85gat), .B1(new_n762_), .B2(new_n397_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n691_), .A2(new_n692_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n640_), .A2(new_n726_), .A3(new_n608_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT114), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT115), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n764_), .A2(KEYINPUT115), .A3(new_n766_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n516_), .A2(new_n517_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n398_), .A2(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n763_), .B1(new_n771_), .B2(new_n773_), .ZN(G1336gat));
  NAND3_X1  g573(.A1(new_n769_), .A2(new_n650_), .A3(new_n770_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(G92gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n762_), .A2(new_n514_), .A3(new_n650_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(G1337gat));
  OAI21_X1  g577(.A(G99gat), .B1(new_n767_), .B2(new_n438_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n762_), .A2(new_n411_), .A3(new_n507_), .A4(new_n511_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g581(.A1(new_n762_), .A2(new_n675_), .A3(new_n510_), .A4(new_n512_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n766_), .B(new_n675_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n784_), .A2(new_n785_), .A3(G106gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n784_), .B2(G106gat), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n783_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT53), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n790_), .B(new_n783_), .C1(new_n786_), .C2(new_n787_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(G1339gat));
  NAND3_X1  g591(.A1(new_n730_), .A2(new_n634_), .A3(new_n581_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(KEYINPUT116), .A2(KEYINPUT54), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n730_), .A2(new_n634_), .A3(new_n581_), .A4(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n576_), .A2(new_n578_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n479_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n473_), .A2(new_n461_), .A3(new_n468_), .ZN(new_n803_));
  AOI22_X1  g602(.A1(new_n476_), .A2(new_n479_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n801_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n483_), .A2(new_n578_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT117), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n556_), .A2(KEYINPUT55), .A3(new_n562_), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT12), .B1(new_n546_), .B2(new_n553_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n810_), .A2(new_n565_), .A3(new_n543_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n809_), .B1(new_n811_), .B2(new_n558_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n558_), .B1(new_n546_), .B2(new_n553_), .ZN(new_n813_));
  NOR4_X1   g612(.A1(new_n813_), .A2(new_n810_), .A3(KEYINPUT70), .A4(new_n543_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n569_), .B1(new_n556_), .B2(new_n562_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n812_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n808_), .B1(new_n818_), .B2(new_n577_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT56), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n807_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n564_), .A2(new_n817_), .A3(new_n570_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n813_), .A2(new_n810_), .A3(new_n543_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n556_), .A2(new_n566_), .ZN(new_n824_));
  AOI22_X1  g623(.A1(new_n823_), .A2(KEYINPUT55), .B1(new_n824_), .B2(new_n559_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n822_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n575_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n827_), .A2(new_n808_), .A3(KEYINPUT56), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n806_), .B1(new_n821_), .B2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n800_), .B1(new_n829_), .B2(new_n685_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n577_), .B1(new_n822_), .B2(new_n825_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n820_), .B1(new_n831_), .B2(KEYINPUT117), .ZN(new_n832_));
  INV_X1    g631(.A(new_n807_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n828_), .A2(new_n832_), .A3(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n805_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n835_), .A2(KEYINPUT57), .A3(new_n632_), .ZN(new_n836_));
  OAI21_X1  g635(.A(KEYINPUT56), .B1(new_n818_), .B2(new_n577_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n831_), .A2(new_n820_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n804_), .A2(new_n578_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n837_), .A2(new_n838_), .A3(KEYINPUT58), .A4(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT118), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n804_), .A2(new_n578_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n827_), .B2(KEYINPUT56), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT118), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n843_), .A2(new_n844_), .A3(KEYINPUT58), .A4(new_n838_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n837_), .A2(new_n838_), .A3(new_n839_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT58), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n841_), .A2(new_n845_), .A3(new_n848_), .A4(new_n686_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n830_), .A2(new_n836_), .A3(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n799_), .B1(new_n850_), .B2(new_n608_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n650_), .A2(new_n675_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n397_), .A2(new_n411_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT59), .B1(new_n851_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(G113gat), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n726_), .A2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n685_), .B1(new_n834_), .B2(new_n805_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n849_), .B1(KEYINPUT57), .B2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(KEYINPUT121), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n830_), .A2(new_n861_), .A3(new_n849_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n860_), .A2(new_n836_), .A3(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n799_), .B1(new_n863_), .B2(new_n608_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n854_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n855_), .B(new_n857_), .C1(new_n864_), .C2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT119), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n851_), .A2(new_n726_), .A3(new_n854_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n870_), .B2(G113gat), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n850_), .A2(new_n608_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n798_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n854_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  OAI211_X1 g674(.A(KEYINPUT119), .B(new_n856_), .C1(new_n875_), .C2(new_n726_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n868_), .A2(new_n871_), .A3(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT122), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT122), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n868_), .A2(new_n871_), .A3(new_n879_), .A4(new_n876_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n880_), .ZN(G1340gat));
  INV_X1    g680(.A(G120gat), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n588_), .B1(new_n875_), .B2(KEYINPUT59), .ZN(new_n883_));
  AOI22_X1  g682(.A1(new_n859_), .A2(KEYINPUT121), .B1(KEYINPUT57), .B2(new_n858_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n609_), .B1(new_n884_), .B2(new_n862_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n866_), .B1(new_n885_), .B2(new_n799_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n882_), .B1(new_n883_), .B2(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n882_), .B1(new_n641_), .B2(KEYINPUT60), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n888_), .B1(KEYINPUT60), .B2(new_n882_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n875_), .A2(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(KEYINPUT123), .B1(new_n887_), .B2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n863_), .A2(new_n608_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n867_), .B1(new_n892_), .B2(new_n798_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n855_), .A2(new_n661_), .ZN(new_n894_));
  OAI21_X1  g693(.A(G120gat), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n896_));
  INV_X1    g695(.A(new_n890_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n895_), .A2(new_n896_), .A3(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n891_), .A2(new_n898_), .ZN(G1341gat));
  NAND2_X1  g698(.A1(new_n886_), .A2(new_n855_), .ZN(new_n900_));
  OAI21_X1  g699(.A(G127gat), .B1(new_n900_), .B2(new_n608_), .ZN(new_n901_));
  OR2_X1    g700(.A1(new_n608_), .A2(G127gat), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n875_), .B2(new_n902_), .ZN(G1342gat));
  OAI21_X1  g702(.A(G134gat), .B1(new_n900_), .B2(new_n634_), .ZN(new_n904_));
  OR2_X1    g703(.A1(new_n632_), .A2(G134gat), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n875_), .B2(new_n905_), .ZN(G1343gat));
  NOR4_X1   g705(.A1(new_n439_), .A2(new_n650_), .A3(new_n398_), .A4(new_n362_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n873_), .A2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(new_n483_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n661_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g712(.A(KEYINPUT124), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n909_), .A2(new_n914_), .A3(new_n609_), .ZN(new_n915_));
  OAI21_X1  g714(.A(KEYINPUT124), .B1(new_n908_), .B2(new_n608_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(KEYINPUT61), .B(G155gat), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n919_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n915_), .A2(new_n916_), .A3(new_n918_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(G1346gat));
  OR3_X1    g721(.A1(new_n908_), .A2(G162gat), .A3(new_n632_), .ZN(new_n923_));
  OAI21_X1  g722(.A(G162gat), .B1(new_n908_), .B2(new_n634_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1347gat));
  NOR3_X1   g724(.A1(new_n438_), .A2(new_n397_), .A3(new_n299_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(new_n362_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  OAI211_X1 g727(.A(new_n483_), .B(new_n928_), .C1(new_n885_), .C2(new_n799_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n930_));
  AND3_X1   g729(.A1(new_n929_), .A2(new_n930_), .A3(G169gat), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n929_), .B2(G169gat), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n928_), .B1(new_n885_), .B2(new_n799_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(KEYINPUT22), .B(G169gat), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n483_), .A2(new_n934_), .ZN(new_n935_));
  XOR2_X1   g734(.A(new_n935_), .B(KEYINPUT125), .Z(new_n936_));
  OAI22_X1  g735(.A1(new_n931_), .A2(new_n932_), .B1(new_n933_), .B2(new_n936_), .ZN(G1348gat));
  AOI21_X1  g736(.A(new_n927_), .B1(new_n892_), .B2(new_n798_), .ZN(new_n938_));
  AOI21_X1  g737(.A(G176gat), .B1(new_n938_), .B2(new_n640_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n873_), .A2(KEYINPUT126), .A3(new_n362_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT126), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n941_), .B1(new_n851_), .B2(new_n675_), .ZN(new_n942_));
  AND3_X1   g741(.A1(new_n940_), .A2(new_n942_), .A3(new_n926_), .ZN(new_n943_));
  AND2_X1   g742(.A1(new_n661_), .A2(G176gat), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n939_), .B1(new_n943_), .B2(new_n944_), .ZN(G1349gat));
  AOI21_X1  g744(.A(new_n244_), .B1(new_n943_), .B2(new_n609_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n608_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n946_), .B1(new_n938_), .B2(new_n947_), .ZN(G1350gat));
  INV_X1    g747(.A(G190gat), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n949_), .B1(new_n938_), .B2(new_n686_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n685_), .A2(new_n210_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n933_), .A2(new_n951_), .ZN(new_n952_));
  OAI21_X1  g751(.A(KEYINPUT127), .B1(new_n950_), .B2(new_n952_), .ZN(new_n953_));
  OAI21_X1  g752(.A(G190gat), .B1(new_n933_), .B2(new_n634_), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n938_), .A2(new_n210_), .A3(new_n685_), .ZN(new_n955_));
  INV_X1    g754(.A(KEYINPUT127), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n954_), .A2(new_n955_), .A3(new_n956_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n953_), .A2(new_n957_), .ZN(G1351gat));
  AND4_X1   g757(.A1(new_n650_), .A2(new_n873_), .A3(new_n436_), .A4(new_n438_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n959_), .A2(new_n483_), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n960_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g760(.A1(new_n959_), .A2(new_n661_), .ZN(new_n962_));
  XNOR2_X1  g761(.A(new_n962_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g762(.A1(new_n959_), .A2(new_n609_), .ZN(new_n964_));
  XNOR2_X1  g763(.A(KEYINPUT63), .B(G211gat), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n964_), .A2(new_n965_), .ZN(new_n966_));
  NOR2_X1   g765(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n966_), .B1(new_n964_), .B2(new_n967_), .ZN(G1354gat));
  INV_X1    g767(.A(G218gat), .ZN(new_n969_));
  NAND3_X1  g768(.A1(new_n959_), .A2(new_n969_), .A3(new_n685_), .ZN(new_n970_));
  AND2_X1   g769(.A1(new_n959_), .A2(new_n686_), .ZN(new_n971_));
  OAI21_X1  g770(.A(new_n970_), .B1(new_n971_), .B2(new_n969_), .ZN(G1355gat));
endmodule


