//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 0 0 0 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 1 1 0 0 0 0 1 1 0 0 0 0 1 1 0 1 0 0 0 0 0 0 0 0 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n886_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_;
  INV_X1    g000(.A(KEYINPUT12), .ZN(new_n202_));
  OR2_X1    g001(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n203_));
  INV_X1    g002(.A(G106gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT64), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT64), .ZN(new_n208_));
  NAND4_X1  g007(.A1(new_n203_), .A2(new_n208_), .A3(new_n204_), .A4(new_n205_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  AND3_X1   g009(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n211_));
  AOI21_X1  g010(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n212_));
  NOR3_X1   g011(.A1(new_n211_), .A2(new_n212_), .A3(KEYINPUT66), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT6), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n214_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n213_), .A2(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  AND2_X1   g020(.A1(G85gat), .A2(G92gat), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n221_), .B1(new_n222_), .B2(KEYINPUT9), .ZN(new_n223_));
  INV_X1    g022(.A(G85gat), .ZN(new_n224_));
  OR2_X1    g023(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n224_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n223_), .B1(new_n227_), .B2(KEYINPUT9), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n210_), .A2(new_n220_), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  NOR3_X1   g031(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n235_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n217_), .A2(KEYINPUT67), .A3(new_n218_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n234_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n222_), .A2(new_n221_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT68), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT68), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n238_), .A2(new_n242_), .A3(new_n239_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(KEYINPUT8), .A3(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n220_), .A2(new_n234_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT8), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(new_n246_), .A3(new_n239_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n230_), .B1(new_n244_), .B2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G57gat), .B(G64gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT69), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT11), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G71gat), .B(G78gat), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n249_), .A2(KEYINPUT69), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT11), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n249_), .A2(KEYINPUT69), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n254_), .A2(new_n255_), .A3(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n251_), .A2(new_n253_), .A3(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n250_), .A2(KEYINPUT11), .A3(new_n252_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n202_), .B1(new_n248_), .B2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G230gat), .A2(G233gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n243_), .A2(KEYINPUT8), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n242_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n247_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(new_n260_), .A3(new_n229_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n229_), .A2(KEYINPUT70), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n210_), .A2(new_n220_), .A3(new_n228_), .A4(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n265_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n258_), .A2(KEYINPUT12), .A3(new_n259_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n261_), .A2(new_n262_), .A3(new_n266_), .A4(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n260_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n248_), .B(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n275_), .B1(new_n277_), .B2(new_n262_), .ZN(new_n278_));
  XOR2_X1   g077(.A(G120gat), .B(G148gat), .Z(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT5), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G176gat), .B(G204gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n278_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n278_), .A2(new_n282_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n283_), .A2(KEYINPUT71), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n284_), .B1(new_n283_), .B2(KEYINPUT71), .ZN(new_n287_));
  NOR3_X1   g086(.A1(new_n286_), .A2(KEYINPUT13), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT13), .B1(new_n286_), .B2(new_n287_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n289_), .A2(KEYINPUT72), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT13), .ZN(new_n293_));
  INV_X1    g092(.A(new_n287_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n293_), .B1(new_n294_), .B2(new_n285_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n292_), .B1(new_n295_), .B2(new_n288_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT74), .B(G8gat), .ZN(new_n297_));
  INV_X1    g096(.A(G1gat), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT14), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G15gat), .B(G22gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT75), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G1gat), .B(G8gat), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n301_), .B(KEYINPUT75), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n304_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G29gat), .B(G36gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G43gat), .B(G50gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n310_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n309_), .A2(new_n313_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G229gat), .A2(G233gat), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n317_), .A2(KEYINPUT77), .A3(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n313_), .B(KEYINPUT15), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n310_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n322_), .A2(new_n318_), .A3(new_n316_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n320_), .A2(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(KEYINPUT77), .B1(new_n317_), .B2(new_n319_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G113gat), .B(G141gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G169gat), .B(G197gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n329_), .A2(KEYINPUT78), .ZN(new_n330_));
  OR3_X1    g129(.A1(new_n324_), .A2(new_n325_), .A3(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n330_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G231gat), .A2(G233gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n260_), .B(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(new_n309_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G127gat), .B(G155gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT16), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT76), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G183gat), .B(G211gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  XOR2_X1   g140(.A(new_n341_), .B(KEYINPUT17), .Z(new_n342_));
  OR2_X1    g141(.A1(new_n336_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(KEYINPUT17), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n336_), .A2(new_n344_), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n291_), .A2(new_n296_), .A3(new_n333_), .A4(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT100), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G127gat), .B(G134gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G113gat), .B(G120gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n354_));
  INV_X1    g153(.A(G169gat), .ZN(new_n355_));
  INV_X1    g154(.A(G176gat), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT80), .B1(G169gat), .B2(G176gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT24), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT81), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT23), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G183gat), .A2(G190gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(KEYINPUT81), .A2(KEYINPUT23), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n364_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n361_), .A2(KEYINPUT82), .A3(new_n367_), .A4(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT82), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n367_), .A2(new_n368_), .ZN(new_n371_));
  AOI21_X1  g170(.A(KEYINPUT24), .B1(new_n357_), .B2(new_n358_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n370_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT25), .B(G183gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT26), .B(G190gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G169gat), .A2(G176gat), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n357_), .A2(KEYINPUT24), .A3(new_n377_), .A4(new_n358_), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n369_), .A2(new_n373_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n365_), .A2(KEYINPUT23), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n364_), .A2(new_n366_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n381_), .B1(new_n382_), .B2(new_n365_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n383_), .B1(G183gat), .B2(G190gat), .ZN(new_n384_));
  INV_X1    g183(.A(new_n377_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT22), .B(G169gat), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n385_), .B1(new_n386_), .B2(new_n356_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n384_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n380_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT30), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G71gat), .B(G99gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(G43gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G227gat), .A2(G233gat), .ZN(new_n393_));
  INV_X1    g192(.A(G15gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n392_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n390_), .B(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT31), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n397_), .A2(KEYINPUT31), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n353_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n397_), .A2(KEYINPUT31), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(new_n352_), .A3(new_n398_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT84), .ZN(new_n404_));
  INV_X1    g203(.A(G155gat), .ZN(new_n405_));
  INV_X1    g204(.A(G162gat), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n404_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G155gat), .A2(G162gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT1), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT85), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n410_), .B2(KEYINPUT1), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT1), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n414_), .A2(KEYINPUT85), .A3(G155gat), .A4(G162gat), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n409_), .A2(new_n411_), .A3(new_n413_), .A4(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(G141gat), .ZN(new_n417_));
  INV_X1    g216(.A(G148gat), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n417_), .A2(new_n418_), .A3(KEYINPUT83), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT83), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n420_), .B1(G141gat), .B2(G148gat), .ZN(new_n421_));
  AOI22_X1  g220(.A1(new_n419_), .A2(new_n421_), .B1(G141gat), .B2(G148gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n416_), .A2(new_n422_), .ZN(new_n423_));
  OR3_X1    g222(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT2), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n425_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n424_), .A2(new_n426_), .A3(new_n427_), .A4(new_n428_), .ZN(new_n429_));
  AOI22_X1  g228(.A1(new_n407_), .A2(new_n408_), .B1(G155gat), .B2(G162gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n423_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT88), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(new_n433_), .A3(new_n353_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT4), .ZN(new_n435_));
  AOI22_X1  g234(.A1(new_n416_), .A2(new_n422_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n435_), .B1(new_n436_), .B2(new_n352_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n434_), .A2(new_n437_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n432_), .A2(new_n433_), .A3(new_n435_), .A4(new_n353_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G225gat), .A2(G233gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT87), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n438_), .A2(new_n439_), .A3(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n353_), .B(new_n436_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n440_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G1gat), .B(G29gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(KEYINPUT0), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(G57gat), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n446_), .A2(G57gat), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n224_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n446_), .A2(G57gat), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n451_), .A2(G85gat), .A3(new_n447_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n442_), .A2(new_n444_), .A3(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n453_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n401_), .A2(new_n403_), .A3(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT97), .ZN(new_n459_));
  XOR2_X1   g258(.A(G8gat), .B(G36gat), .Z(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT18), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G64gat), .B(G92gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT94), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(G197gat), .B(G204gat), .Z(new_n466_));
  XNOR2_X1  g265(.A(G211gat), .B(G218gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n466_), .B1(KEYINPUT21), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(KEYINPUT21), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n470_), .A2(new_n380_), .A3(new_n388_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT20), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n360_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n383_), .A2(new_n376_), .A3(new_n378_), .A4(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(G183gat), .A2(G190gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n387_), .B1(new_n371_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n467_), .A2(KEYINPUT21), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(new_n466_), .A3(new_n469_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n469_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n468_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n472_), .B1(new_n477_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G226gat), .A2(G233gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT19), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n471_), .A2(new_n483_), .A3(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT93), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n380_), .A2(new_n388_), .A3(new_n482_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n470_), .A2(new_n477_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n472_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n491_), .A2(new_n486_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n465_), .B1(new_n488_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n491_), .A2(new_n486_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n471_), .A2(new_n483_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(new_n485_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n494_), .A2(new_n463_), .A3(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT27), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n463_), .ZN(new_n500_));
  AOI211_X1 g299(.A(new_n472_), .B(new_n485_), .C1(new_n489_), .C2(new_n490_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n486_), .B1(new_n471_), .B2(new_n483_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n500_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(new_n497_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT27), .ZN(new_n505_));
  AOI22_X1  g304(.A1(new_n493_), .A2(new_n499_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G78gat), .B(G106gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n432_), .A2(KEYINPUT29), .ZN(new_n508_));
  INV_X1    g307(.A(G228gat), .ZN(new_n509_));
  INV_X1    g308(.A(G233gat), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n508_), .A2(new_n512_), .A3(new_n482_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n512_), .B1(new_n508_), .B2(new_n482_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n507_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n515_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n507_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(new_n513_), .A3(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n516_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n516_), .A2(KEYINPUT86), .ZN(new_n521_));
  XOR2_X1   g320(.A(G22gat), .B(G50gat), .Z(new_n522_));
  INV_X1    g321(.A(KEYINPUT28), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT29), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n436_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n523_), .B1(new_n436_), .B2(new_n524_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n522_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n527_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n522_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(new_n525_), .A3(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n528_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n520_), .A2(new_n521_), .A3(new_n533_), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n516_), .B(new_n519_), .C1(new_n532_), .C2(KEYINPUT86), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n506_), .A2(new_n536_), .ZN(new_n537_));
  OR3_X1    g336(.A1(new_n458_), .A2(new_n459_), .A3(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n459_), .B1(new_n458_), .B2(new_n537_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NOR3_X1   g339(.A1(new_n501_), .A2(new_n500_), .A3(new_n502_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n463_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n505_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT93), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n487_), .B(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n492_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n464_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n543_), .B1(new_n547_), .B2(new_n498_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n534_), .A2(new_n457_), .A3(new_n535_), .ZN(new_n549_));
  OAI21_X1  g348(.A(KEYINPUT95), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n534_), .A2(new_n457_), .A3(new_n535_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT95), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n506_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n550_), .A2(new_n553_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n442_), .A2(new_n444_), .A3(KEYINPUT33), .A4(new_n453_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT89), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n453_), .B1(new_n443_), .B2(new_n441_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n438_), .A2(new_n440_), .A3(new_n439_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(KEYINPUT91), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT91), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n438_), .A2(new_n561_), .A3(new_n440_), .A4(new_n439_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n558_), .A2(new_n560_), .A3(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT90), .B(KEYINPUT33), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n454_), .A2(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n563_), .A2(new_n565_), .A3(new_n497_), .A4(new_n503_), .ZN(new_n566_));
  OAI21_X1  g365(.A(KEYINPUT92), .B1(new_n557_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n457_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n463_), .A2(KEYINPUT32), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n569_), .B1(new_n488_), .B2(new_n492_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n494_), .A2(new_n496_), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n568_), .B(new_n570_), .C1(new_n571_), .C2(new_n569_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n555_), .B(KEYINPUT89), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n563_), .A2(new_n565_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n504_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT92), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .A4(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n567_), .A2(new_n572_), .A3(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n554_), .B1(new_n536_), .B2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n401_), .A2(new_n403_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  OAI21_X1  g380(.A(KEYINPUT96), .B1(new_n579_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n554_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n578_), .A2(new_n536_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT96), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(new_n586_), .A3(new_n580_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n540_), .B1(new_n582_), .B2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n271_), .A2(new_n321_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT34), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n265_), .A2(new_n229_), .ZN(new_n592_));
  OAI221_X1 g391(.A(new_n589_), .B1(KEYINPUT35), .B2(new_n591_), .C1(new_n314_), .C2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(KEYINPUT35), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(G190gat), .B(G218gat), .Z(new_n596_));
  XNOR2_X1  g395(.A(G134gat), .B(G162gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT36), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n595_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n598_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n603_), .A2(KEYINPUT36), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n595_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n602_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n588_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n349_), .A2(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(G1gat), .B1(new_n609_), .B2(new_n457_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n291_), .A2(new_n296_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n612_), .A2(KEYINPUT73), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n291_), .A2(KEYINPUT73), .A3(new_n296_), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n333_), .A2(KEYINPUT79), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT79), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n331_), .A2(new_n617_), .A3(new_n332_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(KEYINPUT98), .B1(new_n588_), .B2(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n538_), .A2(new_n539_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n586_), .B1(new_n585_), .B2(new_n580_), .ZN(new_n623_));
  AOI211_X1 g422(.A(KEYINPUT96), .B(new_n581_), .C1(new_n583_), .C2(new_n584_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n622_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT98), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n625_), .A2(new_n626_), .A3(new_n619_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n621_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT37), .ZN(new_n629_));
  INV_X1    g428(.A(new_n605_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n629_), .B1(new_n630_), .B2(new_n601_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n602_), .A2(KEYINPUT37), .A3(new_n605_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n634_), .A2(new_n346_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n615_), .A2(new_n628_), .A3(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n457_), .A2(G1gat), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT38), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n638_), .A2(KEYINPUT101), .A3(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(KEYINPUT101), .B1(new_n638_), .B2(new_n639_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n638_), .A2(new_n639_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n642_), .A2(KEYINPUT99), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n638_), .A2(new_n644_), .A3(new_n639_), .ZN(new_n645_));
  OAI221_X1 g444(.A(new_n610_), .B1(new_n640_), .B2(new_n641_), .C1(new_n643_), .C2(new_n645_), .ZN(G1324gat));
  NAND3_X1  g445(.A1(new_n636_), .A2(new_n548_), .A3(new_n297_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n349_), .A2(KEYINPUT102), .A3(new_n548_), .A4(new_n608_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n648_), .A2(G8gat), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT39), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n651_), .B1(new_n609_), .B2(new_n506_), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n649_), .A2(new_n650_), .A3(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n650_), .B1(new_n649_), .B2(new_n652_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n647_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  XOR2_X1   g454(.A(KEYINPUT103), .B(KEYINPUT40), .Z(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n656_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n647_), .B(new_n658_), .C1(new_n653_), .C2(new_n654_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(G1325gat));
  NAND3_X1  g459(.A1(new_n636_), .A2(new_n394_), .A3(new_n581_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n349_), .A2(new_n581_), .A3(new_n608_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(G15gat), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n663_), .A2(KEYINPUT105), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(KEYINPUT105), .ZN(new_n665_));
  XOR2_X1   g464(.A(KEYINPUT104), .B(KEYINPUT41), .Z(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n664_), .A2(new_n665_), .A3(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n667_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n661_), .B1(new_n668_), .B2(new_n669_), .ZN(G1326gat));
  OAI21_X1  g469(.A(G22gat), .B1(new_n609_), .B2(new_n536_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT42), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n536_), .A2(G22gat), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT106), .Z(new_n674_));
  NAND2_X1  g473(.A1(new_n636_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n672_), .A2(new_n675_), .ZN(G1327gat));
  NOR2_X1   g475(.A1(new_n606_), .A2(new_n347_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n612_), .A2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n678_), .B1(new_n627_), .B2(new_n621_), .ZN(new_n679_));
  AOI21_X1  g478(.A(G29gat), .B1(new_n679_), .B2(new_n568_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n291_), .A2(new_n333_), .A3(new_n296_), .ZN(new_n681_));
  OAI21_X1  g480(.A(KEYINPUT43), .B1(new_n588_), .B2(new_n633_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n625_), .A2(new_n683_), .A3(new_n634_), .ZN(new_n684_));
  AOI211_X1 g483(.A(new_n347_), .B(new_n681_), .C1(new_n682_), .C2(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n685_), .A2(KEYINPUT44), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n687_), .A2(G29gat), .A3(new_n568_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n682_), .A2(new_n684_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n681_), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n689_), .A2(KEYINPUT44), .A3(new_n346_), .A4(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT107), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n347_), .B1(new_n682_), .B2(new_n684_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n694_), .A2(KEYINPUT107), .A3(KEYINPUT44), .A4(new_n690_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n680_), .B1(new_n688_), .B2(new_n696_), .ZN(G1328gat));
  NOR2_X1   g496(.A1(new_n506_), .A2(G36gat), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n679_), .A2(new_n698_), .ZN(new_n699_));
  XOR2_X1   g498(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n700_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n679_), .A2(new_n698_), .A3(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n548_), .B1(new_n685_), .B2(KEYINPUT44), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n693_), .B2(new_n695_), .ZN(new_n707_));
  INV_X1    g506(.A(G36gat), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n705_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT46), .B1(new_n709_), .B2(KEYINPUT109), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n694_), .A2(new_n690_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n506_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n708_), .B1(new_n696_), .B2(new_n713_), .ZN(new_n714_));
  OAI211_X1 g513(.A(KEYINPUT109), .B(KEYINPUT46), .C1(new_n714_), .C2(new_n704_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n710_), .A2(new_n716_), .ZN(G1329gat));
  NAND4_X1  g516(.A1(new_n696_), .A2(new_n687_), .A3(G43gat), .A4(new_n581_), .ZN(new_n718_));
  AOI21_X1  g517(.A(G43gat), .B1(new_n679_), .B2(new_n581_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g521(.A(new_n536_), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n696_), .A2(new_n687_), .A3(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(G50gat), .ZN(new_n725_));
  INV_X1    g524(.A(new_n679_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n536_), .A2(G50gat), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT110), .ZN(new_n728_));
  OAI22_X1  g527(.A1(new_n724_), .A2(new_n725_), .B1(new_n726_), .B2(new_n728_), .ZN(G1331gat));
  INV_X1    g528(.A(G57gat), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n611_), .A2(new_n635_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT111), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n731_), .B(new_n732_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n588_), .A2(new_n333_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n730_), .B1(new_n735_), .B2(new_n457_), .ZN(new_n736_));
  OR2_X1    g535(.A1(new_n736_), .A2(KEYINPUT112), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(KEYINPUT112), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n613_), .A2(new_n614_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n346_), .B1(new_n616_), .B2(new_n618_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  XOR2_X1   g540(.A(KEYINPUT113), .B(G57gat), .Z(new_n742_));
  NAND4_X1  g541(.A1(new_n741_), .A2(new_n568_), .A3(new_n608_), .A4(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n737_), .A2(new_n738_), .A3(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT114), .ZN(G1332gat));
  NAND3_X1  g544(.A1(new_n741_), .A2(new_n548_), .A3(new_n608_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(G64gat), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n747_), .A2(KEYINPUT48), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(KEYINPUT48), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n506_), .A2(G64gat), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT115), .ZN(new_n751_));
  OAI22_X1  g550(.A1(new_n748_), .A2(new_n749_), .B1(new_n735_), .B2(new_n751_), .ZN(G1333gat));
  OR3_X1    g551(.A1(new_n735_), .A2(G71gat), .A3(new_n580_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n741_), .A2(new_n581_), .A3(new_n608_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(G71gat), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n755_), .A2(KEYINPUT49), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(KEYINPUT49), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n753_), .B1(new_n756_), .B2(new_n757_), .ZN(G1334gat));
  OR3_X1    g557(.A1(new_n735_), .A2(G78gat), .A3(new_n536_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n741_), .A2(new_n723_), .A3(new_n608_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(G78gat), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n761_), .A2(KEYINPUT50), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(KEYINPUT50), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n759_), .B1(new_n762_), .B2(new_n763_), .ZN(G1335gat));
  AND2_X1   g563(.A1(new_n739_), .A2(new_n677_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n765_), .A2(new_n734_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n766_), .A2(new_n224_), .A3(new_n568_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n612_), .A2(new_n333_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n694_), .A2(new_n768_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n769_), .A2(new_n568_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n767_), .B1(new_n224_), .B2(new_n770_), .ZN(G1336gat));
  AOI21_X1  g570(.A(G92gat), .B1(new_n766_), .B2(new_n548_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n506_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n769_), .B2(new_n773_), .ZN(G1337gat));
  NAND4_X1  g573(.A1(new_n766_), .A2(new_n581_), .A3(new_n203_), .A4(new_n205_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n769_), .A2(new_n581_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n776_), .A2(KEYINPUT116), .A3(G99gat), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT116), .B1(new_n776_), .B2(G99gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n775_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT51), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n775_), .B(new_n781_), .C1(new_n777_), .C2(new_n778_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(G1338gat));
  AOI21_X1  g582(.A(new_n204_), .B1(new_n769_), .B2(new_n723_), .ZN(new_n784_));
  OR2_X1    g583(.A1(new_n784_), .A2(KEYINPUT52), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n536_), .A2(G106gat), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n765_), .A2(new_n734_), .A3(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT117), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n765_), .A2(KEYINPUT117), .A3(new_n734_), .A4(new_n786_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n784_), .A2(KEYINPUT52), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n785_), .A2(new_n791_), .A3(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT53), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n785_), .A2(new_n791_), .A3(new_n795_), .A4(new_n792_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(G1339gat));
  NOR3_X1   g596(.A1(new_n580_), .A2(new_n457_), .A3(new_n537_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n333_), .A2(new_n283_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT118), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n275_), .B2(new_n802_), .ZN(new_n803_));
  AOI22_X1  g602(.A1(new_n244_), .A2(new_n247_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n266_), .B1(new_n804_), .B2(new_n272_), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT12), .B1(new_n592_), .B2(new_n276_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n807_), .A2(KEYINPUT118), .A3(KEYINPUT55), .A4(new_n262_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n803_), .A2(new_n808_), .ZN(new_n809_));
  AOI22_X1  g608(.A1(new_n271_), .A2(new_n273_), .B1(new_n248_), .B2(new_n260_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n262_), .B1(new_n810_), .B2(new_n261_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n802_), .B2(new_n275_), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n809_), .A2(KEYINPUT119), .A3(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT119), .B1(new_n809_), .B2(new_n812_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n282_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT56), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  OAI211_X1 g616(.A(KEYINPUT56), .B(new_n282_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n800_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n329_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n322_), .A2(new_n319_), .A3(new_n316_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n319_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n328_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n820_), .A2(new_n823_), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n294_), .A2(new_n285_), .A3(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n606_), .B1(new_n819_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n824_), .A2(new_n283_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n829_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n633_), .B1(new_n830_), .B2(KEYINPUT58), .ZN(new_n831_));
  INV_X1    g630(.A(new_n829_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n809_), .A2(new_n812_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n809_), .A2(KEYINPUT119), .A3(new_n812_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(KEYINPUT56), .B1(new_n837_), .B2(new_n282_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n818_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n832_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT58), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n831_), .A2(new_n842_), .ZN(new_n843_));
  OAI211_X1 g642(.A(KEYINPUT57), .B(new_n606_), .C1(new_n819_), .C2(new_n825_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n828_), .A2(new_n843_), .A3(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n346_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n740_), .A2(new_n633_), .A3(new_n290_), .A4(new_n289_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n847_), .B(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n799_), .B1(new_n846_), .B2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(G113gat), .B1(new_n851_), .B2(new_n333_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT121), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n851_), .B2(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n849_), .B1(new_n845_), .B2(new_n346_), .ZN(new_n857_));
  OAI211_X1 g656(.A(KEYINPUT120), .B(KEYINPUT59), .C1(new_n857_), .C2(new_n799_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n858_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n857_), .A2(KEYINPUT59), .A3(new_n799_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n853_), .B1(new_n859_), .B2(new_n861_), .ZN(new_n862_));
  AOI211_X1 g661(.A(KEYINPUT121), .B(new_n860_), .C1(new_n856_), .C2(new_n858_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n619_), .A2(G113gat), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n852_), .B1(new_n864_), .B2(new_n865_), .ZN(G1340gat));
  AOI211_X1 g665(.A(new_n615_), .B(new_n860_), .C1(new_n856_), .C2(new_n858_), .ZN(new_n867_));
  INV_X1    g666(.A(G120gat), .ZN(new_n868_));
  INV_X1    g667(.A(new_n851_), .ZN(new_n869_));
  NOR3_X1   g668(.A1(new_n612_), .A2(KEYINPUT60), .A3(G120gat), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n870_), .B1(KEYINPUT60), .B2(G120gat), .ZN(new_n871_));
  OAI22_X1  g670(.A1(new_n867_), .A2(new_n868_), .B1(new_n869_), .B2(new_n871_), .ZN(G1341gat));
  AOI21_X1  g671(.A(G127gat), .B1(new_n851_), .B2(new_n347_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n347_), .A2(G127gat), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n873_), .B1(new_n864_), .B2(new_n874_), .ZN(G1342gat));
  AOI21_X1  g674(.A(G134gat), .B1(new_n851_), .B2(new_n607_), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n634_), .A2(G134gat), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n876_), .B1(new_n864_), .B2(new_n877_), .ZN(G1343gat));
  NOR2_X1   g677(.A1(new_n857_), .A2(new_n581_), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n548_), .A2(new_n536_), .A3(new_n457_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n333_), .ZN(new_n883_));
  XOR2_X1   g682(.A(KEYINPUT122), .B(G141gat), .Z(new_n884_));
  XNOR2_X1  g683(.A(new_n883_), .B(new_n884_), .ZN(G1344gat));
  NOR2_X1   g684(.A1(new_n881_), .A2(new_n615_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(new_n418_), .ZN(G1345gat));
  NAND2_X1  g686(.A1(new_n882_), .A2(new_n347_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT61), .B(G155gat), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1346gat));
  OAI21_X1  g689(.A(G162gat), .B1(new_n881_), .B2(new_n633_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n607_), .A2(new_n406_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n881_), .B2(new_n892_), .ZN(G1347gat));
  NAND2_X1  g692(.A1(new_n846_), .A2(new_n850_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n458_), .A2(new_n723_), .A3(new_n506_), .ZN(new_n895_));
  AND2_X1   g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n896_), .A2(new_n386_), .A3(new_n333_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n333_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n898_), .A2(new_n899_), .A3(G169gat), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n898_), .B2(G169gat), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT123), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n900_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  AOI211_X1 g702(.A(KEYINPUT123), .B(new_n899_), .C1(new_n898_), .C2(G169gat), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n897_), .B1(new_n903_), .B2(new_n904_), .ZN(G1348gat));
  NAND3_X1  g704(.A1(new_n896_), .A2(new_n356_), .A3(new_n611_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n894_), .A2(new_n895_), .ZN(new_n907_));
  OAI21_X1  g706(.A(G176gat), .B1(new_n907_), .B2(new_n615_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n908_), .ZN(G1349gat));
  OR2_X1    g708(.A1(KEYINPUT124), .A2(G183gat), .ZN(new_n910_));
  NAND4_X1  g709(.A1(new_n896_), .A2(new_n374_), .A3(new_n347_), .A4(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT124), .ZN(new_n912_));
  OAI22_X1  g711(.A1(new_n907_), .A2(new_n346_), .B1(new_n912_), .B2(G183gat), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n911_), .A2(new_n913_), .ZN(new_n914_));
  XOR2_X1   g713(.A(new_n914_), .B(KEYINPUT125), .Z(G1350gat));
  OAI21_X1  g714(.A(G190gat), .B1(new_n907_), .B2(new_n633_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n607_), .A2(new_n375_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(KEYINPUT126), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n916_), .B1(new_n907_), .B2(new_n918_), .ZN(G1351gat));
  NOR2_X1   g718(.A1(new_n506_), .A2(new_n549_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n879_), .A2(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(new_n333_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g723(.A1(new_n921_), .A2(new_n615_), .ZN(new_n925_));
  XOR2_X1   g724(.A(KEYINPUT127), .B(G204gat), .Z(new_n926_));
  XNOR2_X1  g725(.A(new_n925_), .B(new_n926_), .ZN(G1353gat));
  AOI21_X1  g726(.A(new_n346_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n922_), .A2(new_n928_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n930_));
  XOR2_X1   g729(.A(new_n929_), .B(new_n930_), .Z(G1354gat));
  OR3_X1    g730(.A1(new_n921_), .A2(G218gat), .A3(new_n606_), .ZN(new_n932_));
  OAI21_X1  g731(.A(G218gat), .B1(new_n921_), .B2(new_n633_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1355gat));
endmodule


