//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n884_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n901_, new_n903_, new_n904_, new_n905_, new_n907_,
    new_n908_, new_n909_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_, new_n921_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(KEYINPUT86), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n202_), .B(new_n203_), .ZN(new_n206_));
  AOI21_X1  g005(.A(new_n205_), .B1(new_n206_), .B2(KEYINPUT86), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT87), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT85), .B(G43gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT23), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT24), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n213_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(KEYINPUT24), .A3(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT26), .B(G190gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n220_), .A2(KEYINPUT84), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT25), .B(G183gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT84), .ZN(new_n223_));
  INV_X1    g022(.A(G190gat), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n224_), .A2(KEYINPUT26), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n222_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n216_), .B(new_n219_), .C1(new_n221_), .C2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n212_), .B1(G183gat), .B2(G190gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(G169gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n227_), .A2(KEYINPUT30), .A3(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT30), .B1(new_n227_), .B2(new_n231_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n210_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NOR3_X1   g035(.A1(new_n233_), .A2(new_n234_), .A3(new_n210_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n208_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n237_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n208_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n240_), .A3(new_n235_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G227gat), .A2(G233gat), .ZN(new_n243_));
  INV_X1    g042(.A(G15gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(G71gat), .ZN(new_n246_));
  INV_X1    g045(.A(G99gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT31), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n242_), .A2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n238_), .A2(new_n241_), .A3(new_n249_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G226gat), .A2(G233gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT19), .ZN(new_n256_));
  XOR2_X1   g055(.A(new_n256_), .B(KEYINPUT93), .Z(new_n257_));
  INV_X1    g056(.A(G204gat), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT90), .B1(new_n258_), .B2(G197gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT90), .ZN(new_n260_));
  INV_X1    g059(.A(G197gat), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(new_n261_), .A3(G204gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n258_), .A2(G197gat), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n259_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  XOR2_X1   g063(.A(G211gat), .B(G218gat), .Z(new_n265_));
  NAND3_X1  g064(.A1(new_n264_), .A2(KEYINPUT21), .A3(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n266_), .B(KEYINPUT92), .Z(new_n267_));
  NOR2_X1   g066(.A1(new_n264_), .A2(KEYINPUT21), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT91), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n261_), .A2(G204gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(new_n263_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n265_), .B1(KEYINPUT21), .B2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n267_), .B1(new_n269_), .B2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n222_), .B(KEYINPUT94), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(new_n220_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n219_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT95), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n275_), .A2(KEYINPUT95), .A3(new_n219_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(new_n279_), .A3(new_n216_), .ZN(new_n280_));
  OR2_X1    g079(.A1(new_n228_), .A2(KEYINPUT97), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n228_), .A2(KEYINPUT97), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n230_), .A2(KEYINPUT96), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n230_), .A2(KEYINPUT96), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n281_), .A2(new_n282_), .A3(new_n283_), .A4(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n273_), .B1(new_n280_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n267_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n269_), .A2(new_n272_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n227_), .A2(new_n231_), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT20), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n257_), .B1(new_n286_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT20), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n293_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n273_), .A2(new_n280_), .A3(new_n285_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n256_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n294_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n292_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G8gat), .B(G36gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT18), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G64gat), .B(G92gat), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n300_), .B(new_n301_), .Z(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n298_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n292_), .A2(new_n297_), .A3(new_n302_), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n304_), .A2(KEYINPUT98), .A3(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT98), .B1(new_n304_), .B2(new_n305_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(G1gat), .B(G29gat), .Z(new_n309_));
  XNOR2_X1  g108(.A(G57gat), .B(G85gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n311_), .B(new_n312_), .Z(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(G155gat), .ZN(new_n315_));
  INV_X1    g114(.A(G162gat), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT1), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT1), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(G155gat), .A3(G162gat), .ZN(new_n319_));
  NOR2_X1   g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n317_), .A2(new_n319_), .A3(new_n321_), .ZN(new_n322_));
  OR2_X1    g121(.A1(G141gat), .A2(G148gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G141gat), .A2(G148gat), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n322_), .A2(new_n323_), .A3(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT88), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n315_), .A2(new_n316_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n327_), .A2(new_n320_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n323_), .B(KEYINPUT3), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n324_), .B(KEYINPUT2), .Z(new_n330_));
  OAI21_X1  g129(.A(new_n328_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n326_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n208_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n332_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(new_n206_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT4), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G225gat), .A2(G233gat), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(KEYINPUT4), .B1(new_n208_), .B2(new_n332_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n337_), .A2(new_n339_), .A3(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n336_), .A2(new_n338_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n314_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n314_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n337_), .A2(new_n341_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n345_), .B1(new_n346_), .B2(new_n338_), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT33), .B1(new_n344_), .B2(new_n347_), .ZN(new_n348_));
  AOI211_X1 g147(.A(new_n338_), .B(new_n340_), .C1(new_n336_), .C2(KEYINPUT4), .ZN(new_n349_));
  INV_X1    g148(.A(new_n343_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n313_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT33), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n348_), .A2(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n308_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n342_), .A2(new_n314_), .A3(new_n343_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n351_), .A2(KEYINPUT100), .A3(new_n356_), .ZN(new_n357_));
  NOR3_X1   g156(.A1(new_n286_), .A2(new_n291_), .A3(new_n257_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n296_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n359_));
  OAI211_X1 g158(.A(KEYINPUT32), .B(new_n302_), .C1(new_n358_), .C2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n302_), .A2(KEYINPUT32), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n292_), .A2(new_n297_), .A3(new_n361_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT100), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n364_), .B(new_n313_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n357_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G228gat), .A2(G233gat), .ZN(new_n367_));
  INV_X1    g166(.A(G78gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(G106gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n326_), .A2(new_n372_), .A3(new_n331_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT28), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n373_), .A2(KEYINPUT28), .ZN(new_n376_));
  NOR3_X1   g175(.A1(new_n375_), .A2(new_n376_), .A3(KEYINPUT89), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT89), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n373_), .A2(KEYINPUT28), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n378_), .B1(new_n379_), .B2(new_n374_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n371_), .B1(new_n377_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n332_), .A2(KEYINPUT29), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n289_), .A2(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(G22gat), .B(G50gat), .Z(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n383_), .B(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(KEYINPUT89), .B1(new_n375_), .B2(new_n376_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n371_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n379_), .A2(new_n378_), .A3(new_n374_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n387_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  AND3_X1   g189(.A1(new_n381_), .A2(new_n386_), .A3(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n386_), .B1(new_n381_), .B2(new_n390_), .ZN(new_n392_));
  OR2_X1    g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n366_), .A2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n254_), .B1(new_n355_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT27), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n292_), .A2(new_n297_), .A3(new_n302_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n302_), .B1(new_n292_), .B2(new_n297_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n397_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT102), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT102), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n402_), .B(new_n397_), .C1(new_n398_), .C2(new_n399_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n303_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(KEYINPUT101), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT101), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n406_), .B(new_n303_), .C1(new_n358_), .C2(new_n359_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n398_), .A2(new_n397_), .ZN(new_n409_));
  AOI22_X1  g208(.A1(new_n401_), .A2(new_n403_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n357_), .A2(new_n365_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n393_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT103), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n253_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n415_), .B1(new_n365_), .B2(new_n357_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n414_), .B1(new_n410_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n410_), .A2(new_n416_), .A3(new_n414_), .ZN(new_n419_));
  AOI22_X1  g218(.A1(new_n396_), .A2(new_n413_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G1gat), .B(G8gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT81), .ZN(new_n422_));
  INV_X1    g221(.A(G22gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n244_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G15gat), .A2(G22gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G1gat), .A2(G8gat), .ZN(new_n426_));
  AOI22_X1  g225(.A1(new_n424_), .A2(new_n425_), .B1(KEYINPUT14), .B2(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n422_), .B(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G57gat), .B(G64gat), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n429_), .A2(KEYINPUT11), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(KEYINPUT11), .ZN(new_n431_));
  XOR2_X1   g230(.A(G71gat), .B(G78gat), .Z(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n431_), .A2(new_n432_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n428_), .B(new_n435_), .ZN(new_n436_));
  AND2_X1   g235(.A1(G231gat), .A2(G233gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  XOR2_X1   g238(.A(G127gat), .B(G155gat), .Z(new_n440_));
  XNOR2_X1  g239(.A(G183gat), .B(G211gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(KEYINPUT70), .A3(KEYINPUT17), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n439_), .A2(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n446_), .B1(KEYINPUT17), .B2(new_n445_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n438_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT80), .B(KEYINPUT37), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  XOR2_X1   g252(.A(KEYINPUT10), .B(G99gat), .Z(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n370_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT64), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G99gat), .A2(G106gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(G85gat), .ZN(new_n461_));
  INV_X1    g260(.A(G92gat), .ZN(new_n462_));
  NOR3_X1   g261(.A1(new_n461_), .A2(new_n462_), .A3(KEYINPUT9), .ZN(new_n463_));
  XOR2_X1   g262(.A(G85gat), .B(G92gat), .Z(new_n464_));
  AOI21_X1  g263(.A(new_n463_), .B1(new_n464_), .B2(KEYINPUT9), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n457_), .A2(new_n460_), .A3(new_n465_), .ZN(new_n466_));
  XOR2_X1   g265(.A(KEYINPUT65), .B(KEYINPUT6), .Z(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(new_n459_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n459_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n458_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT66), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n471_), .A2(new_n247_), .A3(new_n370_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT7), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT7), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n471_), .A2(new_n474_), .A3(new_n247_), .A4(new_n370_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n468_), .A2(new_n470_), .A3(new_n473_), .A4(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT8), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n464_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n476_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT67), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n481_), .A2(KEYINPUT6), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT6), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n483_), .A2(KEYINPUT67), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n459_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(KEYINPUT67), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n481_), .A2(KEYINPUT6), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n469_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n485_), .A2(new_n473_), .A3(new_n475_), .A4(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n477_), .B1(new_n489_), .B2(new_n464_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n480_), .B1(new_n490_), .B2(KEYINPUT68), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT68), .ZN(new_n492_));
  AOI211_X1 g291(.A(new_n492_), .B(new_n477_), .C1(new_n489_), .C2(new_n464_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n466_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT69), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(G36gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(G29gat), .ZN(new_n498_));
  INV_X1    g297(.A(G29gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(G36gat), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n498_), .A2(new_n500_), .A3(KEYINPUT76), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT76), .B1(new_n498_), .B2(new_n500_), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT77), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n498_), .A2(new_n500_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT76), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT77), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(new_n508_), .A3(new_n501_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G43gat), .B(G50gat), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n504_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n510_), .B1(new_n504_), .B2(new_n509_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT15), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT15), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n515_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  OAI211_X1 g316(.A(KEYINPUT69), .B(new_n466_), .C1(new_n491_), .C2(new_n493_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n496_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n455_), .B(KEYINPUT64), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n460_), .A2(new_n465_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n473_), .A2(new_n475_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n478_), .B1(new_n460_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n489_), .A2(new_n464_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT8), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n524_), .B1(new_n526_), .B2(new_n492_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n493_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n522_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT35), .ZN(new_n530_));
  NAND2_X1  g329(.A1(G232gat), .A2(G233gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT34), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  AOI22_X1  g332(.A1(new_n529_), .A2(new_n513_), .B1(new_n530_), .B2(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n533_), .A2(new_n530_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n519_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n536_), .B1(new_n519_), .B2(new_n534_), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT79), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT36), .B1(new_n538_), .B2(new_n539_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G190gat), .B(G218gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT78), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(G134gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(G162gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n541_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n545_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT36), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n540_), .B1(new_n546_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT36), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n519_), .A2(new_n534_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n535_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n550_), .B1(new_n552_), .B2(new_n537_), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n540_), .B(new_n548_), .C1(new_n553_), .C2(new_n547_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n453_), .B1(new_n549_), .B2(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n548_), .B1(new_n553_), .B2(new_n547_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n540_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n559_), .A2(new_n554_), .A3(new_n452_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n556_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NOR3_X1   g361(.A1(new_n420_), .A2(new_n451_), .A3(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT12), .B1(new_n435_), .B2(KEYINPUT70), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n564_), .B1(KEYINPUT70), .B2(new_n435_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n496_), .A2(new_n518_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n435_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n494_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT12), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n435_), .B(new_n466_), .C1(new_n491_), .C2(new_n493_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G230gat), .A2(G233gat), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n566_), .A2(new_n570_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT71), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n568_), .A2(new_n571_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n572_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n566_), .A2(new_n570_), .A3(KEYINPUT71), .A4(new_n573_), .ZN(new_n580_));
  XOR2_X1   g379(.A(G120gat), .B(G148gat), .Z(new_n581_));
  XNOR2_X1  g380(.A(G176gat), .B(G204gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n576_), .A2(new_n579_), .A3(new_n580_), .A4(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(KEYINPUT73), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n576_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT74), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n589_), .A2(new_n590_), .A3(new_n585_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n590_), .B1(new_n589_), .B2(new_n585_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n588_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n589_), .A2(new_n585_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT74), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n587_), .A2(KEYINPUT73), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n589_), .A2(new_n590_), .A3(new_n585_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n595_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n593_), .A2(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(KEYINPUT75), .A2(KEYINPUT13), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT75), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT13), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n599_), .A2(new_n601_), .A3(new_n605_), .ZN(new_n606_));
  NAND4_X1  g405(.A1(new_n593_), .A2(new_n598_), .A3(new_n602_), .A4(new_n603_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(G229gat), .A2(G233gat), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n513_), .A2(new_n428_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n513_), .A2(new_n428_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n609_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n428_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n517_), .A2(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n612_), .A2(new_n609_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n613_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G113gat), .B(G141gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G169gat), .B(G197gat), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n618_), .B(new_n619_), .Z(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT83), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n617_), .B(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n608_), .A2(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n563_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(G1gat), .ZN(new_n627_));
  INV_X1    g426(.A(new_n411_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n626_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n559_), .A2(KEYINPUT105), .A3(new_n554_), .ZN(new_n632_));
  AOI21_X1  g431(.A(KEYINPUT105), .B1(new_n559_), .B2(new_n554_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n634_), .A2(KEYINPUT106), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(KEYINPUT106), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n410_), .A2(new_n416_), .A3(new_n414_), .ZN(new_n639_));
  OAI22_X1  g438(.A1(new_n395_), .A2(new_n412_), .B1(new_n639_), .B2(new_n417_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n638_), .A2(new_n450_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n625_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT107), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n644_), .A2(new_n628_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n631_), .B1(new_n645_), .B2(new_n627_), .ZN(G1324gat));
  INV_X1    g445(.A(G8gat), .ZN(new_n647_));
  INV_X1    g446(.A(new_n410_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n626_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n647_), .B1(new_n643_), .B2(new_n648_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n650_), .A2(new_n651_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n649_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT40), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  OAI211_X1 g455(.A(KEYINPUT40), .B(new_n649_), .C1(new_n652_), .C2(new_n653_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1325gat));
  NAND3_X1  g457(.A1(new_n626_), .A2(new_n244_), .A3(new_n253_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n644_), .A2(new_n253_), .ZN(new_n660_));
  AOI21_X1  g459(.A(KEYINPUT41), .B1(new_n660_), .B2(G15gat), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT41), .ZN(new_n662_));
  AOI211_X1 g461(.A(new_n662_), .B(new_n244_), .C1(new_n644_), .C2(new_n253_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n659_), .B1(new_n661_), .B2(new_n663_), .ZN(G1326gat));
  INV_X1    g463(.A(new_n393_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n626_), .A2(new_n423_), .A3(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(KEYINPUT108), .B(KEYINPUT42), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n644_), .A2(new_n665_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n667_), .B1(new_n668_), .B2(G22gat), .ZN(new_n669_));
  INV_X1    g468(.A(new_n667_), .ZN(new_n670_));
  AOI211_X1 g469(.A(new_n423_), .B(new_n670_), .C1(new_n644_), .C2(new_n665_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n666_), .B1(new_n669_), .B2(new_n671_), .ZN(G1327gat));
  NOR2_X1   g471(.A1(new_n634_), .A2(new_n450_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n625_), .A2(new_n640_), .A3(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(G29gat), .B1(new_n674_), .B2(new_n628_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n625_), .A2(new_n451_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT109), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n625_), .A2(KEYINPUT109), .A3(new_n451_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT43), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n640_), .A2(new_n681_), .A3(new_n562_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT110), .ZN(new_n683_));
  OAI21_X1  g482(.A(KEYINPUT43), .B1(new_n420_), .B2(new_n561_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT110), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n640_), .A2(new_n685_), .A3(new_n681_), .A4(new_n562_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n683_), .A2(new_n684_), .A3(new_n686_), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n680_), .A2(new_n687_), .A3(KEYINPUT44), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT44), .B1(new_n680_), .B2(new_n687_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n411_), .A2(new_n499_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n675_), .B1(new_n690_), .B2(new_n691_), .ZN(G1328gat));
  NOR2_X1   g491(.A1(new_n410_), .A2(G36gat), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n674_), .A2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT111), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT111), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n674_), .A2(new_n696_), .A3(new_n693_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n695_), .A2(KEYINPUT45), .A3(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n695_), .A2(new_n697_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT45), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n688_), .A2(new_n689_), .A3(new_n410_), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n698_), .B(new_n701_), .C1(new_n702_), .C2(new_n497_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT46), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n701_), .A2(new_n698_), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n706_), .B(KEYINPUT46), .C1(new_n702_), .C2(new_n497_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(G1329gat));
  INV_X1    g507(.A(G43gat), .ZN(new_n709_));
  NOR4_X1   g508(.A1(new_n688_), .A2(new_n689_), .A3(new_n709_), .A4(new_n254_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n674_), .A2(new_n253_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n709_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n711_), .A2(new_n713_), .A3(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n714_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n713_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(new_n710_), .B2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n715_), .A2(new_n718_), .ZN(G1330gat));
  AOI21_X1  g518(.A(G50gat), .B1(new_n674_), .B2(new_n665_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n665_), .A2(G50gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n690_), .B2(new_n721_), .ZN(G1331gat));
  AOI21_X1  g521(.A(new_n623_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n563_), .A2(new_n723_), .ZN(new_n724_));
  OR3_X1    g523(.A1(new_n724_), .A2(G57gat), .A3(new_n411_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n638_), .A2(new_n450_), .A3(new_n640_), .A4(new_n723_), .ZN(new_n726_));
  OAI21_X1  g525(.A(G57gat), .B1(new_n726_), .B2(new_n411_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(new_n727_), .ZN(G1332gat));
  OAI21_X1  g527(.A(G64gat), .B1(new_n726_), .B2(new_n410_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT48), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n410_), .A2(G64gat), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT113), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n730_), .B1(new_n724_), .B2(new_n732_), .ZN(G1333gat));
  OAI21_X1  g532(.A(G71gat), .B1(new_n726_), .B2(new_n254_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT49), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n254_), .A2(G71gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n735_), .B1(new_n724_), .B2(new_n736_), .ZN(G1334gat));
  OAI21_X1  g536(.A(G78gat), .B1(new_n726_), .B2(new_n393_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT50), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n665_), .A2(new_n368_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n724_), .B2(new_n740_), .ZN(G1335gat));
  NAND2_X1  g540(.A1(new_n723_), .A2(new_n451_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n742_), .A2(KEYINPUT114), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n742_), .A2(KEYINPUT114), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n687_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G85gat), .B1(new_n745_), .B2(new_n411_), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n640_), .A2(new_n723_), .A3(new_n673_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n747_), .A2(new_n461_), .A3(new_n628_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n746_), .A2(new_n748_), .ZN(G1336gat));
  AOI21_X1  g548(.A(G92gat), .B1(new_n747_), .B2(new_n648_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n745_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n410_), .A2(new_n462_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT115), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n750_), .B1(new_n751_), .B2(new_n753_), .ZN(G1337gat));
  NAND2_X1  g553(.A1(new_n751_), .A2(new_n253_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n253_), .A2(new_n454_), .ZN(new_n756_));
  AOI22_X1  g555(.A1(new_n755_), .A2(G99gat), .B1(new_n747_), .B2(new_n756_), .ZN(new_n757_));
  XOR2_X1   g556(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n758_));
  XNOR2_X1  g557(.A(new_n757_), .B(new_n758_), .ZN(G1338gat));
  OAI21_X1  g558(.A(G106gat), .B1(new_n745_), .B2(new_n393_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n747_), .A2(new_n370_), .A3(new_n665_), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT117), .Z(new_n764_));
  OAI211_X1 g563(.A(KEYINPUT52), .B(G106gat), .C1(new_n745_), .C2(new_n393_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n762_), .A2(new_n764_), .A3(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT53), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT53), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n762_), .A2(new_n764_), .A3(new_n768_), .A4(new_n765_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1339gat));
  NAND2_X1  g569(.A1(new_n410_), .A2(new_n628_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n771_), .A2(new_n415_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n612_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n609_), .B1(new_n773_), .B2(new_n610_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n621_), .ZN(new_n775_));
  OR2_X1    g574(.A1(new_n775_), .A2(KEYINPUT119), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n773_), .A2(new_n609_), .ZN(new_n777_));
  AOI22_X1  g576(.A1(new_n775_), .A2(KEYINPUT119), .B1(new_n615_), .B2(new_n777_), .ZN(new_n778_));
  AOI22_X1  g577(.A1(new_n776_), .A2(new_n778_), .B1(new_n620_), .B2(new_n617_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n587_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n576_), .A2(new_n781_), .A3(new_n580_), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n566_), .A2(new_n570_), .A3(new_n573_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n566_), .A2(new_n571_), .A3(new_n570_), .ZN(new_n784_));
  AOI22_X1  g583(.A1(new_n783_), .A2(KEYINPUT55), .B1(new_n784_), .B2(new_n578_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n586_), .B1(new_n782_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT56), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n780_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT58), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT121), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n782_), .A2(new_n785_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n585_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT56), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n788_), .A2(new_n790_), .A3(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n790_), .B1(new_n788_), .B2(new_n793_), .ZN(new_n795_));
  NOR3_X1   g594(.A1(new_n794_), .A2(new_n561_), .A3(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT122), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n593_), .A2(new_n598_), .A3(new_n779_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT118), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n792_), .A2(new_n799_), .A3(KEYINPUT56), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n787_), .B1(new_n786_), .B2(KEYINPUT118), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n623_), .A2(new_n587_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n800_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n798_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n633_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n559_), .A2(KEYINPUT105), .A3(new_n554_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(KEYINPUT57), .A3(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n797_), .B1(new_n804_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT57), .ZN(new_n809_));
  NOR3_X1   g608(.A1(new_n632_), .A2(new_n633_), .A3(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n798_), .A2(new_n803_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n810_), .A2(KEYINPUT122), .A3(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n796_), .B1(new_n808_), .B2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n634_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT120), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT120), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n811_), .A2(new_n634_), .A3(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n815_), .A2(new_n809_), .A3(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n450_), .B1(new_n813_), .B2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n561_), .A2(new_n624_), .A3(new_n450_), .ZN(new_n820_));
  OAI21_X1  g619(.A(KEYINPUT54), .B1(new_n608_), .B2(new_n820_), .ZN(new_n821_));
  AOI211_X1 g620(.A(new_n623_), .B(new_n451_), .C1(new_n556_), .C2(new_n560_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n822_), .A2(new_n823_), .A3(new_n607_), .A4(new_n606_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n821_), .A2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n772_), .B1(new_n819_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(G113gat), .B1(new_n827_), .B2(new_n623_), .ZN(new_n828_));
  OR2_X1    g627(.A1(new_n828_), .A2(KEYINPUT123), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(KEYINPUT123), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n808_), .A2(new_n812_), .ZN(new_n831_));
  OR3_X1    g630(.A1(new_n794_), .A2(new_n561_), .A3(new_n795_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n818_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n825_), .B1(new_n833_), .B2(new_n451_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n772_), .ZN(new_n835_));
  OR2_X1    g634(.A1(new_n835_), .A2(KEYINPUT124), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT59), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(KEYINPUT124), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n836_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(KEYINPUT125), .B1(new_n834_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n839_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT125), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n841_), .B(new_n842_), .C1(new_n819_), .C2(new_n825_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n840_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n826_), .A2(KEYINPUT59), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n623_), .A2(G113gat), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(KEYINPUT126), .ZN(new_n848_));
  AOI22_X1  g647(.A1(new_n829_), .A2(new_n830_), .B1(new_n846_), .B2(new_n848_), .ZN(G1340gat));
  INV_X1    g648(.A(new_n608_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n850_), .B1(new_n826_), .B2(KEYINPUT59), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n815_), .A2(new_n809_), .A3(new_n817_), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n810_), .A2(KEYINPUT122), .A3(new_n811_), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT122), .B1(new_n810_), .B2(new_n811_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n832_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n451_), .B1(new_n852_), .B2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n825_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n842_), .B1(new_n858_), .B2(new_n841_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n843_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n851_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(G120gat), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n850_), .A2(KEYINPUT60), .ZN(new_n863_));
  INV_X1    g662(.A(G120gat), .ZN(new_n864_));
  MUX2_X1   g663(.A(KEYINPUT60), .B(new_n863_), .S(new_n864_), .Z(new_n865_));
  NAND2_X1  g664(.A1(new_n827_), .A2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n862_), .A2(KEYINPUT127), .A3(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT127), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n864_), .B1(new_n844_), .B2(new_n851_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n866_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n868_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n867_), .A2(new_n871_), .ZN(G1341gat));
  NAND3_X1  g671(.A1(new_n844_), .A2(new_n450_), .A3(new_n845_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(G127gat), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n451_), .A2(G127gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n826_), .B2(new_n875_), .ZN(G1342gat));
  NAND3_X1  g675(.A1(new_n844_), .A2(new_n562_), .A3(new_n845_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(G134gat), .ZN(new_n878_));
  OR2_X1    g677(.A1(new_n638_), .A2(G134gat), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n826_), .B2(new_n879_), .ZN(G1343gat));
  NOR4_X1   g679(.A1(new_n834_), .A2(new_n393_), .A3(new_n253_), .A4(new_n771_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n623_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n608_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g684(.A1(new_n881_), .A2(new_n450_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(KEYINPUT61), .B(G155gat), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n886_), .B(new_n887_), .ZN(G1346gat));
  NAND3_X1  g687(.A1(new_n881_), .A2(new_n316_), .A3(new_n637_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n881_), .A2(new_n562_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n889_), .B1(new_n891_), .B2(new_n316_), .ZN(G1347gat));
  NOR3_X1   g691(.A1(new_n410_), .A2(new_n628_), .A3(new_n415_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n858_), .A2(new_n623_), .A3(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(G169gat), .B1(new_n894_), .B2(KEYINPUT62), .ZN(new_n895_));
  OAI21_X1  g694(.A(KEYINPUT62), .B1(new_n894_), .B2(KEYINPUT22), .ZN(new_n896_));
  MUX2_X1   g695(.A(G169gat), .B(new_n895_), .S(new_n896_), .Z(G1348gat));
  AND2_X1   g696(.A1(new_n858_), .A2(new_n893_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n608_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n450_), .ZN(new_n901_));
  MUX2_X1   g700(.A(new_n274_), .B(G183gat), .S(new_n901_), .Z(G1350gat));
  NAND3_X1  g701(.A1(new_n898_), .A2(new_n637_), .A3(new_n220_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n898_), .A2(new_n562_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n903_), .B1(new_n905_), .B2(new_n224_), .ZN(G1351gat));
  NAND3_X1  g705(.A1(new_n411_), .A2(new_n665_), .A3(new_n254_), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n834_), .A2(new_n410_), .A3(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(new_n623_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n608_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g711(.A1(new_n908_), .A2(new_n450_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n914_));
  AND2_X1   g713(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n913_), .A2(new_n914_), .A3(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n916_), .B1(new_n913_), .B2(new_n914_), .ZN(G1354gat));
  INV_X1    g716(.A(G218gat), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n908_), .A2(new_n918_), .A3(new_n637_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n908_), .A2(new_n562_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n919_), .B1(new_n921_), .B2(new_n918_), .ZN(G1355gat));
endmodule


