//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 0 0 0 0 1 0 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n774_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n867_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n909_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_;
  XNOR2_X1  g000(.A(KEYINPUT67), .B(G92gat), .ZN(new_n202_));
  INV_X1    g001(.A(G85gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n203_), .A2(KEYINPUT9), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n202_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  AND2_X1   g005(.A1(new_n206_), .A2(KEYINPUT6), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n206_), .A2(KEYINPUT6), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  XOR2_X1   g008(.A(G85gat), .B(G92gat), .Z(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT9), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n205_), .A2(new_n209_), .A3(new_n211_), .ZN(new_n212_));
  OR2_X1    g011(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n214_));
  NAND2_X1  g013(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  AND2_X1   g015(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT64), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(KEYINPUT65), .B(G106gat), .Z(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT66), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n220_), .A2(KEYINPUT66), .A3(new_n221_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n212_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  OR3_X1    g025(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n228_));
  OAI211_X1 g027(.A(new_n227_), .B(new_n228_), .C1(new_n207_), .C2(new_n208_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT8), .ZN(new_n230_));
  AND3_X1   g029(.A1(new_n229_), .A2(new_n230_), .A3(new_n210_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n230_), .B1(new_n229_), .B2(new_n210_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT69), .B1(new_n226_), .B2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G29gat), .B(G36gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G43gat), .B(G50gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT15), .ZN(new_n238_));
  AND3_X1   g037(.A1(new_n205_), .A2(new_n209_), .A3(new_n211_), .ZN(new_n239_));
  AND3_X1   g038(.A1(new_n220_), .A2(KEYINPUT66), .A3(new_n221_), .ZN(new_n240_));
  AOI21_X1  g039(.A(KEYINPUT66), .B1(new_n220_), .B2(new_n221_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n239_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT69), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n229_), .A2(new_n210_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT8), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n229_), .A2(new_n230_), .A3(new_n210_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n242_), .A2(new_n243_), .A3(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n234_), .A2(new_n238_), .A3(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT74), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT74), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n234_), .A2(new_n248_), .A3(new_n251_), .A4(new_n238_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n242_), .A2(new_n247_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT73), .B(KEYINPUT35), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G232gat), .A2(G233gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  AOI22_X1  g058(.A1(new_n255_), .A2(new_n237_), .B1(new_n256_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n253_), .A2(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n259_), .A2(new_n256_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n253_), .B(new_n260_), .C1(new_n256_), .C2(new_n259_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(KEYINPUT75), .A3(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G190gat), .B(G218gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G134gat), .B(G162gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n268_), .A2(KEYINPUT36), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n265_), .A2(new_n270_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n263_), .A2(KEYINPUT75), .A3(new_n264_), .A4(new_n269_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n268_), .A2(KEYINPUT36), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n274_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n273_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT37), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT37), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n273_), .A2(new_n279_), .A3(new_n276_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G15gat), .B(G22gat), .ZN(new_n282_));
  INV_X1    g081(.A(G1gat), .ZN(new_n283_));
  INV_X1    g082(.A(G8gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT14), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G1gat), .B(G8gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT76), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G231gat), .A2(G233gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT68), .B(G71gat), .ZN(new_n292_));
  INV_X1    g091(.A(G78gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G57gat), .B(G64gat), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n295_), .A2(KEYINPUT11), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n295_), .B(KEYINPUT11), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(new_n294_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n291_), .B(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(G127gat), .B(G155gat), .Z(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT16), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G183gat), .B(G211gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT17), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n306_), .A2(new_n307_), .ZN(new_n309_));
  OR3_X1    g108(.A1(new_n302_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n302_), .A2(new_n308_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n312_), .B(KEYINPUT77), .Z(new_n313_));
  NOR2_X1   g112(.A1(new_n281_), .A2(new_n313_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n234_), .A2(KEYINPUT12), .A3(new_n248_), .A4(new_n300_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n254_), .A2(new_n300_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n254_), .A2(new_n300_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  XOR2_X1   g118(.A(KEYINPUT70), .B(KEYINPUT12), .Z(new_n320_));
  OAI211_X1 g119(.A(new_n315_), .B(new_n317_), .C1(new_n319_), .C2(new_n320_), .ZN(new_n321_));
  AND2_X1   g120(.A1(G230gat), .A2(G233gat), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n322_), .B1(new_n319_), .B2(new_n316_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G120gat), .B(G148gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT5), .ZN(new_n327_));
  XOR2_X1   g126(.A(G176gat), .B(G204gat), .Z(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  OR2_X1    g128(.A1(new_n325_), .A2(new_n329_), .ZN(new_n330_));
  XOR2_X1   g129(.A(new_n329_), .B(KEYINPUT71), .Z(new_n331_));
  NAND2_X1  g130(.A1(new_n325_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n333_), .A2(KEYINPUT13), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(KEYINPUT13), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n314_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT88), .ZN(new_n338_));
  INV_X1    g137(.A(G204gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT89), .ZN(new_n341_));
  NAND2_X1  g140(.A1(KEYINPUT88), .A2(G204gat), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n340_), .A2(new_n341_), .A3(G197gat), .A4(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT21), .ZN(new_n344_));
  INV_X1    g143(.A(G218gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(G211gat), .ZN(new_n346_));
  INV_X1    g145(.A(G211gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(G218gat), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n344_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n349_));
  AND2_X1   g148(.A1(KEYINPUT88), .A2(G204gat), .ZN(new_n350_));
  NOR2_X1   g149(.A1(KEYINPUT88), .A2(G204gat), .ZN(new_n351_));
  INV_X1    g150(.A(G197gat), .ZN(new_n352_));
  NOR3_X1   g151(.A1(new_n350_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT89), .B1(new_n339_), .B2(G197gat), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n343_), .B(new_n349_), .C1(new_n353_), .C2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT91), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n340_), .A2(G197gat), .A3(new_n342_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n354_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n360_), .A2(KEYINPUT91), .A3(new_n343_), .A4(new_n349_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n357_), .A2(new_n361_), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n350_), .A2(new_n351_), .A3(G197gat), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n344_), .B1(G197gat), .B2(G204gat), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n346_), .B(new_n348_), .C1(new_n363_), .C2(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n350_), .A2(new_n351_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n354_), .B1(new_n367_), .B2(G197gat), .ZN(new_n368_));
  INV_X1    g167(.A(new_n343_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n344_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n366_), .B1(new_n370_), .B2(KEYINPUT90), .ZN(new_n371_));
  AOI21_X1  g170(.A(KEYINPUT21), .B1(new_n360_), .B2(new_n343_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT90), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n362_), .B1(new_n371_), .B2(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(G169gat), .A2(G176gat), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT24), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G183gat), .A2(G190gat), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT23), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n378_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  OR2_X1    g182(.A1(new_n383_), .A2(KEYINPUT81), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(KEYINPUT81), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT25), .B(G183gat), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT26), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT80), .B1(new_n387_), .B2(G190gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT26), .B(G190gat), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n386_), .B(new_n388_), .C1(new_n389_), .C2(KEYINPUT80), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G169gat), .A2(G176gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT24), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n376_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n385_), .A2(new_n390_), .A3(new_n395_), .ZN(new_n396_));
  OR2_X1    g195(.A1(G183gat), .A2(G190gat), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT85), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n381_), .A2(new_n397_), .A3(new_n398_), .A4(new_n382_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n391_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n379_), .A2(KEYINPUT23), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n380_), .A2(G183gat), .A3(G190gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(new_n397_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n400_), .B1(new_n404_), .B2(KEYINPUT85), .ZN(new_n405_));
  AND2_X1   g204(.A1(KEYINPUT82), .A2(KEYINPUT22), .ZN(new_n406_));
  NOR2_X1   g205(.A1(KEYINPUT82), .A2(KEYINPUT22), .ZN(new_n407_));
  OAI21_X1  g206(.A(G169gat), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT83), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  OAI211_X1 g209(.A(KEYINPUT83), .B(G169gat), .C1(new_n406_), .C2(new_n407_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT84), .B(G176gat), .ZN(new_n413_));
  INV_X1    g212(.A(G169gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT22), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n412_), .A2(new_n416_), .ZN(new_n417_));
  AOI22_X1  g216(.A1(new_n384_), .A2(new_n396_), .B1(new_n405_), .B2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT20), .B1(new_n375_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n370_), .A2(KEYINPUT90), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n346_), .A2(new_n348_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n363_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n421_), .B1(new_n422_), .B2(new_n364_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n420_), .A2(new_n374_), .A3(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n362_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n383_), .B1(new_n389_), .B2(new_n386_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n376_), .B1(new_n392_), .B2(KEYINPUT96), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n427_), .B1(KEYINPUT96), .B2(new_n392_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT22), .B(G169gat), .ZN(new_n429_));
  AOI22_X1  g228(.A1(new_n413_), .A2(new_n429_), .B1(G169gat), .B2(G176gat), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n426_), .A2(new_n428_), .B1(new_n404_), .B2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n424_), .A2(new_n425_), .A3(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G226gat), .A2(G233gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n432_), .A2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT97), .B1(new_n419_), .B2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT20), .B1(new_n375_), .B2(new_n431_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n423_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n440_));
  AOI211_X1 g239(.A(KEYINPUT90), .B(KEYINPUT21), .C1(new_n360_), .C2(new_n343_), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n357_), .B(new_n361_), .C1(new_n440_), .C2(new_n441_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n384_), .A2(new_n385_), .A3(new_n395_), .A4(new_n390_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n412_), .A2(new_n416_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n404_), .A2(KEYINPUT85), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(new_n391_), .A3(new_n399_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n443_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n442_), .A2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n435_), .B1(new_n439_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT20), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n450_), .B1(new_n442_), .B2(new_n447_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT97), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n451_), .A2(new_n452_), .A3(new_n436_), .A4(new_n432_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n438_), .A2(new_n449_), .A3(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G8gat), .B(G36gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT18), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G64gat), .B(G92gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n454_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n458_), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n438_), .A2(new_n449_), .A3(new_n453_), .A4(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT27), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G127gat), .B(G134gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G113gat), .B(G120gat), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT87), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n465_), .A2(new_n466_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n467_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n465_), .A2(new_n466_), .A3(KEYINPUT87), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT2), .ZN(new_n472_));
  INV_X1    g271(.A(G141gat), .ZN(new_n473_));
  INV_X1    g272(.A(G148gat), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n472_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT3), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n476_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n475_), .A2(new_n477_), .A3(new_n478_), .A4(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G155gat), .A2(G162gat), .ZN(new_n481_));
  OR2_X1    g280(.A1(G155gat), .A2(G162gat), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n480_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  XOR2_X1   g282(.A(G141gat), .B(G148gat), .Z(new_n484_));
  NAND2_X1  g283(.A1(new_n481_), .A2(KEYINPUT1), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n482_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n481_), .A2(KEYINPUT1), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n484_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n470_), .A2(new_n471_), .B1(new_n483_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n467_), .A2(new_n469_), .ZN(new_n490_));
  AND3_X1   g289(.A1(new_n490_), .A2(new_n488_), .A3(new_n483_), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT4), .B1(new_n489_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G225gat), .A2(G233gat), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n470_), .A2(new_n471_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n483_), .A2(new_n488_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT4), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n492_), .A2(new_n494_), .A3(new_n499_), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n489_), .A2(new_n491_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n493_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G1gat), .B(G29gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(G85gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(KEYINPUT0), .B(G57gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n503_), .A2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n500_), .A2(new_n502_), .A3(new_n507_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G22gat), .B(G50gat), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n483_), .A2(new_n488_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT29), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n516_), .A2(KEYINPUT28), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n496_), .A2(KEYINPUT29), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT28), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n513_), .B1(new_n517_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n516_), .A2(KEYINPUT28), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n518_), .A2(new_n519_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(new_n523_), .A3(new_n512_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n521_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G228gat), .A2(G233gat), .ZN(new_n526_));
  XOR2_X1   g325(.A(new_n526_), .B(KEYINPUT92), .Z(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n515_), .B1(new_n483_), .B2(new_n488_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n528_), .B1(new_n375_), .B2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G78gat), .B(G106gat), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n529_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n526_), .A2(KEYINPUT92), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n442_), .A2(new_n533_), .A3(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n530_), .A2(new_n532_), .A3(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n525_), .B1(new_n537_), .B2(KEYINPUT94), .ZN(new_n538_));
  AOI211_X1 g337(.A(new_n529_), .B(new_n534_), .C1(new_n424_), .C2(new_n425_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n527_), .B1(new_n442_), .B2(new_n533_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n531_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT93), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT93), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n543_), .B(new_n531_), .C1(new_n539_), .C2(new_n540_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT94), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n530_), .A2(new_n545_), .A3(new_n536_), .A4(new_n532_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n538_), .A2(new_n542_), .A3(new_n544_), .A4(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n541_), .A2(new_n537_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(new_n525_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n511_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n550_));
  NOR3_X1   g349(.A1(new_n439_), .A2(new_n448_), .A3(new_n435_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n436_), .B1(new_n451_), .B2(new_n432_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n458_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT99), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n432_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n435_), .B1(new_n419_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n431_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n450_), .B1(new_n442_), .B2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n375_), .A2(new_n418_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n559_), .A2(new_n436_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n557_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n562_), .A2(KEYINPUT99), .A3(new_n458_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n555_), .A2(KEYINPUT27), .A3(new_n461_), .A4(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n464_), .A2(new_n550_), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT100), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n464_), .A2(new_n550_), .A3(new_n564_), .A4(KEYINPUT100), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n460_), .A2(KEYINPUT32), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n570_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n438_), .A2(new_n449_), .A3(new_n453_), .A4(new_n569_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n571_), .A2(new_n572_), .A3(new_n511_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(KEYINPUT98), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n503_), .A2(KEYINPUT33), .A3(new_n508_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n507_), .B1(new_n501_), .B2(new_n493_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n494_), .B1(new_n492_), .B2(new_n499_), .ZN(new_n577_));
  OAI21_X1  g376(.A(KEYINPUT33), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n509_), .A2(new_n578_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n459_), .A2(new_n461_), .A3(new_n575_), .A4(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT98), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n572_), .A2(new_n571_), .A3(new_n511_), .A4(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n574_), .A2(new_n580_), .A3(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n547_), .A2(new_n549_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n567_), .A2(new_n568_), .A3(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT30), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n447_), .B(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT86), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G71gat), .B(G99gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(G43gat), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G227gat), .A2(G233gat), .ZN(new_n593_));
  INV_X1    g392(.A(G15gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n592_), .B(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n590_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n589_), .A2(KEYINPUT86), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(new_n596_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n495_), .B(KEYINPUT31), .Z(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n598_), .A2(new_n600_), .A3(new_n602_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n587_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n461_), .A2(KEYINPUT27), .ZN(new_n608_));
  AOI21_X1  g407(.A(KEYINPUT99), .B1(new_n562_), .B2(new_n458_), .ZN(new_n609_));
  AOI211_X1 g408(.A(new_n554_), .B(new_n460_), .C1(new_n557_), .C2(new_n561_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n608_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(KEYINPUT27), .B1(new_n459_), .B2(new_n461_), .ZN(new_n612_));
  OAI21_X1  g411(.A(KEYINPUT101), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT101), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n464_), .A2(new_n614_), .A3(new_n564_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n584_), .B1(new_n613_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n511_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n604_), .A2(new_n605_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n616_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n607_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n238_), .A2(new_n288_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n288_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(new_n237_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(G229gat), .A2(G233gat), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n625_), .A2(KEYINPUT78), .A3(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n288_), .B(new_n237_), .Z(new_n629_));
  AOI21_X1  g428(.A(new_n628_), .B1(new_n627_), .B2(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT78), .B1(new_n625_), .B2(new_n627_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G113gat), .B(G141gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(G169gat), .B(G197gat), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n633_), .B(new_n634_), .Z(new_n635_));
  NAND2_X1  g434(.A1(new_n632_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT79), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n632_), .A2(new_n635_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n621_), .A2(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n337_), .A2(new_n641_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT102), .Z(new_n643_));
  OR2_X1    g442(.A1(new_n617_), .A2(KEYINPUT103), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n617_), .A2(KEYINPUT103), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n643_), .A2(new_n283_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT38), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  XOR2_X1   g449(.A(new_n650_), .B(KEYINPUT105), .Z(new_n651_));
  AOI22_X1  g450(.A1(new_n587_), .A2(new_n606_), .B1(new_n616_), .B2(new_n619_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT104), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n277_), .A2(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n273_), .A2(KEYINPUT104), .A3(new_n276_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n652_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n336_), .A2(new_n640_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n312_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n657_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G1gat), .B1(new_n661_), .B2(new_n617_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n651_), .B(new_n662_), .C1(new_n649_), .C2(new_n648_), .ZN(G1324gat));
  NAND2_X1  g462(.A1(new_n613_), .A2(new_n615_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n643_), .A2(new_n284_), .A3(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(G8gat), .B1(new_n661_), .B2(new_n664_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT39), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(G1325gat));
  OAI21_X1  g470(.A(G15gat), .B1(new_n661_), .B2(new_n606_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT41), .Z(new_n673_));
  INV_X1    g472(.A(new_n606_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n642_), .A2(new_n594_), .A3(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(G1326gat));
  OAI21_X1  g475(.A(G22gat), .B1(new_n661_), .B2(new_n585_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT42), .ZN(new_n678_));
  INV_X1    g477(.A(G22gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n642_), .A2(new_n679_), .A3(new_n584_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(G1327gat));
  INV_X1    g480(.A(new_n656_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n313_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n336_), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n685_), .A2(new_n641_), .A3(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(G29gat), .B1(new_n687_), .B2(new_n511_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n279_), .B1(new_n273_), .B2(new_n276_), .ZN(new_n689_));
  AOI211_X1 g488(.A(KEYINPUT37), .B(new_n275_), .C1(new_n271_), .C2(new_n272_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  OAI211_X1 g490(.A(KEYINPUT107), .B(KEYINPUT43), .C1(new_n652_), .C2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AOI22_X1  g492(.A1(new_n565_), .A2(new_n566_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n674_), .B1(new_n694_), .B2(new_n568_), .ZN(new_n695_));
  AOI211_X1 g494(.A(new_n584_), .B(new_n618_), .C1(new_n613_), .C2(new_n615_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n281_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT107), .B1(new_n697_), .B2(KEYINPUT43), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n691_), .B1(new_n607_), .B2(new_n620_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n700_));
  AOI21_X1  g499(.A(KEYINPUT108), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT108), .ZN(new_n702_));
  NOR4_X1   g501(.A1(new_n652_), .A2(new_n702_), .A3(KEYINPUT43), .A4(new_n691_), .ZN(new_n703_));
  OAI22_X1  g502(.A1(new_n693_), .A2(new_n698_), .B1(new_n701_), .B2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n704_), .A2(new_n313_), .A3(new_n659_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n706_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n647_), .A2(G29gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n688_), .B1(new_n709_), .B2(new_n710_), .ZN(G1328gat));
  NAND3_X1  g510(.A1(new_n707_), .A2(new_n665_), .A3(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(G36gat), .ZN(new_n713_));
  INV_X1    g512(.A(new_n687_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n714_), .A2(G36gat), .A3(new_n664_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT45), .Z(new_n716_));
  NAND2_X1  g515(.A1(new_n713_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT46), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n717_), .B(new_n718_), .ZN(G1329gat));
  NAND3_X1  g518(.A1(new_n709_), .A2(G43gat), .A3(new_n674_), .ZN(new_n720_));
  INV_X1    g519(.A(G43gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n721_), .B1(new_n714_), .B2(new_n606_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT47), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT47), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n720_), .A2(new_n725_), .A3(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1330gat));
  AOI21_X1  g526(.A(G50gat), .B1(new_n687_), .B2(new_n584_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n584_), .A2(G50gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n709_), .B2(new_n729_), .ZN(G1331gat));
  NOR2_X1   g529(.A1(new_n336_), .A2(new_n640_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n621_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(new_n314_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(G57gat), .B1(new_n735_), .B2(new_n647_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n640_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n657_), .A2(new_n737_), .A3(new_n683_), .A4(new_n686_), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT109), .Z(new_n739_));
  XNOR2_X1  g538(.A(KEYINPUT110), .B(G57gat), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n617_), .A2(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n736_), .B1(new_n739_), .B2(new_n741_), .ZN(G1332gat));
  INV_X1    g541(.A(G64gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n739_), .B2(new_n665_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT48), .Z(new_n745_));
  NAND3_X1  g544(.A1(new_n735_), .A2(new_n743_), .A3(new_n665_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1333gat));
  INV_X1    g546(.A(G71gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n739_), .B2(new_n674_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(KEYINPUT111), .B(KEYINPUT49), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n749_), .B(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n735_), .A2(new_n748_), .A3(new_n674_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1334gat));
  AOI21_X1  g552(.A(new_n293_), .B1(new_n739_), .B2(new_n584_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n754_), .B(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n584_), .A2(new_n293_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT113), .Z(new_n758_));
  OAI21_X1  g557(.A(new_n756_), .B1(new_n734_), .B2(new_n758_), .ZN(G1335gat));
  NOR2_X1   g558(.A1(new_n685_), .A2(new_n732_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n760_), .A2(new_n203_), .A3(new_n647_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT107), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n762_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n700_), .B(new_n281_), .C1(new_n695_), .C2(new_n696_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n702_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n621_), .A2(KEYINPUT108), .A3(new_n700_), .A4(new_n281_), .ZN(new_n766_));
  AOI22_X1  g565(.A1(new_n763_), .A2(new_n692_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT114), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n686_), .A2(new_n737_), .A3(new_n313_), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n768_), .A2(new_n617_), .A3(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n761_), .B1(new_n770_), .B2(new_n203_), .ZN(G1336gat));
  AOI21_X1  g570(.A(G92gat), .B1(new_n760_), .B2(new_n665_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n768_), .A2(new_n769_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n664_), .A2(new_n202_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n772_), .B1(new_n773_), .B2(new_n774_), .ZN(G1337gat));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n674_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n606_), .B1(new_n216_), .B2(new_n219_), .ZN(new_n777_));
  AOI22_X1  g576(.A1(new_n776_), .A2(G99gat), .B1(new_n760_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n778_), .B(new_n779_), .ZN(G1338gat));
  NAND3_X1  g579(.A1(new_n760_), .A2(new_n584_), .A3(new_n221_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n769_), .A2(new_n585_), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT115), .B1(new_n704_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT115), .ZN(new_n785_));
  INV_X1    g584(.A(new_n783_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n767_), .A2(new_n785_), .A3(new_n786_), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n782_), .B(G106gat), .C1(new_n784_), .C2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT116), .ZN(new_n789_));
  OAI21_X1  g588(.A(G106gat), .B1(new_n784_), .B2(new_n787_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(new_n791_), .A3(KEYINPUT52), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n789_), .A2(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n785_), .B1(new_n767_), .B2(new_n786_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n704_), .A2(KEYINPUT115), .A3(new_n783_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n796_), .A2(new_n797_), .A3(new_n782_), .A4(G106gat), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n782_), .B1(new_n796_), .B2(G106gat), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(new_n791_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n781_), .B1(new_n793_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT53), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n803_), .B(new_n781_), .C1(new_n793_), .C2(new_n800_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(G1339gat));
  INV_X1    g604(.A(KEYINPUT57), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT120), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n626_), .B1(new_n625_), .B2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n808_), .B1(new_n807_), .B2(new_n625_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n635_), .B1(new_n629_), .B2(new_n626_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n638_), .A2(new_n811_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n812_), .A2(new_n333_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n330_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n321_), .A2(new_n322_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n323_), .A2(KEYINPUT55), .A3(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT119), .ZN(new_n817_));
  OR3_X1    g616(.A1(new_n321_), .A2(KEYINPUT55), .A3(new_n322_), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n816_), .A2(new_n817_), .A3(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n817_), .B1(new_n816_), .B2(new_n818_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n331_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT56), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  OAI211_X1 g622(.A(KEYINPUT56), .B(new_n331_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n814_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n813_), .B1(new_n825_), .B2(new_n640_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n806_), .B1(new_n826_), .B2(new_n656_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n825_), .A2(new_n640_), .ZN(new_n828_));
  OAI211_X1 g627(.A(KEYINPUT57), .B(new_n682_), .C1(new_n828_), .C2(new_n813_), .ZN(new_n829_));
  AOI21_X1  g628(.A(KEYINPUT58), .B1(new_n825_), .B2(new_n812_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n825_), .A2(KEYINPUT58), .A3(new_n812_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n281_), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n827_), .B(new_n829_), .C1(new_n830_), .C2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n312_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n835_), .B1(new_n337_), .B2(new_n640_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(KEYINPUT118), .A2(KEYINPUT54), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n314_), .A2(new_n737_), .A3(new_n336_), .A4(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n834_), .A2(new_n839_), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n616_), .A2(new_n674_), .A3(new_n647_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(G113gat), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n842_), .A2(new_n843_), .A3(new_n640_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n840_), .A2(KEYINPUT59), .A3(new_n841_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT59), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n833_), .A2(new_n313_), .B1(new_n836_), .B2(new_n838_), .ZN(new_n847_));
  XOR2_X1   g646(.A(new_n841_), .B(KEYINPUT121), .Z(new_n848_));
  OAI21_X1  g647(.A(new_n846_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n737_), .B1(new_n845_), .B2(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n844_), .B1(new_n850_), .B2(new_n843_), .ZN(G1340gat));
  INV_X1    g650(.A(G120gat), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n852_), .B1(new_n336_), .B2(KEYINPUT60), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n852_), .A2(KEYINPUT60), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(KEYINPUT122), .B2(new_n854_), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n842_), .B(new_n855_), .C1(KEYINPUT122), .C2(new_n853_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n336_), .B1(new_n845_), .B2(new_n849_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n857_), .A2(KEYINPUT123), .ZN(new_n858_));
  OAI21_X1  g657(.A(G120gat), .B1(new_n857_), .B2(KEYINPUT123), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n856_), .B1(new_n858_), .B2(new_n859_), .ZN(G1341gat));
  INV_X1    g659(.A(G127gat), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n842_), .A2(new_n861_), .A3(new_n683_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n312_), .B1(new_n845_), .B2(new_n849_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n863_), .B2(new_n861_), .ZN(G1342gat));
  INV_X1    g663(.A(G134gat), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n842_), .A2(new_n865_), .A3(new_n656_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n691_), .B1(new_n845_), .B2(new_n849_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(new_n865_), .ZN(G1343gat));
  NOR3_X1   g667(.A1(new_n674_), .A2(new_n585_), .A3(new_n646_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n840_), .A2(new_n664_), .A3(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n870_), .A2(new_n737_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(new_n473_), .ZN(G1344gat));
  NOR2_X1   g671(.A1(new_n870_), .A2(new_n336_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(new_n474_), .ZN(G1345gat));
  NOR2_X1   g673(.A1(new_n870_), .A2(new_n313_), .ZN(new_n875_));
  XOR2_X1   g674(.A(KEYINPUT61), .B(G155gat), .Z(new_n876_));
  XNOR2_X1  g675(.A(new_n875_), .B(new_n876_), .ZN(G1346gat));
  OAI21_X1  g676(.A(G162gat), .B1(new_n870_), .B2(new_n691_), .ZN(new_n878_));
  OR2_X1    g677(.A1(new_n682_), .A2(G162gat), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n870_), .B2(new_n879_), .ZN(G1347gat));
  NAND2_X1  g679(.A1(new_n833_), .A2(new_n313_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n839_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n665_), .A2(new_n674_), .A3(new_n646_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(KEYINPUT124), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n584_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n882_), .A2(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(KEYINPUT125), .B1(new_n886_), .B2(new_n737_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n885_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n847_), .A2(new_n737_), .A3(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT125), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n887_), .A2(new_n891_), .A3(G169gat), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n889_), .A2(new_n429_), .ZN(new_n895_));
  NAND4_X1  g694(.A1(new_n887_), .A2(new_n891_), .A3(KEYINPUT62), .A4(G169gat), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n894_), .A2(new_n895_), .A3(new_n896_), .ZN(G1348gat));
  INV_X1    g696(.A(new_n886_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n686_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n584_), .B1(new_n834_), .B2(new_n839_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n884_), .ZN(new_n901_));
  AND3_X1   g700(.A1(new_n901_), .A2(G176gat), .A3(new_n686_), .ZN(new_n902_));
  AOI22_X1  g701(.A1(new_n899_), .A2(new_n413_), .B1(new_n900_), .B2(new_n902_), .ZN(G1349gat));
  NOR3_X1   g702(.A1(new_n886_), .A2(new_n386_), .A3(new_n312_), .ZN(new_n904_));
  INV_X1    g703(.A(G183gat), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n900_), .A2(new_n683_), .A3(new_n901_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n904_), .B1(new_n905_), .B2(new_n906_), .ZN(G1350gat));
  OAI21_X1  g706(.A(G190gat), .B1(new_n886_), .B2(new_n691_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n656_), .A2(new_n389_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n886_), .B2(new_n909_), .ZN(G1351gat));
  NAND2_X1  g709(.A1(new_n606_), .A2(new_n550_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(KEYINPUT126), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n912_), .A2(new_n664_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n840_), .A2(new_n913_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n914_), .A2(new_n737_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(new_n352_), .ZN(G1352gat));
  INV_X1    g715(.A(KEYINPUT127), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n914_), .A2(new_n336_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n918_), .B2(new_n339_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n367_), .ZN(new_n920_));
  OAI211_X1 g719(.A(KEYINPUT127), .B(G204gat), .C1(new_n914_), .C2(new_n336_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n919_), .A2(new_n920_), .A3(new_n921_), .ZN(G1353gat));
  NOR2_X1   g721(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n923_));
  AND2_X1   g722(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n924_));
  NOR4_X1   g723(.A1(new_n914_), .A2(new_n312_), .A3(new_n923_), .A4(new_n924_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n914_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(new_n660_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n925_), .B1(new_n927_), .B2(new_n923_), .ZN(G1354gat));
  OAI21_X1  g727(.A(G218gat), .B1(new_n914_), .B2(new_n691_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n656_), .A2(new_n345_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n914_), .B2(new_n930_), .ZN(G1355gat));
endmodule


