//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0 1 1 1 0 0 0 1 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n637_, new_n638_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n869_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n909_, new_n910_, new_n911_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G57gat), .B(G64gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G71gat), .B(G78gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n204_), .A2(new_n205_), .A3(KEYINPUT11), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(KEYINPUT11), .ZN(new_n207_));
  INV_X1    g006(.A(new_n205_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n204_), .A2(KEYINPUT11), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n206_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT67), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n213_), .B(new_n206_), .C1(new_n209_), .C2(new_n210_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT6), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT6), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(G99gat), .A3(G106gat), .ZN(new_n219_));
  AND3_X1   g018(.A1(new_n217_), .A2(new_n219_), .A3(KEYINPUT65), .ZN(new_n220_));
  AOI21_X1  g019(.A(KEYINPUT65), .B1(new_n217_), .B2(new_n219_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT9), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n224_), .A2(G85gat), .A3(G92gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G85gat), .B(G92gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT10), .B(G99gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT64), .B(G106gat), .ZN(new_n228_));
  OAI221_X1 g027(.A(new_n225_), .B1(new_n226_), .B2(new_n224_), .C1(new_n227_), .C2(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n223_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n217_), .A2(new_n219_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT7), .ZN(new_n235_));
  INV_X1    g034(.A(G99gat), .ZN(new_n236_));
  INV_X1    g035(.A(G106gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n217_), .A2(new_n219_), .A3(KEYINPUT65), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n234_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n226_), .A2(KEYINPUT8), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n246_));
  AOI22_X1  g045(.A1(new_n240_), .A2(new_n246_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n238_), .A2(KEYINPUT66), .A3(new_n239_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n226_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT8), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n245_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n215_), .A2(new_n231_), .A3(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n215_), .B1(new_n251_), .B2(new_n231_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n203_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT12), .ZN(new_n256_));
  OR2_X1    g055(.A1(new_n211_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n239_), .ZN(new_n259_));
  NOR3_X1   g058(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n246_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(new_n232_), .A3(new_n248_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n226_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n250_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n244_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n265_), .B1(new_n222_), .B2(new_n241_), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT68), .B1(new_n264_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n245_), .B(new_n268_), .C1(new_n249_), .C2(new_n250_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(KEYINPUT69), .B1(new_n270_), .B2(new_n231_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n272_));
  AOI211_X1 g071(.A(new_n272_), .B(new_n230_), .C1(new_n267_), .C2(new_n269_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n258_), .B1(new_n271_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n254_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n275_), .B1(new_n253_), .B2(new_n256_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n255_), .B1(new_n277_), .B2(new_n203_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G120gat), .B(G148gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT5), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G176gat), .B(G204gat), .ZN(new_n281_));
  XOR2_X1   g080(.A(new_n280_), .B(new_n281_), .Z(new_n282_));
  NAND2_X1  g081(.A1(new_n278_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n282_), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n255_), .B(new_n284_), .C1(new_n277_), .C2(new_n203_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n286_), .B1(KEYINPUT70), .B2(KEYINPUT13), .ZN(new_n287_));
  AND2_X1   g086(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n288_));
  NOR2_X1   g087(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n283_), .B(new_n285_), .C1(new_n288_), .C2(new_n289_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n287_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n292_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G127gat), .B(G155gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT16), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G183gat), .B(G211gat), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n297_), .A2(new_n298_), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT17), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(G1gat), .ZN(new_n302_));
  INV_X1    g101(.A(G8gat), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT14), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT73), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  OAI211_X1 g105(.A(KEYINPUT73), .B(KEYINPUT14), .C1(new_n302_), .C2(new_n303_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G15gat), .B(G22gat), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n306_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(G1gat), .B(G8gat), .Z(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n306_), .A2(new_n310_), .A3(new_n307_), .A4(new_n308_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(G231gat), .ZN(new_n315_));
  INV_X1    g114(.A(G233gat), .ZN(new_n316_));
  NOR3_X1   g115(.A1(new_n314_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n315_), .A2(new_n316_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n318_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n211_), .B(KEYINPUT74), .Z(new_n322_));
  AOI21_X1  g121(.A(new_n301_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n323_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n215_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n320_), .B(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n301_), .ZN(new_n327_));
  NOR3_X1   g126(.A1(new_n299_), .A2(new_n300_), .A3(KEYINPUT17), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n326_), .A2(KEYINPUT75), .A3(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(KEYINPUT75), .B1(new_n326_), .B2(new_n329_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n324_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT76), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT76), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n334_), .B(new_n324_), .C1(new_n330_), .C2(new_n331_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G232gat), .A2(G233gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT34), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT35), .ZN(new_n339_));
  XOR2_X1   g138(.A(G29gat), .B(G36gat), .Z(new_n340_));
  XOR2_X1   g139(.A(G43gat), .B(G50gat), .Z(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT15), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n343_), .B1(new_n271_), .B2(new_n273_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n339_), .B1(new_n344_), .B2(KEYINPUT72), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n231_), .A2(new_n251_), .A3(new_n342_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n338_), .A2(KEYINPUT35), .ZN(new_n348_));
  OR3_X1    g147(.A1(new_n345_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT36), .ZN(new_n350_));
  XOR2_X1   g149(.A(G134gat), .B(G162gat), .Z(new_n351_));
  XNOR2_X1  g150(.A(G190gat), .B(G218gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n345_), .A2(new_n347_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n349_), .A2(new_n350_), .A3(new_n353_), .A4(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n353_), .A2(new_n350_), .ZN(new_n356_));
  OR2_X1    g155(.A1(new_n353_), .A2(new_n350_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n354_), .ZN(new_n358_));
  NOR3_X1   g157(.A1(new_n345_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n356_), .B(new_n357_), .C1(new_n358_), .C2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n355_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT37), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n355_), .A2(new_n360_), .A3(KEYINPUT37), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NOR3_X1   g164(.A1(new_n295_), .A2(new_n336_), .A3(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(G169gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G183gat), .A2(G190gat), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n370_), .A2(KEYINPUT23), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n369_), .B(KEYINPUT83), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n371_), .B1(new_n372_), .B2(KEYINPUT23), .ZN(new_n373_));
  INV_X1    g172(.A(G183gat), .ZN(new_n374_));
  OR2_X1    g173(.A1(new_n374_), .A2(KEYINPUT79), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(KEYINPUT79), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n373_), .B1(G190gat), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT23), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n370_), .A2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n380_), .B1(new_n372_), .B2(new_n379_), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(G169gat), .ZN(new_n384_));
  INV_X1    g183(.A(G176gat), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n383_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  OR3_X1    g185(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n381_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT80), .ZN(new_n390_));
  OAI211_X1 g189(.A(KEYINPUT25), .B(new_n376_), .C1(new_n375_), .C2(new_n390_), .ZN(new_n391_));
  AND2_X1   g190(.A1(KEYINPUT81), .A2(KEYINPUT26), .ZN(new_n392_));
  NOR2_X1   g191(.A1(KEYINPUT81), .A2(KEYINPUT26), .ZN(new_n393_));
  OAI21_X1  g192(.A(G190gat), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT82), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT82), .ZN(new_n396_));
  OAI211_X1 g195(.A(new_n396_), .B(G190gat), .C1(new_n392_), .C2(new_n393_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n374_), .A2(KEYINPUT25), .ZN(new_n398_));
  INV_X1    g197(.A(G190gat), .ZN(new_n399_));
  AOI22_X1  g198(.A1(new_n398_), .A2(KEYINPUT80), .B1(KEYINPUT26), .B2(new_n399_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n391_), .A2(new_n395_), .A3(new_n397_), .A4(new_n400_), .ZN(new_n401_));
  AOI22_X1  g200(.A1(new_n368_), .A2(new_n378_), .B1(new_n389_), .B2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT84), .B(G15gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G227gat), .A2(G233gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n402_), .B(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(G127gat), .B(G134gat), .Z(new_n407_));
  XOR2_X1   g206(.A(G113gat), .B(G120gat), .Z(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n406_), .B(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G71gat), .B(G99gat), .ZN(new_n412_));
  INV_X1    g211(.A(G43gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT30), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT31), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n411_), .B(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT85), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G226gat), .A2(G233gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT19), .ZN(new_n420_));
  XOR2_X1   g219(.A(G197gat), .B(G204gat), .Z(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT21), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G197gat), .B(G204gat), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT21), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G211gat), .B(G218gat), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n422_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  OR3_X1    g226(.A1(new_n423_), .A2(new_n426_), .A3(new_n424_), .ZN(new_n428_));
  AND3_X1   g227(.A1(new_n427_), .A2(KEYINPUT90), .A3(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(KEYINPUT90), .B1(new_n427_), .B2(new_n428_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n378_), .A2(new_n368_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n389_), .A2(new_n401_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT20), .B1(new_n431_), .B2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n427_), .A2(new_n428_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT26), .B(G190gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(KEYINPUT25), .B(G183gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(new_n386_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT94), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n441_), .A2(KEYINPUT94), .ZN(new_n444_));
  OAI211_X1 g243(.A(new_n373_), .B(new_n387_), .C1(new_n443_), .C2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(G183gat), .A2(G190gat), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n368_), .B1(new_n381_), .B2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n437_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n420_), .B1(new_n435_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n420_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT20), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT90), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n436_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n427_), .A2(KEYINPUT90), .A3(new_n428_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n452_), .B1(new_n456_), .B2(new_n402_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n373_), .A2(new_n387_), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n441_), .A2(KEYINPUT94), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n458_), .B1(new_n459_), .B2(new_n442_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n447_), .ZN(new_n461_));
  NOR3_X1   g260(.A1(new_n460_), .A2(new_n436_), .A3(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT95), .ZN(new_n463_));
  NOR3_X1   g262(.A1(new_n457_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n451_), .B1(new_n431_), .B2(new_n434_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n445_), .A2(new_n437_), .A3(new_n447_), .ZN(new_n466_));
  AOI21_X1  g265(.A(KEYINPUT95), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n449_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n468_));
  XOR2_X1   g267(.A(G8gat), .B(G36gat), .Z(new_n469_));
  XNOR2_X1  g268(.A(G64gat), .B(G92gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n472_));
  XOR2_X1   g271(.A(new_n471_), .B(new_n472_), .Z(new_n473_));
  NAND2_X1  g272(.A1(new_n468_), .A2(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n463_), .B1(new_n457_), .B2(new_n462_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n465_), .A2(KEYINPUT95), .A3(new_n466_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n473_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(new_n449_), .A3(new_n478_), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n474_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G1gat), .B(G29gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(G85gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT0), .B(G57gat), .ZN(new_n483_));
  XOR2_X1   g282(.A(new_n482_), .B(new_n483_), .Z(new_n484_));
  NAND2_X1  g283(.A1(G225gat), .A2(G233gat), .ZN(new_n485_));
  NOR2_X1   g284(.A1(G155gat), .A2(G162gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G155gat), .A2(G162gat), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n486_), .B1(KEYINPUT1), .B2(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n488_), .B1(KEYINPUT1), .B2(new_n487_), .ZN(new_n489_));
  INV_X1    g288(.A(G141gat), .ZN(new_n490_));
  INV_X1    g289(.A(G148gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G141gat), .A2(G148gat), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n489_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(KEYINPUT3), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT2), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n495_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT86), .B(KEYINPUT3), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT87), .ZN(new_n501_));
  OR3_X1    g300(.A1(new_n500_), .A2(new_n501_), .A3(new_n492_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n501_), .B1(new_n500_), .B2(new_n492_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n499_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n486_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(new_n487_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n494_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(new_n410_), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n409_), .B(new_n494_), .C1(new_n504_), .C2(new_n506_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(KEYINPUT4), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT4), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n507_), .A2(new_n511_), .A3(new_n410_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n485_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n485_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n514_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n484_), .B1(new_n513_), .B2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT33), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n510_), .A2(new_n485_), .A3(new_n512_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n484_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n508_), .A2(new_n509_), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n518_), .B(new_n519_), .C1(new_n485_), .C2(new_n520_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n480_), .A2(new_n517_), .A3(KEYINPUT97), .A4(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT97), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT33), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n516_), .B(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n474_), .A2(new_n479_), .A3(new_n521_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n523_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT99), .ZN(new_n528_));
  XOR2_X1   g327(.A(KEYINPUT98), .B(KEYINPUT20), .Z(new_n529_));
  NAND3_X1  g328(.A1(new_n466_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n530_), .B1(new_n456_), .B2(new_n402_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n528_), .B1(new_n466_), .B2(new_n529_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n420_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  OR3_X1    g332(.A1(new_n435_), .A2(new_n420_), .A3(new_n448_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n478_), .A2(KEYINPUT32), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n535_), .A2(new_n537_), .ZN(new_n538_));
  OR4_X1    g337(.A1(KEYINPUT100), .A2(new_n513_), .A3(new_n484_), .A4(new_n515_), .ZN(new_n539_));
  OR3_X1    g338(.A1(new_n513_), .A2(new_n484_), .A3(new_n515_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n540_), .A2(KEYINPUT100), .A3(new_n516_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n477_), .A2(new_n449_), .A3(new_n536_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n538_), .A2(new_n539_), .A3(new_n541_), .A4(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n522_), .A2(new_n527_), .A3(new_n543_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n507_), .A2(KEYINPUT29), .ZN(new_n545_));
  XOR2_X1   g344(.A(KEYINPUT88), .B(KEYINPUT28), .Z(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(G22gat), .B(G50gat), .Z(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n507_), .A2(KEYINPUT29), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT91), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n507_), .A2(KEYINPUT91), .A3(KEYINPUT29), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n553_), .A2(new_n554_), .A3(new_n436_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT89), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n556_), .A2(G228gat), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(G228gat), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n316_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n456_), .A2(new_n559_), .ZN(new_n560_));
  AOI22_X1  g359(.A1(new_n555_), .A2(new_n559_), .B1(new_n551_), .B2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G78gat), .B(G106gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT92), .Z(new_n563_));
  AOI21_X1  g362(.A(KEYINPUT93), .B1(new_n561_), .B2(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n561_), .A2(new_n563_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n561_), .A2(KEYINPUT93), .A3(new_n563_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n550_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n561_), .A2(new_n563_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n562_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n549_), .B(new_n569_), .C1(new_n570_), .C2(new_n561_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n568_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n544_), .A2(new_n572_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n541_), .A2(new_n539_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n574_), .B1(new_n568_), .B2(new_n571_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n535_), .A2(new_n473_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n479_), .A2(KEYINPUT27), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n474_), .A2(new_n479_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT27), .ZN(new_n579_));
  AOI22_X1  g378(.A1(new_n576_), .A2(new_n577_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n575_), .A2(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n418_), .B1(new_n573_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n572_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n580_), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n574_), .A2(new_n417_), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n583_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n582_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G229gat), .A2(G233gat), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n342_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(new_n314_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n342_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n591_), .A2(KEYINPUT77), .A3(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(KEYINPUT77), .B1(new_n591_), .B2(new_n592_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n589_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n343_), .A2(new_n314_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n596_), .A2(new_n592_), .A3(new_n588_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G113gat), .B(G141gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G169gat), .B(G197gat), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n598_), .B(new_n599_), .Z(new_n600_));
  NAND3_X1  g399(.A1(new_n595_), .A2(new_n597_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT78), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n595_), .A2(new_n597_), .A3(KEYINPUT78), .A4(new_n600_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n595_), .A2(new_n597_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n600_), .ZN(new_n606_));
  AOI22_X1  g405(.A1(new_n603_), .A2(new_n604_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n587_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n366_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n574_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n609_), .A2(G1gat), .A3(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n612_));
  OR2_X1    g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n295_), .A2(new_n607_), .A3(new_n336_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n361_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n587_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(G1gat), .B1(new_n617_), .B2(new_n610_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n611_), .A2(new_n612_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n613_), .A2(new_n618_), .A3(new_n619_), .ZN(G1324gat));
  INV_X1    g419(.A(KEYINPUT39), .ZN(new_n621_));
  INV_X1    g420(.A(new_n617_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(new_n584_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n621_), .B1(new_n623_), .B2(G8gat), .ZN(new_n624_));
  AOI211_X1 g423(.A(KEYINPUT39), .B(new_n303_), .C1(new_n622_), .C2(new_n584_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n584_), .A2(new_n303_), .ZN(new_n626_));
  OAI22_X1  g425(.A1(new_n624_), .A2(new_n625_), .B1(new_n609_), .B2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n627_), .B(new_n629_), .ZN(G1325gat));
  INV_X1    g429(.A(new_n418_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G15gat), .B1(new_n617_), .B2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT41), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n609_), .A2(G15gat), .A3(new_n631_), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n633_), .A2(new_n634_), .ZN(G1326gat));
  OAI21_X1  g434(.A(G22gat), .B1(new_n617_), .B2(new_n572_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT42), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n572_), .A2(G22gat), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n637_), .B1(new_n609_), .B2(new_n638_), .ZN(G1327gat));
  INV_X1    g438(.A(new_n336_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n361_), .A2(new_n640_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n293_), .A2(new_n294_), .A3(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n608_), .A2(new_n642_), .ZN(new_n643_));
  OR3_X1    g442(.A1(new_n643_), .A2(G29gat), .A3(new_n610_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n365_), .B1(new_n582_), .B2(new_n586_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT43), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n640_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n295_), .A2(new_n607_), .ZN(new_n648_));
  OAI211_X1 g447(.A(KEYINPUT43), .B(new_n365_), .C1(new_n582_), .C2(new_n586_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n647_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT44), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n647_), .A2(KEYINPUT44), .A3(new_n648_), .A4(new_n649_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n653_), .A2(KEYINPUT103), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(KEYINPUT103), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n574_), .B(new_n652_), .C1(new_n654_), .C2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT104), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n656_), .A2(new_n657_), .A3(G29gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n656_), .B2(G29gat), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n644_), .B1(new_n658_), .B2(new_n659_), .ZN(G1328gat));
  INV_X1    g459(.A(KEYINPUT46), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n661_), .A2(KEYINPUT106), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n584_), .B(new_n652_), .C1(new_n654_), .C2(new_n655_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(G36gat), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n661_), .A2(KEYINPUT106), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n580_), .A2(G36gat), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n608_), .A2(new_n642_), .A3(new_n667_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n668_), .A2(new_n670_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n666_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n663_), .B1(new_n665_), .B2(new_n674_), .ZN(new_n675_));
  AOI211_X1 g474(.A(new_n662_), .B(new_n673_), .C1(new_n664_), .C2(G36gat), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1329gat));
  AND2_X1   g476(.A1(new_n650_), .A2(new_n651_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n647_), .A2(new_n649_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n679_), .A2(new_n680_), .A3(KEYINPUT44), .A4(new_n648_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n653_), .A2(KEYINPUT103), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n678_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n417_), .A2(new_n413_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n413_), .B1(new_n643_), .B2(new_n631_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT47), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT47), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n685_), .A2(new_n689_), .A3(new_n686_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(G1330gat));
  INV_X1    g490(.A(G50gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n683_), .B2(new_n583_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n643_), .A2(G50gat), .A3(new_n572_), .ZN(new_n694_));
  OAI21_X1  g493(.A(KEYINPUT107), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n652_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n696_));
  OAI21_X1  g495(.A(G50gat), .B1(new_n696_), .B2(new_n572_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT107), .ZN(new_n698_));
  INV_X1    g497(.A(new_n694_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n697_), .A2(new_n698_), .A3(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n695_), .A2(new_n700_), .ZN(G1331gat));
  INV_X1    g500(.A(G57gat), .ZN(new_n702_));
  INV_X1    g501(.A(new_n607_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n587_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n365_), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n704_), .A2(new_n295_), .A3(new_n640_), .A4(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n702_), .B1(new_n706_), .B2(new_n610_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT108), .Z(new_n708_));
  AND2_X1   g507(.A1(new_n293_), .A2(new_n294_), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n709_), .A2(new_n703_), .A3(new_n336_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n710_), .A2(new_n616_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n610_), .A2(new_n702_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n708_), .B1(new_n711_), .B2(new_n712_), .ZN(G1332gat));
  OR3_X1    g512(.A1(new_n706_), .A2(G64gat), .A3(new_n580_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n711_), .ZN(new_n715_));
  OAI21_X1  g514(.A(G64gat), .B1(new_n715_), .B2(new_n580_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n716_), .A2(KEYINPUT48), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n716_), .A2(KEYINPUT48), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n714_), .B1(new_n717_), .B2(new_n718_), .ZN(G1333gat));
  OR3_X1    g518(.A1(new_n706_), .A2(G71gat), .A3(new_n631_), .ZN(new_n720_));
  OAI21_X1  g519(.A(G71gat), .B1(new_n715_), .B2(new_n631_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n721_), .A2(KEYINPUT49), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(KEYINPUT49), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n720_), .B1(new_n722_), .B2(new_n723_), .ZN(G1334gat));
  OR3_X1    g523(.A1(new_n706_), .A2(G78gat), .A3(new_n572_), .ZN(new_n725_));
  OAI21_X1  g524(.A(G78gat), .B1(new_n715_), .B2(new_n572_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(KEYINPUT50), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n726_), .A2(KEYINPUT50), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n725_), .B1(new_n727_), .B2(new_n728_), .ZN(G1335gat));
  NOR2_X1   g528(.A1(new_n709_), .A2(new_n703_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n730_), .A2(new_n647_), .A3(new_n649_), .ZN(new_n731_));
  OAI21_X1  g530(.A(G85gat), .B1(new_n731_), .B2(new_n610_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n704_), .A2(new_n295_), .A3(new_n641_), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n610_), .A2(G85gat), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n732_), .B1(new_n733_), .B2(new_n734_), .ZN(G1336gat));
  OAI21_X1  g534(.A(G92gat), .B1(new_n731_), .B2(new_n580_), .ZN(new_n736_));
  OR2_X1    g535(.A1(new_n580_), .A2(G92gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n736_), .B1(new_n733_), .B2(new_n737_), .ZN(G1337gat));
  INV_X1    g537(.A(new_n733_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n417_), .A2(new_n227_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n730_), .A2(new_n647_), .A3(new_n418_), .A4(new_n649_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT109), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(new_n744_), .A3(G99gat), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n744_), .B1(new_n743_), .B2(G99gat), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n741_), .B(new_n742_), .C1(new_n746_), .C2(new_n747_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n748_), .A2(KEYINPUT111), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n748_), .A2(KEYINPUT111), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n741_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT51), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n749_), .B1(new_n750_), .B2(new_n752_), .ZN(G1338gat));
  OR3_X1    g552(.A1(new_n733_), .A2(new_n572_), .A3(new_n228_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n755_));
  OAI21_X1  g554(.A(G106gat), .B1(new_n731_), .B2(new_n572_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n756_), .A2(KEYINPUT52), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n756_), .A2(KEYINPUT52), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n754_), .B(new_n755_), .C1(new_n757_), .C2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n756_), .B(KEYINPUT52), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n755_), .B1(new_n761_), .B2(new_n754_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1339gat));
  INV_X1    g562(.A(KEYINPUT118), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n703_), .A2(new_n285_), .ZN(new_n765_));
  OAI21_X1  g564(.A(KEYINPUT55), .B1(new_n202_), .B2(KEYINPUT115), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n766_), .B1(KEYINPUT55), .B2(new_n202_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n274_), .A2(new_n276_), .A3(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n254_), .B1(KEYINPUT12), .B2(new_n252_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n270_), .A2(new_n231_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n272_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n270_), .A2(KEYINPUT69), .A3(new_n231_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n770_), .B1(new_n774_), .B2(new_n258_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n282_), .B(new_n769_), .C1(new_n775_), .C2(new_n766_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT56), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT116), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n776_), .A2(new_n777_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n776_), .A2(KEYINPUT116), .A3(new_n777_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n765_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n588_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n592_), .A2(new_n589_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n600_), .B1(new_n596_), .B2(new_n785_), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n603_), .A2(new_n604_), .B1(new_n783_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n788_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n361_), .B1(new_n782_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT57), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  OAI211_X1 g591(.A(KEYINPUT117), .B(new_n361_), .C1(new_n782_), .C2(new_n789_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n764_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT116), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n274_), .A2(new_n276_), .A3(new_n768_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n766_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n797_));
  NOR3_X1   g596(.A1(new_n796_), .A2(new_n797_), .A3(new_n284_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n795_), .B1(new_n798_), .B2(KEYINPUT56), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(KEYINPUT56), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(new_n781_), .A3(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n765_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n789_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n791_), .B1(new_n803_), .B2(new_n615_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n804_), .A2(new_n793_), .A3(new_n764_), .A4(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n801_), .A2(new_n802_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n789_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n615_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n285_), .A2(new_n787_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n776_), .A2(new_n777_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n810_), .B1(new_n800_), .B2(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(KEYINPUT119), .A2(KEYINPUT58), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n812_), .B(new_n813_), .ZN(new_n814_));
  AOI22_X1  g613(.A1(KEYINPUT57), .A2(new_n809_), .B1(new_n814_), .B2(new_n365_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n806_), .A2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n336_), .B1(new_n794_), .B2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(KEYINPUT113), .B1(new_n640_), .B2(new_n607_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT113), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n336_), .A2(new_n819_), .A3(new_n703_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n291_), .A2(new_n818_), .A3(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n705_), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT114), .B1(new_n822_), .B2(KEYINPUT54), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(KEYINPUT54), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT114), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n821_), .A2(new_n705_), .A3(new_n825_), .A4(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n823_), .A2(new_n824_), .A3(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n817_), .A2(new_n828_), .ZN(new_n829_));
  NOR4_X1   g628(.A1(new_n583_), .A2(new_n610_), .A3(new_n584_), .A4(new_n417_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(G113gat), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n832_), .A3(new_n703_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT59), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n831_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n830_), .A2(new_n834_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n804_), .A2(new_n793_), .A3(new_n805_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n814_), .A2(new_n365_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n837_), .A2(new_n838_), .A3(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n809_), .A2(KEYINPUT57), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n838_), .B1(new_n837_), .B2(new_n839_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n336_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n836_), .B1(new_n844_), .B2(new_n828_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n835_), .A2(new_n845_), .A3(new_n607_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n833_), .B1(new_n846_), .B2(new_n832_), .ZN(G1340gat));
  INV_X1    g646(.A(KEYINPUT60), .ZN(new_n848_));
  AOI21_X1  g647(.A(KEYINPUT121), .B1(new_n848_), .B2(G120gat), .ZN(new_n849_));
  AOI21_X1  g648(.A(G120gat), .B1(new_n295_), .B2(new_n848_), .ZN(new_n850_));
  MUX2_X1   g649(.A(new_n849_), .B(KEYINPUT121), .S(new_n850_), .Z(new_n851_));
  NAND2_X1  g650(.A1(new_n831_), .A2(new_n851_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n835_), .A2(new_n845_), .A3(new_n709_), .ZN(new_n853_));
  INV_X1    g652(.A(G120gat), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n852_), .B1(new_n853_), .B2(new_n854_), .ZN(G1341gat));
  INV_X1    g654(.A(G127gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n831_), .A2(new_n856_), .A3(new_n640_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n835_), .A2(new_n845_), .A3(new_n336_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n856_), .ZN(G1342gat));
  INV_X1    g658(.A(G134gat), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n831_), .A2(new_n860_), .A3(new_n615_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n835_), .A2(new_n845_), .A3(new_n705_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n862_), .B2(new_n860_), .ZN(G1343gat));
  AOI21_X1  g662(.A(new_n418_), .B1(new_n817_), .B2(new_n828_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n572_), .A2(new_n584_), .A3(new_n610_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n607_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(new_n490_), .ZN(G1344gat));
  NOR2_X1   g667(.A1(new_n866_), .A2(new_n709_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(new_n491_), .ZN(G1345gat));
  NAND3_X1  g669(.A1(new_n864_), .A2(new_n640_), .A3(new_n865_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(KEYINPUT122), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n864_), .A2(new_n873_), .A3(new_n640_), .A4(new_n865_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(KEYINPUT61), .B(G155gat), .ZN(new_n875_));
  AND3_X1   g674(.A1(new_n872_), .A2(new_n874_), .A3(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1346gat));
  OAI21_X1  g677(.A(G162gat), .B1(new_n866_), .B2(new_n705_), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n361_), .A2(G162gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n866_), .B2(new_n880_), .ZN(G1347gat));
  NAND2_X1  g680(.A1(new_n844_), .A2(new_n828_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT22), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n418_), .A2(new_n610_), .A3(new_n584_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n583_), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n882_), .A2(new_n883_), .A3(new_n703_), .A4(new_n885_), .ZN(new_n886_));
  AND3_X1   g685(.A1(new_n886_), .A2(KEYINPUT62), .A3(new_n384_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(KEYINPUT62), .ZN(new_n888_));
  AND3_X1   g687(.A1(new_n882_), .A2(new_n703_), .A3(new_n885_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n384_), .B1(new_n889_), .B2(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n887_), .B1(new_n888_), .B2(new_n891_), .ZN(G1348gat));
  NAND3_X1  g691(.A1(new_n882_), .A2(new_n295_), .A3(new_n885_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n583_), .B1(new_n817_), .B2(new_n828_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n709_), .A2(new_n385_), .A3(new_n884_), .ZN(new_n895_));
  AOI22_X1  g694(.A1(new_n893_), .A2(new_n385_), .B1(new_n894_), .B2(new_n895_), .ZN(G1349gat));
  NOR2_X1   g695(.A1(new_n336_), .A2(new_n439_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n882_), .A2(new_n885_), .A3(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n884_), .A2(new_n336_), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n829_), .A2(KEYINPUT123), .A3(new_n572_), .A4(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n377_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(KEYINPUT123), .B1(new_n894_), .B2(new_n899_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n898_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  OAI211_X1 g705(.A(KEYINPUT124), .B(new_n898_), .C1(new_n902_), .C2(new_n903_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(G1350gat));
  NAND2_X1  g707(.A1(new_n882_), .A2(new_n885_), .ZN(new_n909_));
  OAI21_X1  g708(.A(G190gat), .B1(new_n909_), .B2(new_n705_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n615_), .A2(new_n438_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n909_), .B2(new_n911_), .ZN(G1351gat));
  NAND2_X1  g711(.A1(new_n575_), .A2(new_n584_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(new_n914_));
  AND2_X1   g713(.A1(new_n864_), .A2(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n703_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g716(.A1(new_n915_), .A2(new_n295_), .ZN(new_n918_));
  XOR2_X1   g717(.A(KEYINPUT125), .B(G204gat), .Z(new_n919_));
  XNOR2_X1  g718(.A(new_n918_), .B(new_n919_), .ZN(G1353gat));
  INV_X1    g719(.A(KEYINPUT63), .ZN(new_n921_));
  INV_X1    g720(.A(G211gat), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n640_), .B1(new_n921_), .B2(new_n922_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(KEYINPUT126), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n915_), .A2(new_n924_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n921_), .A2(new_n922_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n925_), .B(new_n926_), .ZN(G1354gat));
  INV_X1    g726(.A(G218gat), .ZN(new_n928_));
  NAND4_X1  g727(.A1(new_n864_), .A2(new_n928_), .A3(new_n615_), .A4(new_n914_), .ZN(new_n929_));
  AND3_X1   g728(.A1(new_n864_), .A2(new_n365_), .A3(new_n914_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n930_), .B2(new_n928_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT127), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  OAI211_X1 g732(.A(new_n929_), .B(KEYINPUT127), .C1(new_n930_), .C2(new_n928_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(G1355gat));
endmodule


