//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 0 0 0 0 0 1 1 0 1 1 1 0 0 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n762_, new_n763_, new_n764_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n777_, new_n778_,
    new_n779_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n900_, new_n902_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_, new_n927_, new_n929_,
    new_n930_, new_n932_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n949_, new_n950_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_;
  INV_X1    g000(.A(KEYINPUT68), .ZN(new_n202_));
  XOR2_X1   g001(.A(G120gat), .B(G148gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(G176gat), .B(G204gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(KEYINPUT10), .B(G99gat), .Z(new_n208_));
  INV_X1    g007(.A(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT65), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G99gat), .A2(G106gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G85gat), .ZN(new_n216_));
  INV_X1    g015(.A(G92gat), .ZN(new_n217_));
  NOR3_X1   g016(.A1(new_n216_), .A2(new_n217_), .A3(KEYINPUT9), .ZN(new_n218_));
  XOR2_X1   g017(.A(G85gat), .B(G92gat), .Z(new_n219_));
  AOI21_X1  g018(.A(new_n218_), .B1(new_n219_), .B2(KEYINPUT9), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n211_), .A2(new_n215_), .A3(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G99gat), .A2(G106gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT7), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n219_), .B1(new_n224_), .B2(new_n214_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT8), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n221_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G57gat), .B(G64gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT11), .ZN(new_n229_));
  XOR2_X1   g028(.A(G71gat), .B(G78gat), .Z(new_n230_));
  OR2_X1    g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n228_), .A2(KEYINPUT11), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n229_), .A2(new_n230_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n231_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n227_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT12), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G230gat), .A2(G233gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n238_), .B(KEYINPUT64), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n227_), .A2(new_n234_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n227_), .A2(new_n236_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n234_), .B(KEYINPUT66), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n237_), .A2(new_n240_), .A3(new_n241_), .A4(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n235_), .A2(new_n241_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(new_n239_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n207_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n245_), .A2(new_n247_), .A3(new_n207_), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT13), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n250_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT13), .ZN(new_n253_));
  NOR3_X1   g052(.A1(new_n252_), .A2(new_n253_), .A3(new_n248_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n202_), .B1(new_n251_), .B2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n253_), .B1(new_n252_), .B2(new_n248_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n249_), .A2(KEYINPUT13), .A3(new_n250_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(new_n257_), .A3(KEYINPUT68), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n255_), .A2(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(G127gat), .B(G155gat), .Z(new_n260_));
  XNOR2_X1  g059(.A(G183gat), .B(G211gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(KEYINPUT73), .B(KEYINPUT16), .Z(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT17), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G1gat), .B(G8gat), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n267_), .A2(KEYINPUT71), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(KEYINPUT71), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G15gat), .B(G22gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G1gat), .A2(G8gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT14), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n270_), .A2(new_n274_), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n268_), .A2(new_n273_), .A3(new_n271_), .A4(new_n269_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G231gat), .A2(G233gat), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n278_), .B(KEYINPUT72), .Z(new_n279_));
  XNOR2_X1  g078(.A(new_n277_), .B(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n266_), .B1(new_n234_), .B2(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n281_), .B1(new_n234_), .B2(new_n280_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n280_), .A2(new_n243_), .ZN(new_n283_));
  NOR3_X1   g082(.A1(new_n283_), .A2(new_n265_), .A3(new_n264_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n280_), .A2(new_n243_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n282_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(G29gat), .B(G36gat), .Z(new_n289_));
  XOR2_X1   g088(.A(G43gat), .B(G50gat), .Z(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n277_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT74), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n293_), .B1(new_n277_), .B2(new_n291_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G229gat), .A2(G233gat), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT75), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n294_), .A2(KEYINPUT75), .A3(new_n296_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT74), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n292_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n277_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n291_), .B(KEYINPUT15), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n302_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n295_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n299_), .A2(new_n300_), .A3(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(G113gat), .B(G141gat), .Z(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT76), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G169gat), .B(G197gat), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n309_), .B(new_n310_), .Z(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n307_), .A2(new_n312_), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n299_), .A2(new_n300_), .A3(new_n306_), .A4(new_n311_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n259_), .A2(new_n288_), .A3(new_n315_), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n316_), .A2(KEYINPUT101), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G226gat), .A2(G233gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT19), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G211gat), .B(G218gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT21), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G197gat), .B(G204gat), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n321_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(G197gat), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n325_), .A2(KEYINPUT87), .A3(G204gat), .ZN(new_n326_));
  INV_X1    g125(.A(new_n323_), .ZN(new_n327_));
  OAI211_X1 g126(.A(KEYINPUT21), .B(new_n326_), .C1(new_n327_), .C2(KEYINPUT87), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n323_), .A2(new_n322_), .ZN(new_n329_));
  AOI22_X1  g128(.A1(new_n324_), .A2(new_n328_), .B1(new_n321_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(G183gat), .ZN(new_n331_));
  INV_X1    g130(.A(G190gat), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT23), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n331_), .A2(KEYINPUT23), .ZN(new_n334_));
  AOI21_X1  g133(.A(KEYINPUT79), .B1(new_n334_), .B2(G190gat), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT23), .ZN(new_n336_));
  NAND4_X1  g135(.A1(new_n336_), .A2(KEYINPUT79), .A3(G183gat), .A4(G190gat), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n333_), .B1(new_n335_), .B2(new_n338_), .ZN(new_n339_));
  NOR3_X1   g138(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(KEYINPUT80), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT80), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n336_), .B1(G183gat), .B2(G190gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n336_), .A2(G183gat), .A3(G190gat), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT79), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n344_), .B1(new_n347_), .B2(new_n337_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n343_), .B1(new_n348_), .B2(new_n340_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n331_), .A2(KEYINPUT25), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT25), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(G183gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT26), .ZN(new_n354_));
  AOI21_X1  g153(.A(KEYINPUT77), .B1(new_n354_), .B2(G190gat), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(G190gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n332_), .A2(KEYINPUT26), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT77), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G169gat), .A2(G176gat), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AOI22_X1  g164(.A1(new_n356_), .A2(new_n360_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n342_), .A2(new_n349_), .A3(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT22), .B(G169gat), .ZN(new_n368_));
  INV_X1    g167(.A(G176gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n363_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT81), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n333_), .A2(new_n345_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(G183gat), .A2(G190gat), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT81), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n370_), .A2(new_n363_), .A3(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n372_), .A2(new_n376_), .A3(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n330_), .B1(new_n367_), .B2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n340_), .B1(new_n333_), .B2(new_n345_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n357_), .A2(new_n358_), .A3(new_n350_), .A4(new_n352_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n361_), .A2(KEYINPUT89), .A3(KEYINPUT24), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n383_), .B1(G169gat), .B2(G176gat), .ZN(new_n384_));
  AOI21_X1  g183(.A(KEYINPUT89), .B1(new_n361_), .B2(KEYINPUT24), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n381_), .B(new_n382_), .C1(new_n384_), .C2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n348_), .A2(new_n374_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n386_), .B1(new_n387_), .B2(new_n371_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n329_), .A2(new_n321_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n320_), .B1(new_n327_), .B2(KEYINPUT21), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n326_), .A2(KEYINPUT21), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT87), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n391_), .B1(new_n392_), .B2(new_n323_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n389_), .B1(new_n390_), .B2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT20), .B1(new_n388_), .B2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n319_), .B1(new_n380_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT96), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n367_), .A2(new_n330_), .A3(new_n379_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT20), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n400_), .B1(new_n388_), .B2(new_n394_), .ZN(new_n401_));
  XOR2_X1   g200(.A(new_n319_), .B(KEYINPUT88), .Z(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n399_), .A2(new_n401_), .A3(new_n403_), .ZN(new_n404_));
  OAI211_X1 g203(.A(KEYINPUT96), .B(new_n319_), .C1(new_n380_), .C2(new_n395_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n398_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(G8gat), .B(G36gat), .Z(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G64gat), .B(G92gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n406_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT98), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT27), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n367_), .A2(new_n379_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n394_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n319_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n339_), .A2(new_n375_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n371_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n381_), .A2(new_n382_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n385_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n421_), .B(new_n383_), .C1(G169gat), .C2(G176gat), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n418_), .A2(new_n419_), .B1(new_n420_), .B2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n400_), .B1(new_n423_), .B2(new_n330_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n416_), .A2(KEYINPUT90), .A3(new_n417_), .A4(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n399_), .A2(new_n401_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(new_n402_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n380_), .A2(new_n395_), .ZN(new_n429_));
  AOI21_X1  g228(.A(KEYINPUT90), .B1(new_n429_), .B2(new_n417_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n428_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n411_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n414_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT98), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n406_), .A2(new_n434_), .A3(new_n411_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n413_), .A2(new_n433_), .A3(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G22gat), .B(G50gat), .ZN(new_n437_));
  INV_X1    g236(.A(G141gat), .ZN(new_n438_));
  INV_X1    g237(.A(G148gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G141gat), .A2(G148gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(G155gat), .A2(G162gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G155gat), .A2(G162gat), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n443_), .B1(KEYINPUT1), .B2(new_n444_), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n444_), .A2(KEYINPUT1), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n442_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT3), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n448_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT84), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n441_), .A2(KEYINPUT2), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT2), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n453_), .A2(G141gat), .A3(G148gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n440_), .A2(KEYINPUT3), .ZN(new_n456_));
  NOR2_X1   g255(.A1(G141gat), .A2(G148gat), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n457_), .A2(KEYINPUT84), .A3(new_n448_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n451_), .A2(new_n455_), .A3(new_n456_), .A4(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n444_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n460_), .A2(new_n443_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n447_), .B1(new_n459_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT29), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT28), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n464_), .A2(KEYINPUT28), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n437_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n467_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n437_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n469_), .A2(new_n465_), .A3(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n468_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n459_), .A2(new_n461_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n447_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n463_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(G78gat), .B1(new_n475_), .B2(new_n330_), .ZN(new_n476_));
  INV_X1    g275(.A(G78gat), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n394_), .B(new_n477_), .C1(new_n462_), .C2(new_n463_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n476_), .A2(G106gat), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(G106gat), .B1(new_n476_), .B2(new_n478_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G228gat), .A2(G233gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT86), .ZN(new_n482_));
  OR2_X1    g281(.A1(new_n481_), .A2(KEYINPUT86), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n482_), .B(new_n483_), .C1(new_n330_), .C2(KEYINPUT85), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NOR3_X1   g284(.A1(new_n479_), .A2(new_n480_), .A3(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n478_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n461_), .ZN(new_n488_));
  NOR4_X1   g287(.A1(new_n450_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n489_));
  AOI21_X1  g288(.A(KEYINPUT84), .B1(new_n457_), .B2(new_n448_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  AOI22_X1  g290(.A1(new_n452_), .A2(new_n454_), .B1(new_n440_), .B2(KEYINPUT3), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n488_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT29), .B1(new_n493_), .B2(new_n447_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n477_), .B1(new_n494_), .B2(new_n394_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n209_), .B1(new_n487_), .B2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n476_), .A2(G106gat), .A3(new_n478_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n484_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n472_), .B1(new_n486_), .B2(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n485_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n496_), .A2(new_n497_), .A3(new_n484_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n500_), .A2(new_n501_), .A3(new_n471_), .A4(new_n468_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n499_), .A2(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n411_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n416_), .A2(new_n417_), .A3(new_n424_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT90), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n507_), .A2(new_n432_), .A3(new_n427_), .A4(new_n425_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n504_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n414_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n436_), .A2(new_n503_), .A3(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(G1gat), .B(G29gat), .Z(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G57gat), .B(G85gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G225gat), .A2(G233gat), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT92), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G127gat), .B(G134gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G113gat), .B(G120gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n519_), .B1(new_n462_), .B2(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(new_n520_), .B(new_n521_), .Z(new_n524_));
  OAI211_X1 g323(.A(new_n524_), .B(KEYINPUT92), .C1(new_n493_), .C2(new_n447_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n473_), .A2(new_n474_), .A3(new_n522_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT93), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT93), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n462_), .A2(new_n529_), .A3(new_n522_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT4), .B1(new_n526_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n473_), .A2(new_n474_), .ZN(new_n533_));
  AOI21_X1  g332(.A(KEYINPUT4), .B1(new_n533_), .B2(new_n524_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n518_), .B1(new_n532_), .B2(new_n535_), .ZN(new_n536_));
  AND4_X1   g335(.A1(new_n529_), .A2(new_n473_), .A3(new_n474_), .A4(new_n522_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n529_), .B1(new_n462_), .B2(new_n522_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n523_), .A2(new_n525_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n539_), .A2(new_n518_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n517_), .B1(new_n536_), .B2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(KEYINPUT92), .B1(new_n533_), .B2(new_n524_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n462_), .A2(new_n519_), .A3(new_n522_), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n528_), .B(new_n530_), .C1(new_n544_), .C2(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n534_), .B1(new_n546_), .B2(KEYINPUT4), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n516_), .B(new_n541_), .C1(new_n547_), .C2(new_n518_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n543_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G71gat), .B(G99gat), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n367_), .A2(KEYINPUT30), .A3(new_n379_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(KEYINPUT30), .B1(new_n367_), .B2(new_n379_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n551_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n554_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n551_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n556_), .A2(new_n557_), .A3(new_n552_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n555_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G227gat), .A2(G233gat), .ZN(new_n560_));
  INV_X1    g359(.A(G15gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(G43gat), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n559_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT83), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n522_), .B(KEYINPUT31), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT82), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n565_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n563_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n555_), .A2(new_n558_), .A3(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n564_), .A2(new_n568_), .A3(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n568_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n570_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n569_), .B1(new_n555_), .B2(new_n558_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n572_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n550_), .A2(new_n571_), .A3(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(KEYINPUT99), .B1(new_n511_), .B2(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n434_), .B1(new_n406_), .B2(new_n411_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n508_), .A2(KEYINPUT27), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  AOI22_X1  g379(.A1(new_n580_), .A2(new_n435_), .B1(new_n414_), .B2(new_n509_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT99), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n575_), .A2(new_n571_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n583_), .A2(new_n549_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n581_), .A2(new_n582_), .A3(new_n503_), .A4(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n577_), .A2(new_n585_), .ZN(new_n586_));
  AND4_X1   g385(.A1(new_n548_), .A2(new_n543_), .A3(new_n502_), .A4(new_n499_), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n587_), .A2(new_n436_), .A3(new_n510_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n518_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT4), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n590_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n589_), .B1(new_n591_), .B2(new_n534_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n592_), .A2(KEYINPUT33), .A3(new_n516_), .A4(new_n541_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n546_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n516_), .B1(new_n594_), .B2(new_n589_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n595_), .B1(new_n589_), .B2(new_n547_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n593_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT33), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n548_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT95), .ZN(new_n600_));
  INV_X1    g399(.A(new_n509_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT95), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n548_), .A2(new_n602_), .A3(new_n598_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n597_), .A2(new_n600_), .A3(new_n601_), .A4(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n432_), .A2(KEYINPUT32), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n431_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n406_), .A2(KEYINPUT32), .A3(new_n432_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n548_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n516_), .B1(new_n592_), .B2(new_n541_), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n606_), .B(new_n607_), .C1(new_n608_), .C2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT97), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT97), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n549_), .A2(new_n612_), .A3(new_n606_), .A4(new_n607_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n604_), .A2(new_n611_), .A3(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n588_), .B1(new_n614_), .B2(new_n503_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n583_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n586_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n291_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n227_), .A2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n620_));
  NAND2_X1  g419(.A1(G232gat), .A2(G233gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT35), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n619_), .B(new_n624_), .C1(new_n304_), .C2(new_n227_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT70), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n227_), .A2(new_n304_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT70), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n627_), .A2(new_n628_), .A3(new_n624_), .A4(new_n619_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n619_), .B1(new_n304_), .B2(new_n227_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n622_), .B(KEYINPUT35), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n626_), .A2(new_n629_), .A3(new_n632_), .ZN(new_n633_));
  XOR2_X1   g432(.A(G134gat), .B(G162gat), .Z(new_n634_));
  XNOR2_X1  g433(.A(G190gat), .B(G218gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT36), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n636_), .A2(new_n637_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n633_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  AOI22_X1  g439(.A1(new_n625_), .A2(KEYINPUT70), .B1(new_n630_), .B2(new_n631_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n641_), .A2(new_n637_), .A3(new_n636_), .A4(new_n629_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT102), .Z(new_n644_));
  AND2_X1   g443(.A1(new_n617_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n316_), .A2(KEYINPUT101), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n317_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT103), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(new_n549_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(G1gat), .ZN(new_n650_));
  INV_X1    g449(.A(new_n259_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n617_), .A2(new_n315_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT100), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n617_), .A2(KEYINPUT100), .A3(new_n315_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n651_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT37), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n643_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n640_), .A2(KEYINPUT37), .A3(new_n642_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n660_), .A2(new_n287_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n656_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT38), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n550_), .A2(G1gat), .ZN(new_n664_));
  OR3_X1    g463(.A1(new_n662_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n663_), .B1(new_n662_), .B2(new_n664_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n650_), .A2(new_n665_), .A3(new_n666_), .ZN(G1324gat));
  OAI21_X1  g466(.A(G8gat), .B1(new_n647_), .B2(new_n581_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT39), .ZN(new_n669_));
  OR3_X1    g468(.A1(new_n662_), .A2(G8gat), .A3(new_n581_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n669_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1325gat));
  INV_X1    g473(.A(new_n662_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n675_), .A2(new_n561_), .A3(new_n616_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n648_), .A2(new_n616_), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n677_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(KEYINPUT41), .B1(new_n677_), .B2(G15gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n676_), .B1(new_n678_), .B2(new_n679_), .ZN(G1326gat));
  INV_X1    g479(.A(G22gat), .ZN(new_n681_));
  INV_X1    g480(.A(new_n503_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n675_), .A2(new_n681_), .A3(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n648_), .A2(new_n682_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n685_), .B2(G22gat), .ZN(new_n686_));
  AOI211_X1 g485(.A(KEYINPUT42), .B(new_n681_), .C1(new_n648_), .C2(new_n682_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n683_), .B1(new_n686_), .B2(new_n687_), .ZN(G1327gat));
  NOR2_X1   g487(.A1(new_n643_), .A2(new_n288_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n656_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(G29gat), .B1(new_n691_), .B2(new_n549_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n617_), .A2(new_n694_), .A3(new_n660_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n614_), .A2(new_n503_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n588_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n616_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n577_), .A2(new_n585_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n696_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  OAI211_X1 g500(.A(new_n586_), .B(KEYINPUT105), .C1(new_n615_), .C2(new_n616_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n703_));
  INV_X1    g502(.A(new_n659_), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT37), .B1(new_n640_), .B2(new_n642_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n703_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n658_), .A2(KEYINPUT106), .A3(new_n659_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n701_), .A2(new_n702_), .A3(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n695_), .B1(new_n710_), .B2(KEYINPUT43), .ZN(new_n711_));
  INV_X1    g510(.A(new_n315_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n651_), .A2(new_n288_), .A3(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n693_), .B1(new_n711_), .B2(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n708_), .B1(new_n617_), .B2(new_n696_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n694_), .B1(new_n716_), .B2(new_n702_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n713_), .B(KEYINPUT44), .C1(new_n717_), .C2(new_n695_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n715_), .A2(new_n718_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n549_), .A2(G29gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n692_), .B1(new_n719_), .B2(new_n720_), .ZN(G1328gat));
  INV_X1    g520(.A(new_n581_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n715_), .A2(new_n722_), .A3(new_n718_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G36gat), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n581_), .A2(G36gat), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  OAI21_X1  g525(.A(KEYINPUT45), .B1(new_n690_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT45), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n656_), .A2(new_n728_), .A3(new_n689_), .A4(new_n725_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n724_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT46), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n724_), .A2(new_n730_), .A3(KEYINPUT46), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1329gat));
  NAND4_X1  g534(.A1(new_n715_), .A2(G43gat), .A3(new_n616_), .A4(new_n718_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(KEYINPUT107), .B(G43gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n737_), .B1(new_n690_), .B2(new_n583_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g539(.A(G50gat), .B1(new_n691_), .B2(new_n682_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n682_), .A2(G50gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n719_), .B2(new_n742_), .ZN(G1331gat));
  NAND4_X1  g542(.A1(new_n645_), .A2(new_n288_), .A3(new_n651_), .A4(new_n712_), .ZN(new_n744_));
  INV_X1    g543(.A(G57gat), .ZN(new_n745_));
  NOR3_X1   g544(.A1(new_n744_), .A2(new_n745_), .A3(new_n550_), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n617_), .A2(new_n651_), .A3(new_n712_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(new_n661_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n749_), .A2(KEYINPUT108), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(KEYINPUT108), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(new_n549_), .A3(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n746_), .B1(new_n752_), .B2(new_n745_), .ZN(G1332gat));
  OAI21_X1  g552(.A(G64gat), .B1(new_n744_), .B2(new_n581_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT48), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n581_), .A2(G64gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n755_), .B1(new_n748_), .B2(new_n756_), .ZN(G1333gat));
  OAI21_X1  g556(.A(G71gat), .B1(new_n744_), .B2(new_n583_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT49), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n583_), .A2(G71gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n759_), .B1(new_n748_), .B2(new_n760_), .ZN(G1334gat));
  OAI21_X1  g560(.A(G78gat), .B1(new_n744_), .B2(new_n503_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT50), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n749_), .A2(new_n477_), .A3(new_n682_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(G1335gat));
  NAND2_X1  g564(.A1(new_n712_), .A2(new_n287_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n259_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n767_), .B(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n769_), .B1(new_n717_), .B2(new_n695_), .ZN(new_n770_));
  OAI21_X1  g569(.A(G85gat), .B1(new_n770_), .B2(new_n550_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n747_), .A2(new_n689_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n772_), .A2(G85gat), .A3(new_n550_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n771_), .A2(new_n774_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT110), .ZN(G1336gat));
  OAI21_X1  g575(.A(G92gat), .B1(new_n770_), .B2(new_n581_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n772_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(new_n217_), .A3(new_n722_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(G1337gat));
  XNOR2_X1  g579(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n616_), .B(new_n769_), .C1(new_n717_), .C2(new_n695_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(G99gat), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n782_), .A2(KEYINPUT111), .A3(G99gat), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n747_), .A2(new_n208_), .A3(new_n616_), .A4(new_n689_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT112), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n781_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n782_), .A2(KEYINPUT111), .A3(G99gat), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT111), .B1(new_n782_), .B2(G99gat), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n789_), .B(new_n781_), .C1(new_n791_), .C2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n790_), .A2(new_n794_), .ZN(G1338gat));
  NAND3_X1  g594(.A1(new_n778_), .A2(new_n209_), .A3(new_n682_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n682_), .B(new_n769_), .C1(new_n717_), .C2(new_n695_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n797_), .A2(new_n798_), .A3(G106gat), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n797_), .B2(G106gat), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n796_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT53), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n803_), .B(new_n796_), .C1(new_n799_), .C2(new_n800_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(G1339gat));
  NAND4_X1  g604(.A1(new_n712_), .A2(new_n288_), .A3(new_n256_), .A4(new_n257_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n806_), .A2(new_n660_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT54), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n311_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n305_), .A2(new_n296_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n314_), .A2(new_n250_), .A3(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT56), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n245_), .A2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n237_), .A2(new_n241_), .A3(new_n244_), .ZN(new_n817_));
  AOI22_X1  g616(.A1(new_n816_), .A2(KEYINPUT55), .B1(new_n239_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n245_), .A2(new_n815_), .A3(new_n819_), .ZN(new_n820_));
  AOI211_X1 g619(.A(new_n814_), .B(new_n207_), .C1(new_n818_), .C2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n816_), .A2(KEYINPUT55), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n817_), .A2(new_n239_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n822_), .A2(new_n820_), .A3(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n207_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT56), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n813_), .B(KEYINPUT116), .C1(new_n821_), .C2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT58), .B1(new_n827_), .B2(KEYINPUT117), .ZN(new_n828_));
  AND3_X1   g627(.A1(new_n245_), .A2(new_n815_), .A3(new_n819_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n819_), .B1(new_n245_), .B2(new_n815_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n817_), .A2(new_n239_), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n829_), .A2(new_n830_), .A3(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n814_), .B1(new_n832_), .B2(new_n207_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n824_), .A2(KEYINPUT56), .A3(new_n825_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n812_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n836_), .B1(KEYINPUT117), .B2(KEYINPUT58), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n835_), .A2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n660_), .B1(new_n828_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n840_));
  INV_X1    g639(.A(new_n643_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n252_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(new_n821_), .B2(new_n826_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n252_), .A2(new_n248_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n314_), .A2(new_n811_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n841_), .B1(new_n843_), .B2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n840_), .B1(new_n848_), .B2(KEYINPUT57), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(KEYINPUT57), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n315_), .A2(new_n250_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n851_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n643_), .B1(new_n852_), .B2(new_n846_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(KEYINPUT115), .A3(new_n854_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n839_), .A2(new_n849_), .A3(new_n850_), .A4(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n808_), .B1(new_n856_), .B2(new_n287_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n511_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n550_), .A2(new_n583_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n857_), .A2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(G113gat), .B1(new_n861_), .B2(new_n315_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT59), .B1(new_n857_), .B2(new_n860_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n860_), .A2(KEYINPUT59), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n853_), .A2(new_n854_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n813_), .B1(new_n821_), .B2(new_n826_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n837_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT117), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n869_), .B1(new_n835_), .B2(KEYINPUT116), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n868_), .B1(new_n870_), .B2(KEYINPUT58), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n865_), .B1(new_n871_), .B2(new_n660_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n853_), .A2(new_n854_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n288_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n864_), .B1(new_n874_), .B2(new_n808_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n863_), .A2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n315_), .A2(G113gat), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(KEYINPUT118), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n862_), .B1(new_n876_), .B2(new_n878_), .ZN(G1340gat));
  NAND3_X1  g678(.A1(new_n863_), .A2(new_n875_), .A3(new_n651_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(G120gat), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT60), .ZN(new_n882_));
  AOI21_X1  g681(.A(G120gat), .B1(new_n651_), .B2(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n883_), .B1(new_n882_), .B2(G120gat), .ZN(new_n884_));
  AOI21_X1  g683(.A(KEYINPUT119), .B1(new_n861_), .B2(new_n884_), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n861_), .A2(KEYINPUT119), .A3(new_n884_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n881_), .B1(new_n885_), .B2(new_n886_), .ZN(G1341gat));
  AOI21_X1  g686(.A(G127gat), .B1(new_n861_), .B2(new_n288_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n288_), .A2(G127gat), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(KEYINPUT120), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n888_), .B1(new_n876_), .B2(new_n890_), .ZN(G1342gat));
  NAND3_X1  g690(.A1(new_n863_), .A2(new_n875_), .A3(new_n660_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(G134gat), .ZN(new_n893_));
  INV_X1    g692(.A(G134gat), .ZN(new_n894_));
  INV_X1    g693(.A(new_n644_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n861_), .A2(new_n894_), .A3(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n893_), .A2(new_n896_), .ZN(G1343gat));
  INV_X1    g696(.A(new_n857_), .ZN(new_n898_));
  NOR4_X1   g697(.A1(new_n722_), .A2(new_n550_), .A3(new_n503_), .A4(new_n616_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n898_), .A2(new_n315_), .A3(new_n899_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g700(.A1(new_n898_), .A2(new_n651_), .A3(new_n899_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g702(.A1(new_n898_), .A2(new_n288_), .A3(new_n899_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(KEYINPUT61), .B(G155gat), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n904_), .B(new_n905_), .ZN(G1346gat));
  AND4_X1   g705(.A1(G162gat), .A2(new_n898_), .A3(new_n709_), .A4(new_n899_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n898_), .A2(new_n895_), .A3(new_n899_), .ZN(new_n908_));
  INV_X1    g707(.A(G162gat), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n907_), .B1(new_n908_), .B2(new_n909_), .ZN(G1347gat));
  NAND3_X1  g709(.A1(new_n839_), .A2(new_n873_), .A3(new_n850_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n808_), .B1(new_n911_), .B2(new_n287_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n581_), .A2(new_n576_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n914_), .A2(new_n682_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n912_), .A2(new_n712_), .A3(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n918_));
  INV_X1    g717(.A(G169gat), .ZN(new_n919_));
  OR3_X1    g718(.A1(new_n917_), .A2(new_n918_), .A3(new_n919_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n918_), .B1(new_n917_), .B2(new_n919_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n917_), .A2(new_n368_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n920_), .A2(new_n921_), .A3(new_n922_), .ZN(G1348gat));
  NOR2_X1   g722(.A1(new_n912_), .A2(new_n916_), .ZN(new_n924_));
  AOI21_X1  g723(.A(G176gat), .B1(new_n924_), .B2(new_n651_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n857_), .A2(new_n682_), .ZN(new_n926_));
  NOR3_X1   g725(.A1(new_n259_), .A2(new_n369_), .A3(new_n914_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n925_), .B1(new_n926_), .B2(new_n927_), .ZN(G1349gat));
  NAND3_X1  g727(.A1(new_n926_), .A2(new_n288_), .A3(new_n913_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n287_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n930_));
  AOI22_X1  g729(.A1(new_n929_), .A2(new_n331_), .B1(new_n924_), .B2(new_n930_), .ZN(G1350gat));
  NAND4_X1  g730(.A1(new_n924_), .A2(new_n357_), .A3(new_n358_), .A4(new_n895_), .ZN(new_n932_));
  OAI211_X1 g731(.A(new_n660_), .B(new_n915_), .C1(new_n874_), .C2(new_n808_), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT121), .ZN(new_n934_));
  AND3_X1   g733(.A1(new_n933_), .A2(new_n934_), .A3(G190gat), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n934_), .B1(new_n933_), .B2(G190gat), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n932_), .B1(new_n935_), .B2(new_n936_), .ZN(G1351gat));
  AND2_X1   g736(.A1(new_n587_), .A2(new_n583_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n722_), .A2(new_n938_), .ZN(new_n939_));
  INV_X1    g738(.A(new_n939_), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n898_), .A2(new_n315_), .A3(new_n940_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n325_), .A2(KEYINPUT122), .ZN(new_n942_));
  INV_X1    g741(.A(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n325_), .A2(KEYINPUT122), .ZN(new_n944_));
  XOR2_X1   g743(.A(new_n944_), .B(KEYINPUT123), .Z(new_n945_));
  AND3_X1   g744(.A1(new_n941_), .A2(new_n943_), .A3(new_n945_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n945_), .B1(new_n941_), .B2(new_n943_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n946_), .A2(new_n947_), .ZN(G1352gat));
  NOR2_X1   g747(.A1(new_n857_), .A2(new_n939_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n949_), .A2(new_n651_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g750(.A(new_n287_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n952_), .B(KEYINPUT124), .ZN(new_n953_));
  NOR3_X1   g752(.A1(KEYINPUT125), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n953_), .A2(new_n954_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n949_), .A2(new_n955_), .ZN(new_n956_));
  OAI21_X1  g755(.A(KEYINPUT125), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n957_));
  INV_X1    g756(.A(new_n957_), .ZN(new_n958_));
  XNOR2_X1  g757(.A(new_n956_), .B(new_n958_), .ZN(G1354gat));
  INV_X1    g758(.A(new_n660_), .ZN(new_n960_));
  XOR2_X1   g759(.A(KEYINPUT127), .B(G218gat), .Z(new_n961_));
  NOR4_X1   g760(.A1(new_n857_), .A2(new_n960_), .A3(new_n939_), .A4(new_n961_), .ZN(new_n962_));
  NOR3_X1   g761(.A1(new_n848_), .A2(new_n840_), .A3(KEYINPUT57), .ZN(new_n963_));
  AOI21_X1  g762(.A(KEYINPUT115), .B1(new_n853_), .B2(new_n854_), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n963_), .A2(new_n964_), .ZN(new_n965_));
  AOI21_X1  g764(.A(new_n288_), .B1(new_n872_), .B2(new_n965_), .ZN(new_n966_));
  OAI211_X1 g765(.A(new_n895_), .B(new_n940_), .C1(new_n966_), .C2(new_n808_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n967_), .A2(KEYINPUT126), .ZN(new_n968_));
  INV_X1    g767(.A(KEYINPUT126), .ZN(new_n969_));
  NAND4_X1  g768(.A1(new_n898_), .A2(new_n969_), .A3(new_n895_), .A4(new_n940_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n968_), .A2(new_n970_), .ZN(new_n971_));
  AOI21_X1  g770(.A(new_n962_), .B1(new_n971_), .B2(new_n961_), .ZN(G1355gat));
endmodule


