//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 1 0 0 1 1 1 0 1 1 0 0 1 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0 0 1 1 1 1 0 1 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 0 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n930_,
    new_n932_, new_n933_, new_n935_, new_n936_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n960_, new_n961_, new_n963_, new_n964_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n971_, new_n972_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n979_, new_n980_;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G211gat), .B(G218gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(G197gat), .A2(G204gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G197gat), .A2(G204gat), .ZN(new_n208_));
  NAND4_X1  g007(.A1(new_n205_), .A2(KEYINPUT21), .A3(new_n207_), .A4(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n207_), .A2(KEYINPUT21), .A3(new_n208_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT21), .ZN(new_n211_));
  INV_X1    g010(.A(new_n208_), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n211_), .B1(new_n212_), .B2(new_n206_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n210_), .A2(new_n213_), .A3(new_n204_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n209_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT29), .ZN(new_n216_));
  INV_X1    g015(.A(G141gat), .ZN(new_n217_));
  INV_X1    g016(.A(G148gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT1), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n219_), .B(new_n220_), .C1(new_n221_), .C2(new_n222_), .ZN(new_n223_));
  AND2_X1   g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G155gat), .A2(G162gat), .ZN(new_n225_));
  NOR3_X1   g024(.A1(new_n224_), .A2(new_n225_), .A3(KEYINPUT1), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n223_), .A2(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n224_), .A2(new_n225_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT87), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT2), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n220_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT3), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n232_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n231_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n230_), .B1(new_n220_), .B2(new_n229_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n228_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT88), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n227_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  OAI211_X1 g038(.A(KEYINPUT88), .B(new_n228_), .C1(new_n235_), .C2(new_n236_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n216_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT90), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n215_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  AOI211_X1 g042(.A(KEYINPUT90), .B(new_n216_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n203_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT91), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G78gat), .B(G106gat), .ZN(new_n247_));
  XOR2_X1   g046(.A(new_n247_), .B(KEYINPUT92), .Z(new_n248_));
  INV_X1    g047(.A(KEYINPUT91), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n249_), .B(new_n203_), .C1(new_n243_), .C2(new_n244_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT89), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n209_), .A2(new_n214_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n252_), .A2(new_n203_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n251_), .B1(new_n254_), .B2(new_n241_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n237_), .A2(new_n238_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n227_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(new_n240_), .A3(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT29), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n259_), .A2(KEYINPUT89), .A3(new_n253_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n255_), .A2(new_n260_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n246_), .A2(new_n248_), .A3(new_n250_), .A4(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT93), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n250_), .A2(new_n261_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT93), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n264_), .A2(new_n265_), .A3(new_n248_), .A4(new_n246_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n258_), .A2(KEYINPUT29), .ZN(new_n267_));
  XOR2_X1   g066(.A(new_n267_), .B(KEYINPUT28), .Z(new_n268_));
  XNOR2_X1  g067(.A(G22gat), .B(G50gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n250_), .A2(new_n261_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n252_), .B1(new_n259_), .B2(KEYINPUT90), .ZN(new_n272_));
  INV_X1    g071(.A(new_n244_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n249_), .B1(new_n274_), .B2(new_n203_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n247_), .B1(new_n271_), .B2(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n263_), .A2(new_n266_), .A3(new_n270_), .A4(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n248_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n278_), .B1(new_n271_), .B2(new_n275_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n262_), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n268_), .B(new_n269_), .Z(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n277_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT27), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G8gat), .B(G36gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT18), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G64gat), .B(G92gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT94), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G226gat), .A2(G233gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT19), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G169gat), .A2(G176gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT77), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT77), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(G169gat), .A3(G176gat), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n295_), .A2(new_n297_), .A3(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(G183gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT25), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT25), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(G183gat), .ZN(new_n304_));
  INV_X1    g103(.A(G190gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT26), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT26), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(G190gat), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n302_), .A2(new_n304_), .A3(new_n306_), .A4(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(G169gat), .A2(G176gat), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT24), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G183gat), .A2(G190gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT23), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT23), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n315_), .A2(G183gat), .A3(G190gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n300_), .A2(new_n309_), .A3(new_n312_), .A4(new_n317_), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n297_), .A2(new_n299_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n313_), .A2(new_n315_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n301_), .A2(new_n305_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(G169gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT22), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT22), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(G169gat), .ZN(new_n327_));
  INV_X1    g126(.A(G176gat), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n325_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n319_), .A2(new_n323_), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n318_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT78), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT78), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n318_), .A2(new_n333_), .A3(new_n330_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n332_), .A2(new_n252_), .A3(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT20), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT25), .B(G183gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT26), .B(G190gat), .ZN(new_n338_));
  AOI22_X1  g137(.A1(new_n337_), .A2(new_n338_), .B1(new_n311_), .B2(new_n310_), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n295_), .A2(new_n296_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(new_n330_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n336_), .B1(new_n342_), .B2(new_n215_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n293_), .B1(new_n335_), .B2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT20), .B1(new_n342_), .B2(new_n215_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n332_), .A2(new_n334_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n345_), .B1(new_n346_), .B2(new_n215_), .ZN(new_n347_));
  AOI22_X1  g146(.A1(new_n290_), .A2(new_n344_), .B1(new_n347_), .B2(new_n293_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n335_), .A2(new_n343_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n290_), .B1(new_n349_), .B2(new_n292_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n289_), .B1(new_n348_), .B2(new_n351_), .ZN(new_n352_));
  AND3_X1   g151(.A1(new_n318_), .A2(new_n333_), .A3(new_n330_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n333_), .B1(new_n318_), .B2(new_n330_), .ZN(new_n354_));
  NOR3_X1   g153(.A1(new_n353_), .A2(new_n354_), .A3(new_n215_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n319_), .A2(new_n329_), .ZN(new_n356_));
  AOI22_X1  g155(.A1(new_n356_), .A2(new_n323_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT20), .B1(new_n357_), .B2(new_n252_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n290_), .B(new_n292_), .C1(new_n355_), .C2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n215_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n336_), .B1(new_n357_), .B2(new_n252_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(new_n361_), .A3(new_n293_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n359_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n289_), .ZN(new_n364_));
  NOR3_X1   g163(.A1(new_n363_), .A2(new_n364_), .A3(new_n350_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n284_), .B1(new_n352_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT98), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT97), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n289_), .B(KEYINPUT96), .ZN(new_n369_));
  NOR3_X1   g168(.A1(new_n355_), .A2(new_n358_), .A3(new_n292_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n293_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n369_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT27), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n368_), .B1(new_n365_), .B2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n348_), .A2(new_n351_), .A3(new_n289_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n335_), .A2(new_n293_), .A3(new_n343_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n376_), .B1(new_n347_), .B2(new_n293_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n284_), .B1(new_n377_), .B2(new_n369_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n375_), .A2(KEYINPUT97), .A3(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n374_), .A2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n364_), .B1(new_n363_), .B2(new_n350_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n375_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT98), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(new_n383_), .A3(new_n284_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n367_), .A2(new_n380_), .A3(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G225gat), .A2(G233gat), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(G127gat), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n388_), .A2(G134gat), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n388_), .A2(G134gat), .ZN(new_n390_));
  INV_X1    g189(.A(G113gat), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n391_), .A2(G120gat), .ZN(new_n392_));
  INV_X1    g191(.A(G120gat), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n393_), .A2(G113gat), .ZN(new_n394_));
  OAI22_X1  g193(.A1(new_n389_), .A2(new_n390_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G127gat), .B(G134gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G113gat), .B(G120gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n395_), .A2(KEYINPUT84), .A3(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(KEYINPUT84), .B1(new_n395_), .B2(new_n398_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n258_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n395_), .A2(new_n398_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n239_), .A2(new_n240_), .A3(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n387_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(KEYINPUT4), .B1(new_n258_), .B2(new_n401_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n402_), .A2(new_n404_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n406_), .B1(new_n407_), .B2(KEYINPUT4), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n405_), .B1(new_n408_), .B2(new_n387_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G1gat), .B(G29gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(G85gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT0), .B(G57gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n409_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n413_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n416_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n417_));
  NOR3_X1   g216(.A1(new_n417_), .A2(new_n386_), .A3(new_n406_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n415_), .B1(new_n418_), .B2(new_n405_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n414_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT80), .B(KEYINPUT82), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT79), .B(KEYINPUT30), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n332_), .A2(new_n334_), .A3(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n423_), .B1(new_n332_), .B2(new_n334_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n422_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n423_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n346_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n422_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n429_), .A2(new_n424_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n427_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G227gat), .A2(G233gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT81), .ZN(new_n434_));
  XOR2_X1   g233(.A(G71gat), .B(G99gat), .Z(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G15gat), .B(G43gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n432_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT84), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n396_), .A2(new_n397_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n396_), .A2(new_n397_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n440_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n395_), .A2(new_n398_), .A3(KEYINPUT84), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(KEYINPUT31), .ZN(new_n446_));
  AOI21_X1  g245(.A(KEYINPUT85), .B1(new_n446_), .B2(KEYINPUT83), .ZN(new_n447_));
  INV_X1    g246(.A(new_n438_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n427_), .A2(new_n448_), .A3(new_n431_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n439_), .A2(new_n447_), .A3(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n447_), .B1(KEYINPUT85), .B2(new_n446_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n449_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n448_), .B1(new_n427_), .B2(new_n431_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n451_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n421_), .A2(new_n450_), .A3(new_n454_), .ZN(new_n455_));
  NOR3_X1   g254(.A1(new_n283_), .A2(new_n385_), .A3(new_n455_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n367_), .A2(new_n380_), .A3(new_n421_), .A4(new_n384_), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n457_), .A2(new_n283_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT86), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n454_), .A2(new_n459_), .A3(new_n450_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n459_), .B1(new_n454_), .B2(new_n450_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n377_), .A2(KEYINPUT32), .A3(new_n289_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n289_), .A2(KEYINPUT32), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n348_), .A2(new_n351_), .A3(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n420_), .A2(new_n463_), .A3(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n402_), .A2(new_n404_), .A3(new_n387_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(new_n413_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT95), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n445_), .B1(new_n240_), .B2(new_n239_), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n239_), .A2(new_n240_), .A3(new_n403_), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT4), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n406_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n470_), .B1(new_n475_), .B2(new_n386_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n470_), .B(new_n386_), .C1(new_n417_), .C2(new_n406_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n469_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n479_), .A2(new_n375_), .A3(new_n381_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT33), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n419_), .A2(new_n481_), .ZN(new_n482_));
  OAI211_X1 g281(.A(KEYINPUT33), .B(new_n415_), .C1(new_n418_), .C2(new_n405_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n466_), .B1(new_n480_), .B2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n462_), .B1(new_n283_), .B2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT99), .B1(new_n458_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n457_), .A2(new_n283_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n484_), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT95), .B1(new_n408_), .B2(new_n387_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n468_), .B1(new_n490_), .B2(new_n477_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n382_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n489_), .A2(new_n492_), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n493_), .A2(new_n282_), .A3(new_n277_), .A4(new_n466_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT99), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n488_), .A2(new_n494_), .A3(new_n495_), .A4(new_n462_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n456_), .B1(new_n487_), .B2(new_n496_), .ZN(new_n497_));
  XOR2_X1   g296(.A(G29gat), .B(G36gat), .Z(new_n498_));
  XOR2_X1   g297(.A(G43gat), .B(G50gat), .Z(new_n499_));
  OR2_X1    g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n499_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT75), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G15gat), .B(G22gat), .ZN(new_n505_));
  INV_X1    g304(.A(G1gat), .ZN(new_n506_));
  INV_X1    g305(.A(G8gat), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT14), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n505_), .A2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G1gat), .B(G8gat), .ZN(new_n510_));
  XOR2_X1   g309(.A(new_n509_), .B(new_n510_), .Z(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n504_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n503_), .A2(new_n511_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n513_), .A2(new_n514_), .A3(KEYINPUT76), .ZN(new_n515_));
  OR3_X1    g314(.A1(new_n503_), .A2(KEYINPUT76), .A3(new_n511_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G229gat), .A2(G233gat), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n502_), .B(KEYINPUT15), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(new_n512_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n514_), .A2(new_n523_), .A3(new_n519_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n521_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G113gat), .B(G141gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G169gat), .B(G197gat), .ZN(new_n527_));
  XOR2_X1   g326(.A(new_n526_), .B(new_n527_), .Z(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n525_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n521_), .A2(new_n524_), .A3(new_n528_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n497_), .A2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G120gat), .B(G148gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT5), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G176gat), .B(G204gat), .ZN(new_n537_));
  XOR2_X1   g336(.A(new_n536_), .B(new_n537_), .Z(new_n538_));
  XNOR2_X1  g337(.A(G57gat), .B(G64gat), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT70), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT11), .ZN(new_n542_));
  XOR2_X1   g341(.A(G71gat), .B(G78gat), .Z(new_n543_));
  OR2_X1    g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n539_), .B(KEYINPUT70), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT11), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n542_), .A2(new_n547_), .A3(new_n543_), .ZN(new_n548_));
  AND2_X1   g347(.A1(new_n544_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(KEYINPUT66), .B(KEYINPUT6), .ZN(new_n550_));
  INV_X1    g349(.A(G99gat), .ZN(new_n551_));
  INV_X1    g350(.A(G106gat), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n550_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n551_), .A2(new_n552_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n550_), .A2(new_n553_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(KEYINPUT67), .A2(KEYINPUT7), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n554_), .A2(new_n557_), .A3(new_n558_), .A4(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT69), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G85gat), .B(G92gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT68), .ZN(new_n563_));
  AND3_X1   g362(.A1(new_n560_), .A2(new_n561_), .A3(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n561_), .B1(new_n560_), .B2(new_n563_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT8), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n564_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n560_), .A2(new_n563_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n568_), .A2(KEYINPUT69), .A3(new_n566_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n554_), .A2(new_n558_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT9), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n571_), .A2(G85gat), .A3(G92gat), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n572_), .B1(new_n562_), .B2(new_n571_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n570_), .A2(new_n573_), .ZN(new_n574_));
  OR2_X1    g373(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n575_));
  NAND2_X1  g374(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT64), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n575_), .A2(KEYINPUT64), .A3(new_n576_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n581_), .A2(KEYINPUT65), .A3(new_n552_), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT65), .B1(new_n581_), .B2(new_n552_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n574_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n569_), .A2(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n549_), .B1(new_n567_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n568_), .A2(KEYINPUT69), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n560_), .A2(new_n561_), .A3(new_n563_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(KEYINPUT8), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n544_), .A2(new_n548_), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n589_), .A2(new_n590_), .A3(new_n569_), .A4(new_n584_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n586_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G230gat), .A2(G233gat), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT71), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n592_), .A2(KEYINPUT71), .A3(new_n594_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n586_), .A2(KEYINPUT12), .A3(new_n591_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n569_), .A2(new_n584_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(new_n589_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT12), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n602_), .A2(new_n603_), .A3(new_n549_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n594_), .B1(new_n600_), .B2(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n538_), .B1(new_n599_), .B2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n600_), .A2(new_n604_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(new_n593_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n538_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n608_), .A2(new_n597_), .A3(new_n598_), .A4(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT13), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT72), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(KEYINPUT72), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  AOI22_X1  g413(.A1(new_n606_), .A2(new_n610_), .B1(new_n612_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n606_), .A2(new_n610_), .A3(new_n614_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT37), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n602_), .A2(new_n522_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n502_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n620_), .B1(new_n621_), .B2(new_n602_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G232gat), .A2(G233gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT34), .ZN(new_n624_));
  INV_X1    g423(.A(new_n522_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n625_), .B1(new_n601_), .B2(new_n589_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT73), .ZN(new_n627_));
  OAI211_X1 g426(.A(KEYINPUT35), .B(new_n624_), .C1(new_n626_), .C2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G190gat), .B(G218gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G134gat), .B(G162gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  AOI22_X1  g430(.A1(new_n622_), .A2(new_n628_), .B1(KEYINPUT36), .B2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n602_), .A2(new_n621_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n633_), .A2(new_n626_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n624_), .A2(KEYINPUT35), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n620_), .B2(KEYINPUT73), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n624_), .A2(KEYINPUT35), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n634_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n631_), .A2(KEYINPUT36), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n632_), .A2(new_n638_), .A3(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n640_), .B1(new_n632_), .B2(new_n638_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n619_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n632_), .A2(new_n638_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(new_n639_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n632_), .A2(new_n638_), .A3(new_n640_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n645_), .A2(KEYINPUT37), .A3(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n590_), .B(new_n511_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(G231gat), .A2(G233gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n648_), .B(new_n649_), .ZN(new_n650_));
  XOR2_X1   g449(.A(G127gat), .B(G155gat), .Z(new_n651_));
  XNOR2_X1  g450(.A(G183gat), .B(G211gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(new_n653_));
  XOR2_X1   g452(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n650_), .A2(KEYINPUT17), .A3(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n655_), .B(KEYINPUT17), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n650_), .A2(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n643_), .A2(new_n647_), .A3(new_n659_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n534_), .A2(new_n618_), .A3(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n661_), .A2(new_n506_), .A3(new_n420_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT100), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT38), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n664_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT101), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n618_), .A2(new_n667_), .A3(new_n532_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n617_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n532_), .B1(new_n670_), .B2(new_n615_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT101), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n659_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n669_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n645_), .A2(new_n646_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n497_), .A2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n675_), .A2(new_n420_), .A3(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(G1gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n665_), .A2(new_n666_), .A3(new_n680_), .ZN(G1324gat));
  NAND3_X1  g480(.A1(new_n661_), .A2(new_n507_), .A3(new_n385_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n675_), .A2(new_n385_), .A3(new_n678_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT39), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n683_), .A2(new_n684_), .A3(G8gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n683_), .B2(G8gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n682_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  XOR2_X1   g486(.A(KEYINPUT102), .B(KEYINPUT40), .Z(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(G1325gat));
  INV_X1    g488(.A(new_n461_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n454_), .A2(new_n459_), .A3(new_n450_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n675_), .A2(new_n692_), .A3(new_n678_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n693_), .A2(new_n694_), .A3(G15gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n693_), .B2(G15gat), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT41), .ZN(new_n697_));
  OR3_X1    g496(.A1(new_n695_), .A2(new_n696_), .A3(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n697_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n699_));
  INV_X1    g498(.A(G15gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n661_), .A2(new_n700_), .A3(new_n692_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n698_), .A2(new_n699_), .A3(new_n701_), .ZN(G1326gat));
  AND2_X1   g501(.A1(new_n277_), .A2(new_n282_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT104), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n704_), .A2(G22gat), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT105), .Z(new_n706_));
  NAND2_X1  g505(.A1(new_n661_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n704_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n675_), .A2(new_n678_), .A3(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(G22gat), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n710_), .A2(KEYINPUT42), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(KEYINPUT42), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n707_), .B1(new_n711_), .B2(new_n712_), .ZN(G1327gat));
  NOR2_X1   g512(.A1(new_n676_), .A2(new_n659_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n618_), .A2(new_n714_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n534_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(G29gat), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n420_), .A2(new_n717_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT107), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n716_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT106), .ZN(new_n721_));
  INV_X1    g520(.A(new_n456_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n485_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n692_), .B1(new_n703_), .B2(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n495_), .B1(new_n724_), .B2(new_n488_), .ZN(new_n725_));
  AND4_X1   g524(.A1(new_n495_), .A2(new_n488_), .A3(new_n494_), .A4(new_n462_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n722_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT43), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n643_), .A2(new_n647_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n727_), .A2(new_n728_), .A3(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n729_), .ZN(new_n731_));
  OAI21_X1  g530(.A(KEYINPUT43), .B1(new_n497_), .B2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n668_), .A2(new_n672_), .A3(new_n674_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(KEYINPUT44), .B1(new_n733_), .B2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n737_));
  AOI211_X1 g536(.A(new_n737_), .B(new_n734_), .C1(new_n730_), .C2(new_n732_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n736_), .A2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n420_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n721_), .B1(new_n740_), .B2(G29gat), .ZN(new_n741_));
  AOI211_X1 g540(.A(KEYINPUT106), .B(new_n717_), .C1(new_n739_), .C2(new_n420_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n720_), .B1(new_n741_), .B2(new_n742_), .ZN(G1328gat));
  XNOR2_X1  g542(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n744_));
  INV_X1    g543(.A(G36gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n739_), .B2(new_n385_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n534_), .A2(new_n745_), .A3(new_n385_), .A4(new_n715_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT45), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n747_), .B(new_n748_), .ZN(new_n749_));
  OAI211_X1 g548(.A(KEYINPUT108), .B(new_n744_), .C1(new_n746_), .C2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n744_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n728_), .B1(new_n727_), .B2(new_n729_), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n497_), .A2(KEYINPUT43), .A3(new_n731_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n735_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(new_n737_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n733_), .A2(KEYINPUT44), .A3(new_n735_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n755_), .A2(new_n385_), .A3(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n749_), .B1(new_n757_), .B2(G36gat), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n751_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n750_), .A2(new_n760_), .ZN(G1329gat));
  AOI21_X1  g560(.A(G43gat), .B1(new_n716_), .B2(new_n692_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n454_), .A2(G43gat), .A3(new_n450_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n739_), .B2(new_n763_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT47), .Z(G1330gat));
  NOR2_X1   g564(.A1(new_n704_), .A2(G50gat), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT110), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n716_), .A2(new_n767_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n736_), .A2(new_n738_), .A3(new_n703_), .ZN(new_n769_));
  INV_X1    g568(.A(G50gat), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n768_), .B1(new_n769_), .B2(new_n770_), .ZN(G1331gat));
  NOR3_X1   g570(.A1(new_n618_), .A2(new_n532_), .A3(new_n674_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n678_), .A2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(G57gat), .B1(new_n773_), .B2(new_n421_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n618_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n660_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT111), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n497_), .A2(new_n532_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  OR2_X1    g578(.A1(new_n421_), .A2(G57gat), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n774_), .B1(new_n779_), .B2(new_n780_), .ZN(G1332gat));
  INV_X1    g580(.A(new_n385_), .ZN(new_n782_));
  OR3_X1    g581(.A1(new_n779_), .A2(G64gat), .A3(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n678_), .A2(new_n385_), .A3(new_n772_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n784_), .A2(G64gat), .ZN(new_n785_));
  XNOR2_X1  g584(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n785_), .A2(new_n786_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n783_), .B1(new_n787_), .B2(new_n788_), .ZN(G1333gat));
  OAI21_X1  g588(.A(G71gat), .B1(new_n773_), .B2(new_n462_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT49), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n462_), .A2(G71gat), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n791_), .B1(new_n779_), .B2(new_n792_), .ZN(G1334gat));
  OAI21_X1  g592(.A(G78gat), .B1(new_n773_), .B2(new_n704_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT50), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n704_), .A2(G78gat), .ZN(new_n796_));
  XOR2_X1   g595(.A(new_n796_), .B(KEYINPUT113), .Z(new_n797_));
  OAI21_X1  g596(.A(new_n795_), .B1(new_n779_), .B2(new_n797_), .ZN(G1335gat));
  NAND2_X1  g597(.A1(new_n533_), .A2(new_n674_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n618_), .A2(new_n799_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n733_), .A2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n420_), .A2(G85gat), .ZN(new_n802_));
  XOR2_X1   g601(.A(new_n802_), .B(KEYINPUT115), .Z(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n778_), .A2(new_n775_), .A3(new_n714_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n806_));
  OR2_X1    g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n806_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n421_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n804_), .B1(new_n809_), .B2(G85gat), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT116), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n810_), .B(new_n811_), .ZN(G1336gat));
  INV_X1    g611(.A(G92gat), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n807_), .A2(new_n808_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n813_), .B1(new_n815_), .B2(new_n782_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT117), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT117), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n818_), .B(new_n813_), .C1(new_n815_), .C2(new_n782_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n782_), .A2(new_n813_), .ZN(new_n820_));
  AOI22_X1  g619(.A1(new_n817_), .A2(new_n819_), .B1(new_n801_), .B2(new_n820_), .ZN(G1337gat));
  NAND3_X1  g620(.A1(new_n454_), .A2(new_n450_), .A3(new_n581_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n815_), .A2(new_n822_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n801_), .A2(new_n692_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n824_), .A2(new_n551_), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT51), .B1(new_n823_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT51), .ZN(new_n827_));
  OAI221_X1 g626(.A(new_n827_), .B1(new_n824_), .B2(new_n551_), .C1(new_n815_), .C2(new_n822_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(G1338gat));
  NAND3_X1  g628(.A1(new_n814_), .A2(new_n552_), .A3(new_n283_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT52), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n733_), .A2(new_n283_), .A3(new_n800_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(G106gat), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n832_), .A2(new_n831_), .A3(G106gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n830_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT53), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n830_), .B(new_n837_), .C1(new_n833_), .C2(new_n834_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(G1339gat));
  NAND3_X1  g638(.A1(new_n660_), .A2(new_n533_), .A3(new_n618_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n840_), .B(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT57), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n517_), .A2(new_n520_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n514_), .A2(new_n523_), .A3(new_n520_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n529_), .ZN(new_n846_));
  OR3_X1    g645(.A1(new_n844_), .A2(KEYINPUT120), .A3(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT120), .B1(new_n844_), .B2(new_n846_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(new_n531_), .A3(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n849_), .B1(new_n606_), .B2(new_n610_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT56), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n600_), .A2(new_n594_), .A3(new_n604_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT55), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n852_), .A2(new_n605_), .A3(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n607_), .A2(new_n853_), .A3(new_n593_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n538_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n851_), .B1(new_n854_), .B2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(KEYINPUT118), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n600_), .A2(new_n604_), .A3(new_n594_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n608_), .A2(KEYINPUT55), .A3(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n609_), .B1(new_n605_), .B2(new_n853_), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT56), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n860_), .A2(KEYINPUT56), .A3(new_n861_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT119), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n860_), .A2(new_n861_), .A3(new_n867_), .A4(KEYINPUT56), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n858_), .A2(new_n864_), .A3(new_n866_), .A4(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n532_), .A2(new_n610_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n850_), .B1(new_n869_), .B2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n843_), .B1(new_n872_), .B2(new_n677_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n866_), .A2(new_n868_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n860_), .A2(new_n861_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n863_), .B1(new_n875_), .B2(new_n851_), .ZN(new_n876_));
  AOI211_X1 g675(.A(KEYINPUT118), .B(KEYINPUT56), .C1(new_n860_), .C2(new_n861_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n870_), .B1(new_n874_), .B2(new_n878_), .ZN(new_n879_));
  OAI211_X1 g678(.A(KEYINPUT57), .B(new_n676_), .C1(new_n879_), .C2(new_n850_), .ZN(new_n880_));
  AND4_X1   g679(.A1(new_n531_), .A2(new_n847_), .A3(new_n610_), .A4(new_n848_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n865_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n862_), .B2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT58), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n881_), .B(KEYINPUT58), .C1(new_n862_), .C2(new_n882_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n885_), .A2(new_n729_), .A3(new_n886_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n873_), .A2(new_n880_), .A3(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n842_), .B1(new_n888_), .B2(new_n674_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n454_), .A2(new_n450_), .ZN(new_n890_));
  NOR4_X1   g689(.A1(new_n283_), .A2(new_n385_), .A3(new_n421_), .A4(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n889_), .A2(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(G113gat), .B1(new_n893_), .B2(new_n532_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT121), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n888_), .A2(new_n674_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n842_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(KEYINPUT59), .B1(new_n898_), .B2(new_n891_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n889_), .A2(new_n900_), .A3(new_n892_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n895_), .B1(new_n899_), .B2(new_n901_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n898_), .A2(KEYINPUT59), .A3(new_n891_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n900_), .B1(new_n889_), .B2(new_n892_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n903_), .A2(new_n904_), .A3(KEYINPUT121), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n902_), .A2(new_n905_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n391_), .B1(new_n532_), .B2(KEYINPUT122), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n907_), .B1(KEYINPUT122), .B2(new_n391_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n894_), .B1(new_n906_), .B2(new_n908_), .ZN(G1340gat));
  OAI21_X1  g708(.A(new_n393_), .B1(new_n618_), .B2(KEYINPUT60), .ZN(new_n910_));
  OAI211_X1 g709(.A(new_n893_), .B(new_n910_), .C1(KEYINPUT60), .C2(new_n393_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n618_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT123), .ZN(new_n913_));
  OAI21_X1  g712(.A(G120gat), .B1(new_n912_), .B2(new_n913_), .ZN(new_n914_));
  AOI211_X1 g713(.A(KEYINPUT123), .B(new_n618_), .C1(new_n903_), .C2(new_n904_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n911_), .B1(new_n914_), .B2(new_n915_), .ZN(G1341gat));
  NAND3_X1  g715(.A1(new_n893_), .A2(new_n388_), .A3(new_n659_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n674_), .B1(new_n902_), .B2(new_n905_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n918_), .B2(new_n388_), .ZN(G1342gat));
  AOI21_X1  g718(.A(G134gat), .B1(new_n893_), .B2(new_n677_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(KEYINPUT124), .B(G134gat), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n731_), .A2(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n920_), .B1(new_n906_), .B2(new_n922_), .ZN(G1343gat));
  NOR2_X1   g722(.A1(new_n703_), .A2(new_n692_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n924_), .A2(new_n420_), .A3(new_n782_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(KEYINPUT125), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n898_), .A2(new_n926_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n927_), .A2(new_n533_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(new_n217_), .ZN(G1344gat));
  NOR2_X1   g728(.A1(new_n927_), .A2(new_n618_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(new_n218_), .ZN(G1345gat));
  NOR2_X1   g730(.A1(new_n927_), .A2(new_n674_), .ZN(new_n932_));
  XOR2_X1   g731(.A(KEYINPUT61), .B(G155gat), .Z(new_n933_));
  XNOR2_X1  g732(.A(new_n932_), .B(new_n933_), .ZN(G1346gat));
  OAI21_X1  g733(.A(G162gat), .B1(new_n927_), .B2(new_n731_), .ZN(new_n935_));
  OR2_X1    g734(.A1(new_n676_), .A2(G162gat), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n935_), .B1(new_n927_), .B2(new_n936_), .ZN(G1347gat));
  INV_X1    g736(.A(KEYINPUT126), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n782_), .A2(new_n420_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(new_n692_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n708_), .A2(new_n940_), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n898_), .A2(new_n532_), .A3(new_n941_), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n942_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n943_));
  AND2_X1   g742(.A1(new_n325_), .A2(new_n327_), .ZN(new_n944_));
  NAND4_X1  g743(.A1(new_n898_), .A2(new_n944_), .A3(new_n532_), .A4(new_n941_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n943_), .A2(new_n945_), .ZN(new_n946_));
  AOI21_X1  g745(.A(KEYINPUT62), .B1(new_n942_), .B2(G169gat), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n938_), .B1(new_n946_), .B2(new_n947_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n942_), .A2(G169gat), .ZN(new_n949_));
  INV_X1    g748(.A(KEYINPUT62), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n949_), .A2(new_n950_), .ZN(new_n951_));
  NAND4_X1  g750(.A1(new_n951_), .A2(KEYINPUT126), .A3(new_n945_), .A4(new_n943_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n948_), .A2(new_n952_), .ZN(G1348gat));
  NAND2_X1  g752(.A1(new_n898_), .A2(new_n941_), .ZN(new_n954_));
  INV_X1    g753(.A(new_n954_), .ZN(new_n955_));
  AOI21_X1  g754(.A(G176gat), .B1(new_n955_), .B2(new_n775_), .ZN(new_n956_));
  NOR2_X1   g755(.A1(new_n889_), .A2(new_n283_), .ZN(new_n957_));
  NOR3_X1   g756(.A1(new_n940_), .A2(new_n618_), .A3(new_n328_), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n956_), .B1(new_n957_), .B2(new_n958_), .ZN(G1349gat));
  NOR3_X1   g758(.A1(new_n954_), .A2(new_n337_), .A3(new_n674_), .ZN(new_n960_));
  NAND4_X1  g759(.A1(new_n957_), .A2(new_n692_), .A3(new_n659_), .A4(new_n939_), .ZN(new_n961_));
  AOI21_X1  g760(.A(new_n960_), .B1(new_n301_), .B2(new_n961_), .ZN(G1350gat));
  OAI21_X1  g761(.A(G190gat), .B1(new_n954_), .B2(new_n731_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n677_), .A2(new_n338_), .ZN(new_n964_));
  OAI21_X1  g763(.A(new_n963_), .B1(new_n954_), .B2(new_n964_), .ZN(G1351gat));
  AND2_X1   g764(.A1(new_n939_), .A2(new_n924_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n898_), .A2(new_n966_), .ZN(new_n967_));
  NOR2_X1   g766(.A1(new_n967_), .A2(new_n533_), .ZN(new_n968_));
  XOR2_X1   g767(.A(KEYINPUT127), .B(G197gat), .Z(new_n969_));
  XNOR2_X1  g768(.A(new_n968_), .B(new_n969_), .ZN(G1352gat));
  INV_X1    g769(.A(new_n967_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n971_), .A2(new_n775_), .ZN(new_n972_));
  XNOR2_X1  g771(.A(new_n972_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g772(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n974_));
  AND2_X1   g773(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n975_));
  NOR4_X1   g774(.A1(new_n967_), .A2(new_n674_), .A3(new_n974_), .A4(new_n975_), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n971_), .A2(new_n659_), .ZN(new_n977_));
  AOI21_X1  g776(.A(new_n976_), .B1(new_n977_), .B2(new_n974_), .ZN(G1354gat));
  OR3_X1    g777(.A1(new_n967_), .A2(G218gat), .A3(new_n676_), .ZN(new_n979_));
  OAI21_X1  g778(.A(G218gat), .B1(new_n967_), .B2(new_n731_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n979_), .A2(new_n980_), .ZN(G1355gat));
endmodule


