//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 0 1 0 0 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 0 0 0 0 0 1 1 0 0 1 0 1 0 1 1 1 0 1 0 0 1 0 1 1 1 0 1 0 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n795_, new_n796_,
    new_n797_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n902_, new_n903_, new_n904_, new_n906_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n933_, new_n934_, new_n936_,
    new_n937_, new_n938_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n955_, new_n956_, new_n957_;
  INV_X1    g000(.A(KEYINPUT6), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT67), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT67), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT6), .ZN(new_n205_));
  AND2_X1   g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  AND3_X1   g005(.A1(new_n203_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n206_), .B1(new_n203_), .B2(new_n205_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  XOR2_X1   g008(.A(KEYINPUT10), .B(G99gat), .Z(new_n210_));
  INV_X1    g009(.A(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G85gat), .A2(G92gat), .ZN(new_n215_));
  XOR2_X1   g014(.A(G85gat), .B(G92gat), .Z(new_n216_));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(new_n217_), .A3(KEYINPUT9), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT9), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G85gat), .B(G92gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n219_), .B1(new_n220_), .B2(KEYINPUT65), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n215_), .B1(new_n218_), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT66), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n222_), .A2(KEYINPUT66), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n209_), .B(new_n214_), .C1(new_n224_), .C2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G99gat), .A2(G106gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT7), .ZN(new_n228_));
  AOI211_X1 g027(.A(KEYINPUT8), .B(new_n220_), .C1(new_n209_), .C2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT8), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT68), .B1(new_n207_), .B2(new_n208_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n206_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n204_), .A2(KEYINPUT6), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n202_), .A2(KEYINPUT67), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n233_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n203_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n232_), .A2(new_n239_), .A3(new_n228_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n231_), .B1(new_n240_), .B2(new_n216_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n230_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  AOI211_X1 g042(.A(KEYINPUT69), .B(new_n231_), .C1(new_n240_), .C2(new_n216_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n226_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G57gat), .B(G64gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT11), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G71gat), .B(G78gat), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n247_), .A2(new_n249_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n246_), .A2(KEYINPUT11), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n251_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n245_), .A2(new_n255_), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n226_), .B(new_n254_), .C1(new_n243_), .C2(new_n244_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(G230gat), .A3(G233gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT70), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G230gat), .A2(G233gat), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n257_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT12), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n245_), .A2(new_n263_), .A3(new_n255_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n263_), .B1(new_n245_), .B2(new_n255_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n262_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n260_), .B1(new_n257_), .B2(new_n261_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n259_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(KEYINPUT71), .B(KEYINPUT5), .Z(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT72), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G120gat), .B(G148gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G176gat), .B(G204gat), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n272_), .B(new_n273_), .Z(new_n274_));
  NAND2_X1  g073(.A1(new_n268_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT73), .ZN(new_n276_));
  INV_X1    g075(.A(new_n274_), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n259_), .B(new_n277_), .C1(new_n266_), .C2(new_n267_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n275_), .A2(new_n276_), .A3(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n268_), .A2(KEYINPUT73), .A3(new_n274_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT74), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT13), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(KEYINPUT74), .A2(KEYINPUT13), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n281_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n279_), .A2(new_n282_), .A3(new_n283_), .A4(new_n280_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G15gat), .B(G22gat), .ZN(new_n289_));
  INV_X1    g088(.A(G1gat), .ZN(new_n290_));
  INV_X1    g089(.A(G8gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT14), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G1gat), .B(G8gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G231gat), .A2(G233gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(new_n255_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G127gat), .B(G155gat), .Z(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT16), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G183gat), .B(G211gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(KEYINPUT79), .A2(KEYINPUT17), .ZN(new_n304_));
  OR3_X1    g103(.A1(new_n299_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  MUX2_X1   g104(.A(new_n304_), .B(KEYINPUT17), .S(new_n303_), .Z(new_n306_));
  NAND2_X1  g105(.A1(new_n299_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT37), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G190gat), .B(G218gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G134gat), .B(G162gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n312_), .B(KEYINPUT36), .Z(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(G29gat), .B(G36gat), .Z(new_n315_));
  XOR2_X1   g114(.A(G43gat), .B(G50gat), .Z(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT15), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n245_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT75), .B(KEYINPUT34), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G232gat), .A2(G233gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT35), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n226_), .B(new_n317_), .C1(new_n243_), .C2(new_n244_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n319_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n322_), .A2(new_n323_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n327_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n319_), .A2(new_n329_), .A3(new_n324_), .A4(new_n325_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n314_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT78), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(KEYINPUT76), .B(KEYINPUT36), .Z(new_n335_));
  NOR2_X1   g134(.A1(new_n312_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n328_), .A2(new_n330_), .A3(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n337_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n309_), .B1(new_n334_), .B2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n328_), .A2(new_n330_), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n313_), .B(KEYINPUT77), .Z(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(KEYINPUT37), .A3(new_n337_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n339_), .A2(new_n343_), .ZN(new_n344_));
  NOR3_X1   g143(.A1(new_n288_), .A2(new_n308_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n317_), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n346_), .A2(new_n295_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G229gat), .A2(G233gat), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n318_), .A2(new_n295_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n346_), .B(new_n295_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n348_), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n349_), .A2(new_n350_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G113gat), .B(G141gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT80), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G169gat), .B(G197gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n353_), .B(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G8gat), .B(G36gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT18), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G64gat), .B(G92gat), .ZN(new_n362_));
  XOR2_X1   g161(.A(new_n361_), .B(new_n362_), .Z(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G226gat), .A2(G233gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n367_), .B(KEYINPUT99), .Z(new_n368_));
  XOR2_X1   g167(.A(KEYINPUT22), .B(G169gat), .Z(new_n369_));
  INV_X1    g168(.A(KEYINPUT101), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(G176gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(KEYINPUT22), .B(G169gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT101), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n371_), .A2(new_n372_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G169gat), .A2(G176gat), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT83), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT23), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n379_), .B1(G183gat), .B2(G190gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G183gat), .A2(G190gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT84), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT84), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n383_), .A2(G183gat), .A3(G190gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n380_), .B1(new_n385_), .B2(new_n379_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(G183gat), .A2(G190gat), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n375_), .B(new_n378_), .C1(new_n386_), .C2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n379_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n381_), .A2(new_n379_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  NOR3_X1   g191(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n393_), .B1(new_n395_), .B2(new_n376_), .ZN(new_n396_));
  XOR2_X1   g195(.A(KEYINPUT25), .B(G183gat), .Z(new_n397_));
  INV_X1    g196(.A(G190gat), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n398_), .A2(KEYINPUT26), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(KEYINPUT26), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n392_), .B(new_n396_), .C1(new_n397_), .C2(new_n401_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n388_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT21), .ZN(new_n404_));
  INV_X1    g203(.A(G204gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(G197gat), .ZN(new_n406_));
  INV_X1    g205(.A(G197gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(G204gat), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n404_), .B1(new_n406_), .B2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT93), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n406_), .A2(KEYINPUT94), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT94), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n412_), .A2(new_n405_), .A3(G197gat), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n411_), .A2(new_n413_), .A3(new_n404_), .A4(new_n408_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G211gat), .B(G218gat), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n411_), .A2(new_n408_), .A3(new_n413_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n415_), .A2(new_n404_), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n410_), .A2(new_n416_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n403_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT20), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT85), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n373_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(G169gat), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n424_), .A2(KEYINPUT22), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n372_), .B1(new_n425_), .B2(KEYINPUT85), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n378_), .B1(new_n423_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n385_), .A2(KEYINPUT23), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT81), .B(G183gat), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n428_), .B(new_n390_), .C1(G190gat), .C2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT86), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n427_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n429_), .A2(G190gat), .ZN(new_n433_));
  NOR3_X1   g232(.A1(new_n433_), .A2(new_n389_), .A3(new_n391_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT86), .ZN(new_n435_));
  OR2_X1    g234(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n436_));
  XOR2_X1   g235(.A(KEYINPUT81), .B(G183gat), .Z(new_n437_));
  INV_X1    g236(.A(KEYINPUT25), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n436_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n400_), .A2(KEYINPUT82), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n400_), .A2(KEYINPUT82), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n439_), .A2(new_n440_), .A3(new_n399_), .A4(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n376_), .B(KEYINPUT83), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n443_), .A2(new_n394_), .ZN(new_n444_));
  NOR3_X1   g243(.A1(new_n444_), .A2(new_n386_), .A3(new_n393_), .ZN(new_n445_));
  AOI22_X1  g244(.A1(new_n432_), .A2(new_n435_), .B1(new_n442_), .B2(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n421_), .B1(new_n446_), .B2(new_n419_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT100), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n420_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n386_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n393_), .B1(new_n378_), .B2(new_n395_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n442_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n430_), .A2(new_n431_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n369_), .A2(KEYINPUT85), .ZN(new_n454_));
  INV_X1    g253(.A(new_n426_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n443_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n456_), .B1(new_n434_), .B2(KEYINPUT86), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n419_), .B(new_n452_), .C1(new_n453_), .C2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT20), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT100), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n368_), .B1(new_n449_), .B2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n421_), .B1(new_n403_), .B2(new_n419_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n452_), .B1(new_n457_), .B2(new_n453_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n410_), .A2(new_n416_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n418_), .A2(new_n417_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n463_), .A2(new_n466_), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n462_), .A2(new_n367_), .A3(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n364_), .B1(new_n461_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n368_), .ZN(new_n470_));
  OR2_X1    g269(.A1(new_n403_), .A2(new_n419_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n458_), .A2(new_n448_), .A3(KEYINPUT20), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n448_), .B1(new_n458_), .B2(KEYINPUT20), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n470_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n468_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n475_), .A2(new_n476_), .A3(new_n363_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n469_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT27), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n460_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n468_), .B1(new_n480_), .B2(new_n470_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n479_), .B1(new_n481_), .B2(new_n363_), .ZN(new_n482_));
  AND2_X1   g281(.A1(new_n462_), .A2(new_n467_), .ZN(new_n483_));
  OAI22_X1  g282(.A1(new_n480_), .A2(new_n470_), .B1(new_n367_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n364_), .ZN(new_n485_));
  AOI22_X1  g284(.A1(new_n478_), .A2(new_n479_), .B1(new_n482_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT87), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n446_), .A2(KEYINPUT30), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT30), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n463_), .A2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n487_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n491_));
  XOR2_X1   g290(.A(G127gat), .B(G134gat), .Z(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT89), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G127gat), .B(G134gat), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT89), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G113gat), .B(G120gat), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n493_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n497_), .B1(new_n493_), .B2(new_n496_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(KEYINPUT31), .ZN(new_n502_));
  INV_X1    g301(.A(new_n500_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(new_n498_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT31), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n502_), .A2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n491_), .A2(KEYINPUT88), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n446_), .A2(KEYINPUT30), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n463_), .A2(new_n489_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n509_), .A2(new_n510_), .A3(KEYINPUT87), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G71gat), .B(G99gat), .ZN(new_n512_));
  INV_X1    g311(.A(G43gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G227gat), .A2(G233gat), .ZN(new_n515_));
  INV_X1    g314(.A(G15gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n514_), .B(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n509_), .A2(new_n510_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n507_), .A2(KEYINPUT88), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n519_), .A2(new_n487_), .A3(new_n520_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n508_), .A2(new_n511_), .A3(new_n518_), .A4(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n511_), .A2(new_n518_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n521_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n520_), .B1(new_n519_), .B2(new_n487_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n523_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n522_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G225gat), .A2(G233gat), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G155gat), .A2(G162gat), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT91), .ZN(new_n531_));
  NOR3_X1   g330(.A1(new_n531_), .A2(G155gat), .A3(G162gat), .ZN(new_n532_));
  INV_X1    g331(.A(G155gat), .ZN(new_n533_));
  INV_X1    g332(.A(G162gat), .ZN(new_n534_));
  AOI21_X1  g333(.A(KEYINPUT91), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n530_), .B1(new_n532_), .B2(new_n535_), .ZN(new_n536_));
  AND3_X1   g335(.A1(KEYINPUT90), .A2(G141gat), .A3(G148gat), .ZN(new_n537_));
  AOI21_X1  g336(.A(KEYINPUT90), .B1(G141gat), .B2(G148gat), .ZN(new_n538_));
  NOR3_X1   g337(.A1(new_n537_), .A2(new_n538_), .A3(KEYINPUT2), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(G141gat), .A2(G148gat), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT3), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n544_));
  NAND3_X1  g343(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n543_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n536_), .B1(new_n540_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n530_), .A2(KEYINPUT1), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT1), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n550_), .A2(G155gat), .A3(G162gat), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n549_), .B(new_n551_), .C1(new_n532_), .C2(new_n535_), .ZN(new_n552_));
  NOR3_X1   g351(.A1(new_n537_), .A2(new_n538_), .A3(new_n541_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT92), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n552_), .A2(KEYINPUT92), .A3(new_n553_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n548_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n501_), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n552_), .A2(KEYINPUT92), .A3(new_n553_), .ZN(new_n560_));
  AOI21_X1  g359(.A(KEYINPUT92), .B1(new_n552_), .B2(new_n553_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n539_), .A2(new_n546_), .ZN(new_n562_));
  OAI22_X1  g361(.A1(new_n560_), .A2(new_n561_), .B1(new_n562_), .B2(new_n536_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(new_n504_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n529_), .B1(new_n559_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT102), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n566_), .B1(new_n564_), .B2(KEYINPUT4), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n559_), .A2(new_n564_), .A3(KEYINPUT4), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT4), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n563_), .A2(new_n504_), .A3(KEYINPUT102), .A4(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n567_), .A2(new_n568_), .A3(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n565_), .B1(new_n571_), .B2(new_n529_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G1gat), .B(G29gat), .ZN(new_n573_));
  INV_X1    g372(.A(G85gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT0), .B(G57gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n572_), .A2(new_n578_), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n572_), .A2(new_n578_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n527_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G228gat), .A2(G233gat), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT29), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n466_), .B(new_n582_), .C1(new_n558_), .C2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT96), .ZN(new_n585_));
  XOR2_X1   g384(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n586_));
  AOI21_X1  g385(.A(new_n419_), .B1(new_n563_), .B2(new_n586_), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n584_), .B(new_n585_), .C1(new_n587_), .C2(new_n582_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n586_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n466_), .B1(new_n558_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n582_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n585_), .B1(new_n593_), .B2(new_n584_), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n589_), .A2(new_n594_), .A3(G78gat), .ZN(new_n595_));
  INV_X1    g394(.A(G78gat), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n584_), .B1(new_n587_), .B2(new_n582_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(KEYINPUT96), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n596_), .B1(new_n598_), .B2(new_n588_), .ZN(new_n599_));
  OAI21_X1  g398(.A(G106gat), .B1(new_n595_), .B2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G22gat), .B(G50gat), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NOR3_X1   g401(.A1(new_n563_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT28), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n604_), .B1(new_n558_), .B2(new_n583_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n602_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n603_), .A2(new_n605_), .A3(new_n602_), .ZN(new_n608_));
  OAI21_X1  g407(.A(KEYINPUT97), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(G78gat), .B1(new_n589_), .B2(new_n594_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n598_), .A2(new_n596_), .A3(new_n588_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(new_n211_), .A3(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n600_), .A2(new_n610_), .A3(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  OR3_X1    g414(.A1(new_n607_), .A2(KEYINPUT97), .A3(new_n608_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n609_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n617_), .B1(new_n600_), .B2(new_n613_), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n486_), .B(new_n581_), .C1(new_n615_), .C2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT105), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n616_), .A2(new_n609_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n595_), .A2(new_n599_), .A3(G106gat), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n211_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n621_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(new_n614_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT105), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n625_), .A2(new_n626_), .A3(new_n486_), .A4(new_n581_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n620_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n527_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n580_), .A2(new_n579_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n624_), .A2(new_n631_), .A3(new_n614_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n482_), .A2(new_n485_), .ZN(new_n633_));
  AND3_X1   g432(.A1(new_n475_), .A2(new_n363_), .A3(new_n476_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n363_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n633_), .B1(new_n636_), .B2(KEYINPUT27), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n632_), .A2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n572_), .A2(new_n578_), .ZN(new_n639_));
  OAI21_X1  g438(.A(KEYINPUT103), .B1(new_n639_), .B2(KEYINPUT33), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n571_), .A2(new_n529_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n559_), .A2(new_n564_), .A3(new_n529_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(new_n578_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n639_), .B2(KEYINPUT33), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT103), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT33), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n646_), .B(new_n647_), .C1(new_n572_), .C2(new_n578_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n636_), .A2(new_n640_), .A3(new_n645_), .A4(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n363_), .A2(KEYINPUT32), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n484_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n475_), .A2(new_n476_), .A3(new_n650_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n653_), .A2(KEYINPUT104), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT104), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n655_), .B1(new_n481_), .B2(new_n650_), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n630_), .B(new_n652_), .C1(new_n654_), .C2(new_n656_), .ZN(new_n657_));
  AOI22_X1  g456(.A1(new_n649_), .A2(new_n657_), .B1(new_n614_), .B2(new_n624_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n629_), .B1(new_n638_), .B2(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n359_), .B1(new_n628_), .B2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n345_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n662_), .A2(new_n290_), .A3(new_n630_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT38), .ZN(new_n664_));
  INV_X1    g463(.A(new_n288_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n308_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n665_), .A2(new_n358_), .A3(new_n666_), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n667_), .A2(KEYINPUT106), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n331_), .A2(new_n332_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n333_), .A3(new_n337_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n671_), .B1(new_n628_), .B2(new_n659_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n667_), .A2(KEYINPUT106), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n668_), .A2(new_n672_), .A3(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G1gat), .B1(new_n674_), .B2(new_n631_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n664_), .A2(new_n675_), .ZN(G1324gat));
  NAND3_X1  g475(.A1(new_n662_), .A2(new_n291_), .A3(new_n637_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n668_), .A2(new_n672_), .A3(new_n673_), .A4(new_n637_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT39), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n678_), .A2(new_n679_), .A3(G8gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n678_), .B2(G8gat), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n677_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT40), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI211_X1 g483(.A(KEYINPUT40), .B(new_n677_), .C1(new_n680_), .C2(new_n681_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1325gat));
  NAND4_X1  g485(.A1(new_n668_), .A2(new_n672_), .A3(new_n673_), .A4(new_n527_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(G15gat), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT107), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT107), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n687_), .A2(new_n690_), .A3(G15gat), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT41), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n662_), .A2(new_n516_), .A3(new_n527_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n689_), .A2(KEYINPUT41), .A3(new_n691_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n694_), .A2(new_n695_), .A3(new_n696_), .ZN(G1326gat));
  OR3_X1    g496(.A1(new_n661_), .A2(G22gat), .A3(new_n625_), .ZN(new_n698_));
  OAI21_X1  g497(.A(G22gat), .B1(new_n674_), .B2(new_n625_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(KEYINPUT108), .B(KEYINPUT42), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n699_), .A2(new_n700_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n698_), .B1(new_n701_), .B2(new_n702_), .ZN(G1327gat));
  NOR2_X1   g502(.A1(new_n670_), .A2(new_n666_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n660_), .A2(new_n665_), .A3(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT110), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n706_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(G29gat), .B1(new_n709_), .B2(new_n630_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n628_), .A2(new_n659_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT109), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n339_), .A2(new_n714_), .A3(new_n343_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n339_), .B2(new_n343_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n712_), .B1(new_n713_), .B2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n344_), .A2(new_n712_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n719_), .B1(new_n628_), .B2(new_n659_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n288_), .A2(new_n359_), .A3(new_n666_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n711_), .B1(new_n721_), .B2(new_n723_), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n722_), .B(KEYINPUT44), .C1(new_n718_), .C2(new_n720_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n630_), .A2(G29gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n710_), .B1(new_n726_), .B2(new_n727_), .ZN(G1328gat));
  NOR2_X1   g527(.A1(new_n486_), .A2(G36gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n707_), .A2(new_n708_), .A3(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT45), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT45), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n707_), .A2(new_n732_), .A3(new_n708_), .A4(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n724_), .A2(new_n637_), .A3(new_n725_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(G36gat), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT46), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n734_), .A2(KEYINPUT46), .A3(new_n736_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1329gat));
  NAND4_X1  g540(.A1(new_n724_), .A2(G43gat), .A3(new_n527_), .A4(new_n725_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n707_), .A2(new_n527_), .A3(new_n708_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT111), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n743_), .A2(new_n744_), .A3(new_n513_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n743_), .B2(new_n513_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n742_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT47), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT47), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n749_), .B(new_n742_), .C1(new_n745_), .C2(new_n746_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(G1330gat));
  INV_X1    g550(.A(new_n625_), .ZN(new_n752_));
  AOI21_X1  g551(.A(G50gat), .B1(new_n709_), .B2(new_n752_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n752_), .A2(G50gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n726_), .B2(new_n754_), .ZN(G1331gat));
  NAND4_X1  g554(.A1(new_n672_), .A2(new_n359_), .A3(new_n288_), .A4(new_n666_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n757_), .A2(G57gat), .A3(new_n630_), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n713_), .A2(new_n359_), .A3(new_n288_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n344_), .A2(new_n308_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n759_), .A2(new_n630_), .A3(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(G57gat), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n761_), .A2(KEYINPUT112), .A3(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT112), .B1(new_n761_), .B2(new_n762_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n758_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT113), .Z(G1332gat));
  INV_X1    g565(.A(KEYINPUT48), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n757_), .A2(new_n637_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(G64gat), .ZN(new_n769_));
  INV_X1    g568(.A(G64gat), .ZN(new_n770_));
  AOI211_X1 g569(.A(KEYINPUT48), .B(new_n770_), .C1(new_n757_), .C2(new_n637_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n759_), .A2(new_n760_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n637_), .A2(new_n770_), .ZN(new_n773_));
  OAI22_X1  g572(.A1(new_n769_), .A2(new_n771_), .B1(new_n772_), .B2(new_n773_), .ZN(G1333gat));
  OR3_X1    g573(.A1(new_n772_), .A2(G71gat), .A3(new_n629_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n757_), .A2(new_n527_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT49), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n776_), .A2(new_n777_), .A3(G71gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n776_), .B2(G71gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(G1334gat));
  INV_X1    g579(.A(KEYINPUT50), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n757_), .A2(new_n752_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n782_), .B2(G78gat), .ZN(new_n783_));
  AOI211_X1 g582(.A(KEYINPUT50), .B(new_n596_), .C1(new_n757_), .C2(new_n752_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n752_), .A2(new_n596_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT114), .ZN(new_n786_));
  OAI22_X1  g585(.A1(new_n783_), .A2(new_n784_), .B1(new_n772_), .B2(new_n786_), .ZN(G1335gat));
  NAND2_X1  g586(.A1(new_n759_), .A2(new_n704_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n789_), .A2(new_n574_), .A3(new_n630_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n288_), .A2(new_n359_), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n721_), .A2(new_n791_), .A3(new_n666_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n792_), .A2(new_n630_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n790_), .B1(new_n793_), .B2(new_n574_), .ZN(G1336gat));
  AOI21_X1  g593(.A(G92gat), .B1(new_n789_), .B2(new_n637_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n637_), .A2(G92gat), .ZN(new_n796_));
  XOR2_X1   g595(.A(new_n796_), .B(KEYINPUT115), .Z(new_n797_));
  AOI21_X1  g596(.A(new_n795_), .B1(new_n792_), .B2(new_n797_), .ZN(G1337gat));
  NAND2_X1  g597(.A1(new_n792_), .A2(new_n527_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n527_), .A2(new_n210_), .ZN(new_n800_));
  AOI22_X1  g599(.A1(new_n799_), .A2(G99gat), .B1(new_n789_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT51), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n801_), .B(new_n803_), .ZN(G1338gat));
  NAND3_X1  g603(.A1(new_n789_), .A2(new_n211_), .A3(new_n752_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n791_), .A2(new_n666_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n752_), .B(new_n806_), .C1(new_n718_), .C2(new_n720_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(G106gat), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(new_n809_), .A3(KEYINPUT52), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n807_), .A2(new_n811_), .A3(G106gat), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT117), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n810_), .A2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n811_), .B1(new_n807_), .B2(G106gat), .ZN(new_n816_));
  OAI22_X1  g615(.A1(new_n816_), .A2(new_n809_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n805_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n805_), .B(new_n819_), .C1(new_n815_), .C2(new_n817_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(G1339gat));
  NAND2_X1  g622(.A1(new_n278_), .A2(new_n358_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n825_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n256_), .A2(KEYINPUT12), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n245_), .A2(new_n263_), .A3(new_n255_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n267_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n829_), .A2(KEYINPUT55), .A3(new_n830_), .A4(new_n262_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n257_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(G230gat), .A3(G233gat), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n826_), .A2(new_n831_), .A3(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n274_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT56), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n834_), .A2(KEYINPUT56), .A3(new_n274_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n824_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n350_), .A2(new_n347_), .A3(new_n352_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n357_), .B1(new_n351_), .B2(new_n348_), .ZN(new_n841_));
  AOI22_X1  g640(.A1(new_n353_), .A2(new_n357_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n279_), .A2(new_n280_), .A3(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n670_), .B1(new_n839_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  OAI211_X1 g645(.A(KEYINPUT57), .B(new_n670_), .C1(new_n839_), .C2(new_n843_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n278_), .A2(new_n842_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n834_), .A2(KEYINPUT56), .A3(new_n274_), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT56), .B1(new_n834_), .B2(new_n274_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n848_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT58), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  OAI211_X1 g652(.A(KEYINPUT58), .B(new_n848_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n344_), .A3(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n846_), .A2(new_n847_), .A3(new_n855_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n760_), .A2(new_n286_), .A3(new_n359_), .A4(new_n287_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(KEYINPUT54), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n665_), .A2(new_n859_), .A3(new_n359_), .A4(new_n760_), .ZN(new_n860_));
  AOI22_X1  g659(.A1(new_n856_), .A2(new_n308_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n625_), .A2(new_n630_), .A3(new_n486_), .A4(new_n527_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(G113gat), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n863_), .A2(new_n864_), .A3(new_n358_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n866_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n862_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n343_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n869_), .B1(new_n670_), .B2(new_n309_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n870_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n871_));
  AOI22_X1  g670(.A1(new_n845_), .A2(new_n844_), .B1(new_n871_), .B2(new_n854_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n666_), .B1(new_n872_), .B2(new_n847_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n858_), .A2(new_n860_), .ZN(new_n874_));
  OAI211_X1 g673(.A(KEYINPUT59), .B(new_n868_), .C1(new_n873_), .C2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n359_), .B1(new_n867_), .B2(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n865_), .B1(new_n876_), .B2(new_n864_), .ZN(G1340gat));
  INV_X1    g676(.A(G120gat), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n867_), .A2(new_n875_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n878_), .B1(new_n879_), .B2(new_n288_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n863_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n878_), .B1(new_n665_), .B2(KEYINPUT60), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n882_), .B1(KEYINPUT60), .B2(new_n878_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n881_), .A2(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(KEYINPUT120), .B1(new_n880_), .B2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n665_), .B1(new_n867_), .B2(new_n875_), .ZN(new_n887_));
  OAI221_X1 g686(.A(new_n886_), .B1(new_n881_), .B2(new_n883_), .C1(new_n887_), .C2(new_n878_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n885_), .A2(new_n888_), .ZN(G1341gat));
  AOI21_X1  g688(.A(G127gat), .B1(new_n863_), .B2(new_n666_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n666_), .A2(G127gat), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(KEYINPUT121), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n890_), .B1(new_n879_), .B2(new_n892_), .ZN(G1342gat));
  XOR2_X1   g692(.A(KEYINPUT122), .B(G134gat), .Z(new_n894_));
  NAND2_X1  g693(.A1(new_n344_), .A2(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n895_), .B1(new_n867_), .B2(new_n875_), .ZN(new_n896_));
  AOI21_X1  g695(.A(G134gat), .B1(new_n863_), .B2(new_n671_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT123), .ZN(new_n898_));
  OR3_X1    g697(.A1(new_n896_), .A2(new_n897_), .A3(new_n898_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(G1343gat));
  NAND3_X1  g700(.A1(new_n752_), .A2(new_n630_), .A3(new_n629_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n861_), .A2(new_n637_), .A3(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n358_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n288_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g706(.A1(new_n903_), .A2(new_n666_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT61), .B(G155gat), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n908_), .B(new_n909_), .ZN(G1346gat));
  AOI21_X1  g709(.A(G162gat), .B1(new_n903_), .B2(new_n671_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n715_), .A2(new_n716_), .A3(new_n534_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n911_), .B1(new_n903_), .B2(new_n912_), .ZN(G1347gat));
  AND2_X1   g712(.A1(new_n371_), .A2(new_n374_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n861_), .A2(new_n486_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT124), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n625_), .A2(new_n581_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n915_), .A2(new_n916_), .A3(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n916_), .B1(new_n915_), .B2(new_n917_), .ZN(new_n920_));
  OAI211_X1 g719(.A(new_n358_), .B(new_n914_), .C1(new_n919_), .C2(new_n920_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n915_), .A2(new_n358_), .A3(new_n917_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n923_));
  AND3_X1   g722(.A1(new_n922_), .A2(new_n923_), .A3(G169gat), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n923_), .B1(new_n922_), .B2(G169gat), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n921_), .B1(new_n924_), .B2(new_n925_), .ZN(G1348gat));
  NAND2_X1  g725(.A1(new_n915_), .A2(new_n917_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(KEYINPUT124), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(new_n918_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n929_), .A2(new_n372_), .A3(new_n288_), .ZN(new_n930_));
  OAI21_X1  g729(.A(G176gat), .B1(new_n927_), .B2(new_n665_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1349gat));
  AND2_X1   g731(.A1(new_n666_), .A2(new_n397_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n915_), .A2(new_n666_), .A3(new_n917_), .ZN(new_n934_));
  AOI22_X1  g733(.A1(new_n929_), .A2(new_n933_), .B1(new_n437_), .B2(new_n934_), .ZN(G1350gat));
  NOR2_X1   g734(.A1(new_n670_), .A2(new_n401_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n936_), .B1(new_n919_), .B2(new_n920_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n870_), .B1(new_n928_), .B2(new_n918_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n938_), .B2(new_n398_), .ZN(G1351gat));
  NOR2_X1   g738(.A1(new_n632_), .A2(new_n527_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n915_), .A2(new_n940_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n941_), .ZN(new_n942_));
  AOI21_X1  g741(.A(G197gat), .B1(new_n942_), .B2(new_n358_), .ZN(new_n943_));
  NAND4_X1  g742(.A1(new_n915_), .A2(G197gat), .A3(new_n358_), .A4(new_n940_), .ZN(new_n944_));
  AND2_X1   g743(.A1(new_n944_), .A2(KEYINPUT125), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n944_), .A2(KEYINPUT125), .ZN(new_n946_));
  NOR3_X1   g745(.A1(new_n943_), .A2(new_n945_), .A3(new_n946_), .ZN(G1352gat));
  NOR2_X1   g746(.A1(new_n941_), .A2(new_n665_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(new_n405_), .ZN(G1353gat));
  XOR2_X1   g748(.A(KEYINPUT63), .B(G211gat), .Z(new_n950_));
  NAND3_X1  g749(.A1(new_n942_), .A2(new_n666_), .A3(new_n950_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n952_), .B1(new_n941_), .B2(new_n308_), .ZN(new_n953_));
  AND2_X1   g752(.A1(new_n951_), .A2(new_n953_), .ZN(G1354gat));
  AOI21_X1  g753(.A(G218gat), .B1(new_n942_), .B2(new_n671_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n344_), .A2(G218gat), .ZN(new_n956_));
  XOR2_X1   g755(.A(new_n956_), .B(KEYINPUT126), .Z(new_n957_));
  AOI21_X1  g756(.A(new_n955_), .B1(new_n942_), .B2(new_n957_), .ZN(G1355gat));
endmodule


