//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 1 1 1 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n859_, new_n861_, new_n862_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n902_, new_n904_, new_n905_, new_n907_,
    new_n908_, new_n909_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT36), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT7), .ZN(new_n206_));
  INV_X1    g005(.A(G99gat), .ZN(new_n207_));
  INV_X1    g006(.A(G106gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT6), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n209_), .A2(new_n212_), .A3(new_n213_), .A4(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(G85gat), .B(G92gat), .Z(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT8), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  XOR2_X1   g019(.A(KEYINPUT10), .B(G99gat), .Z(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(new_n208_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n216_), .A2(KEYINPUT9), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n212_), .A2(new_n213_), .ZN(new_n224_));
  INV_X1    g023(.A(G85gat), .ZN(new_n225_));
  INV_X1    g024(.A(G92gat), .ZN(new_n226_));
  OR3_X1    g025(.A1(new_n225_), .A2(new_n226_), .A3(KEYINPUT9), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .A4(new_n227_), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n220_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n217_), .A2(new_n218_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n215_), .A2(KEYINPUT65), .A3(new_n216_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n230_), .A2(KEYINPUT8), .A3(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n229_), .A2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G29gat), .B(G36gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(G50gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT69), .B(G43gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(G50gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n234_), .B(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n236_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n237_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT70), .B1(new_n233_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT70), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n229_), .A2(new_n242_), .A3(new_n245_), .A4(new_n232_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT71), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n237_), .A2(new_n241_), .A3(KEYINPUT15), .ZN(new_n249_));
  AOI21_X1  g048(.A(KEYINPUT15), .B1(new_n237_), .B2(new_n241_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n248_), .B1(new_n251_), .B2(new_n233_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n247_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G232gat), .A2(G233gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT34), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n253_), .A2(KEYINPUT35), .A3(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT73), .ZN(new_n257_));
  INV_X1    g056(.A(new_n255_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT35), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n259_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n247_), .A2(new_n252_), .A3(new_n261_), .A4(new_n262_), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n256_), .A2(new_n257_), .A3(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n257_), .B1(new_n256_), .B2(new_n263_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n205_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT74), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT37), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT36), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n256_), .A2(new_n270_), .A3(new_n204_), .A4(new_n263_), .ZN(new_n271_));
  OAI211_X1 g070(.A(KEYINPUT74), .B(new_n205_), .C1(new_n264_), .C2(new_n265_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n268_), .A2(new_n269_), .A3(new_n271_), .A4(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT72), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n271_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n256_), .A2(new_n263_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(new_n205_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n271_), .A2(new_n274_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n275_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT37), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n273_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G15gat), .B(G22gat), .ZN(new_n282_));
  INV_X1    g081(.A(G1gat), .ZN(new_n283_));
  INV_X1    g082(.A(G8gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT14), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n282_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G1gat), .B(G8gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G231gat), .A2(G233gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G57gat), .B(G64gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT11), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G71gat), .B(G78gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n292_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n291_), .A2(KEYINPUT11), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n294_), .B1(new_n297_), .B2(new_n293_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n290_), .B(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n299_), .A2(KEYINPUT17), .ZN(new_n300_));
  XOR2_X1   g099(.A(KEYINPUT75), .B(KEYINPUT16), .Z(new_n301_));
  XNOR2_X1  g100(.A(G127gat), .B(G155gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G183gat), .B(G211gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  MUX2_X1   g104(.A(KEYINPUT17), .B(new_n300_), .S(new_n305_), .Z(new_n306_));
  INV_X1    g105(.A(KEYINPUT76), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n299_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n306_), .B(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n281_), .A2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT77), .ZN(new_n311_));
  XOR2_X1   g110(.A(G64gat), .B(G92gat), .Z(new_n312_));
  XNOR2_X1  g111(.A(G8gat), .B(G36gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT101), .B(KEYINPUT18), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(G183gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT79), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT79), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(G183gat), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n319_), .A2(new_n321_), .A3(KEYINPUT25), .ZN(new_n322_));
  OR2_X1    g121(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT26), .B(G190gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G183gat), .A2(G190gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT23), .ZN(new_n328_));
  NOR2_X1   g127(.A1(G169gat), .A2(G176gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT80), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT80), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n331_), .B1(G169gat), .B2(G176gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G169gat), .A2(G176gat), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n333_), .A2(KEYINPUT24), .A3(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT24), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n330_), .A2(new_n332_), .A3(new_n336_), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n326_), .A2(new_n328_), .A3(new_n335_), .A4(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(G204gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(G197gat), .ZN(new_n340_));
  INV_X1    g139(.A(G197gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(G204gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT21), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n340_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G211gat), .B(G218gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G197gat), .B(G204gat), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n343_), .A2(KEYINPUT91), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n344_), .B(new_n345_), .C1(new_n346_), .C2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n345_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n340_), .A2(new_n342_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(new_n351_), .A3(new_n347_), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n349_), .A2(new_n352_), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n319_), .A2(new_n321_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n328_), .B1(new_n354_), .B2(G190gat), .ZN(new_n355_));
  INV_X1    g154(.A(G176gat), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT81), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT22), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n356_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(G169gat), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n329_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n355_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n338_), .A2(new_n353_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT20), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT96), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT25), .B(G183gat), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n325_), .A2(KEYINPUT97), .ZN(new_n368_));
  INV_X1    g167(.A(G190gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT26), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT26), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(G190gat), .ZN(new_n372_));
  AND3_X1   g171(.A1(new_n370_), .A2(new_n372_), .A3(KEYINPUT97), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n367_), .B1(new_n368_), .B2(new_n373_), .ZN(new_n374_));
  XOR2_X1   g173(.A(KEYINPUT98), .B(KEYINPUT24), .Z(new_n375_));
  NAND3_X1  g174(.A1(new_n333_), .A2(new_n375_), .A3(new_n334_), .ZN(new_n376_));
  OR2_X1    g175(.A1(new_n333_), .A2(new_n375_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n374_), .A2(new_n376_), .A3(new_n377_), .A4(new_n328_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n328_), .B1(G183gat), .B2(G190gat), .ZN(new_n379_));
  XOR2_X1   g178(.A(new_n334_), .B(KEYINPUT99), .Z(new_n380_));
  XOR2_X1   g179(.A(KEYINPUT22), .B(G169gat), .Z(new_n381_));
  OAI211_X1 g180(.A(new_n379_), .B(new_n380_), .C1(G176gat), .C2(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n353_), .B1(new_n378_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n363_), .A2(KEYINPUT96), .A3(KEYINPUT20), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n366_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G226gat), .A2(G233gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT19), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n388_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n353_), .B1(new_n338_), .B2(new_n362_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT100), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT20), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n378_), .A2(new_n382_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n393_), .B1(new_n394_), .B2(new_n353_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n390_), .B1(new_n392_), .B2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n317_), .B1(new_n389_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n386_), .A2(new_n388_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n338_), .A2(new_n362_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n349_), .A2(new_n352_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT100), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT100), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n399_), .A2(new_n403_), .A3(new_n400_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n395_), .A2(new_n390_), .A3(new_n402_), .A4(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n398_), .A2(new_n316_), .A3(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n397_), .A2(KEYINPUT27), .A3(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT104), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n363_), .A2(KEYINPUT96), .A3(KEYINPUT20), .ZN(new_n409_));
  AOI21_X1  g208(.A(KEYINPUT96), .B1(new_n363_), .B2(KEYINPUT20), .ZN(new_n410_));
  NOR3_X1   g209(.A1(new_n409_), .A2(new_n410_), .A3(new_n383_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n405_), .B1(new_n411_), .B2(new_n390_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(new_n317_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n406_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT27), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT104), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n397_), .A2(new_n417_), .A3(KEYINPUT27), .A4(new_n406_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n408_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G1gat), .B(G29gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(G85gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT0), .B(G57gat), .ZN(new_n422_));
  XOR2_X1   g221(.A(new_n421_), .B(new_n422_), .Z(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G225gat), .A2(G233gat), .ZN(new_n425_));
  INV_X1    g224(.A(G155gat), .ZN(new_n426_));
  INV_X1    g225(.A(G162gat), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT1), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT1), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n429_), .A2(G155gat), .A3(G162gat), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n428_), .B(new_n430_), .C1(G155gat), .C2(G162gat), .ZN(new_n431_));
  INV_X1    g230(.A(G141gat), .ZN(new_n432_));
  INV_X1    g231(.A(G148gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G141gat), .A2(G148gat), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n431_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(G127gat), .ZN(new_n438_));
  INV_X1    g237(.A(G134gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(G113gat), .ZN(new_n441_));
  INV_X1    g240(.A(G120gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G127gat), .A2(G134gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G113gat), .A2(G120gat), .ZN(new_n445_));
  AND4_X1   g244(.A1(new_n440_), .A2(new_n443_), .A3(new_n444_), .A4(new_n445_), .ZN(new_n446_));
  AOI22_X1  g245(.A1(new_n440_), .A2(new_n444_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT102), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n440_), .A2(new_n444_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n443_), .A2(new_n445_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT102), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n440_), .A2(new_n443_), .A3(new_n444_), .A4(new_n445_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n451_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n448_), .A2(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n456_));
  XOR2_X1   g255(.A(new_n456_), .B(KEYINPUT87), .Z(new_n457_));
  INV_X1    g256(.A(KEYINPUT2), .ZN(new_n458_));
  OAI211_X1 g257(.A(G141gat), .B(G148gat), .C1(new_n458_), .C2(KEYINPUT88), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT88), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n435_), .A2(new_n460_), .A3(KEYINPUT2), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n459_), .A2(new_n461_), .B1(KEYINPUT88), .B2(new_n458_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT84), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT84), .B1(G141gat), .B2(G148gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  AND2_X1   g265(.A1(KEYINPUT85), .A2(KEYINPUT3), .ZN(new_n467_));
  NOR2_X1   g266(.A1(KEYINPUT85), .A2(KEYINPUT3), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n466_), .A2(KEYINPUT86), .A3(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(KEYINPUT86), .B1(new_n466_), .B2(new_n469_), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n457_), .B(new_n462_), .C1(new_n470_), .C2(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(G155gat), .B(G162gat), .Z(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT89), .ZN(new_n474_));
  AOI211_X1 g273(.A(new_n437_), .B(new_n455_), .C1(new_n472_), .C2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT83), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n451_), .A2(new_n476_), .A3(new_n453_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n446_), .A2(KEYINPUT83), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n472_), .A2(new_n474_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n480_), .B1(new_n481_), .B2(new_n436_), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT4), .B1(new_n475_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n436_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n479_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT4), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n425_), .B1(new_n483_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n455_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n481_), .A2(new_n436_), .A3(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n485_), .A2(new_n425_), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n424_), .B1(new_n488_), .B2(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(KEYINPUT4), .B1(new_n484_), .B2(new_n479_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n437_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n490_), .B1(new_n480_), .B2(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n494_), .B1(new_n496_), .B2(KEYINPUT4), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n491_), .B(new_n423_), .C1(new_n497_), .C2(new_n425_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n493_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G71gat), .B(G99gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G227gat), .A2(G233gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  XOR2_X1   g302(.A(G15gat), .B(G43gat), .Z(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n399_), .B(KEYINPUT30), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT82), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n505_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n506_), .B(new_n507_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n508_), .B1(new_n509_), .B2(new_n505_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n479_), .B(KEYINPUT31), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n512_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  XOR2_X1   g315(.A(G78gat), .B(G106gat), .Z(new_n517_));
  INV_X1    g316(.A(KEYINPUT29), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n400_), .B1(new_n495_), .B2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n400_), .A2(KEYINPUT92), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G228gat), .A2(G233gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT90), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n521_), .A2(KEYINPUT90), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n520_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n519_), .B(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT95), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n517_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT28), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n528_), .B1(new_n495_), .B2(new_n518_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n495_), .A2(new_n528_), .A3(new_n518_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G22gat), .B(G50gat), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n530_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n524_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n519_), .B(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT95), .ZN(new_n536_));
  INV_X1    g335(.A(new_n532_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n531_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n537_), .B1(new_n538_), .B2(new_n529_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n527_), .A2(new_n533_), .A3(new_n536_), .A4(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n533_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT94), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n517_), .B(KEYINPUT93), .Z(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n542_), .A2(new_n525_), .A3(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n535_), .A2(new_n543_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n525_), .A2(new_n544_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n546_), .A2(new_n547_), .A3(KEYINPUT94), .A4(new_n541_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n540_), .A2(new_n545_), .A3(new_n548_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n419_), .A2(new_n500_), .A3(new_n516_), .A4(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n408_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n500_), .A2(new_n548_), .A3(new_n540_), .A4(new_n545_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n488_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT33), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n556_), .A2(new_n557_), .A3(new_n491_), .A4(new_n423_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n498_), .A2(KEYINPUT33), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n425_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n485_), .A2(new_n561_), .A3(new_n490_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n424_), .B(new_n562_), .C1(new_n497_), .C2(new_n561_), .ZN(new_n563_));
  AND3_X1   g362(.A1(new_n413_), .A2(new_n563_), .A3(new_n406_), .ZN(new_n564_));
  AND3_X1   g363(.A1(new_n560_), .A2(new_n564_), .A3(KEYINPUT103), .ZN(new_n565_));
  AOI21_X1  g364(.A(KEYINPUT103), .B1(new_n560_), .B2(new_n564_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n316_), .A2(KEYINPUT32), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n398_), .A2(new_n567_), .A3(new_n405_), .ZN(new_n568_));
  OAI211_X1 g367(.A(KEYINPUT32), .B(new_n316_), .C1(new_n389_), .C2(new_n396_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n499_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n565_), .A2(new_n566_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n549_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n555_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n551_), .B1(new_n574_), .B2(new_n515_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n311_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT68), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n233_), .A2(new_n298_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n298_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n579_), .A2(new_n229_), .A3(new_n232_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n578_), .A2(KEYINPUT12), .A3(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT12), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n233_), .A2(new_n582_), .A3(new_n298_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G230gat), .A2(G233gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT64), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT66), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n586_), .B1(new_n578_), .B2(new_n580_), .ZN(new_n588_));
  AOI22_X1  g387(.A1(new_n584_), .A2(new_n586_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n588_), .A2(new_n587_), .ZN(new_n590_));
  XOR2_X1   g389(.A(G176gat), .B(G204gat), .Z(new_n591_));
  XNOR2_X1  g390(.A(G120gat), .B(G148gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n589_), .A2(new_n590_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n595_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n577_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n598_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n600_), .A2(KEYINPUT68), .A3(new_n596_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT13), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n599_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n602_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n288_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n249_), .A2(new_n250_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT78), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G229gat), .A2(G233gat), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n242_), .A2(new_n607_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n608_), .A2(new_n609_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n610_), .A2(new_n611_), .A3(new_n612_), .A4(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n242_), .B(new_n607_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n611_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n614_), .A2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G113gat), .B(G141gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G169gat), .B(G197gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n618_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n618_), .A2(new_n621_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n606_), .A2(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n576_), .A2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n627_), .A2(new_n283_), .A3(new_n499_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT38), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n268_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(new_n309_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n575_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(new_n626_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G1gat), .B1(new_n633_), .B2(new_n500_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT105), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n629_), .A2(new_n635_), .ZN(G1324gat));
  INV_X1    g435(.A(KEYINPUT107), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n632_), .A2(new_n626_), .A3(new_n552_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT106), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(new_n639_), .A3(G8gat), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n639_), .B1(new_n638_), .B2(G8gat), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n637_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n638_), .A2(G8gat), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT106), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n645_), .A2(KEYINPUT107), .A3(new_n640_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n643_), .A2(new_n646_), .A3(KEYINPUT39), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n627_), .A2(new_n284_), .A3(new_n552_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT39), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n637_), .B(new_n649_), .C1(new_n641_), .C2(new_n642_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n647_), .A2(new_n648_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT40), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n647_), .A2(KEYINPUT40), .A3(new_n648_), .A4(new_n650_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1325gat));
  OAI21_X1  g454(.A(G15gat), .B1(new_n633_), .B2(new_n515_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT41), .Z(new_n657_));
  INV_X1    g456(.A(G15gat), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n627_), .A2(new_n658_), .A3(new_n516_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(G1326gat));
  OAI21_X1  g459(.A(G22gat), .B1(new_n633_), .B2(new_n549_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT42), .ZN(new_n662_));
  INV_X1    g461(.A(G22gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n627_), .A2(new_n663_), .A3(new_n573_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT108), .ZN(G1327gat));
  NAND2_X1  g465(.A1(new_n281_), .A2(KEYINPUT109), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT109), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n273_), .A2(new_n668_), .A3(new_n280_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(KEYINPUT43), .B1(new_n575_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT110), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n281_), .A2(KEYINPUT43), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n672_), .B1(new_n575_), .B2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n483_), .A2(new_n487_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n492_), .B1(new_n677_), .B2(new_n561_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n557_), .B1(new_n678_), .B2(new_n423_), .ZN(new_n679_));
  NOR4_X1   g478(.A1(new_n488_), .A2(new_n492_), .A3(KEYINPUT33), .A4(new_n424_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n413_), .A2(new_n563_), .A3(new_n406_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n676_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n560_), .A2(new_n564_), .A3(KEYINPUT103), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n683_), .A2(new_n570_), .A3(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n554_), .B1(new_n685_), .B2(new_n549_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n550_), .B1(new_n686_), .B2(new_n516_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n687_), .A2(KEYINPUT110), .A3(new_n673_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n671_), .A2(new_n675_), .A3(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n309_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n626_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n689_), .A2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(KEYINPUT111), .B(KEYINPUT44), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n689_), .A2(KEYINPUT44), .A3(new_n692_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n695_), .A2(new_n499_), .A3(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(G29gat), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n691_), .A2(new_n575_), .A3(new_n630_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n700_), .A2(G29gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n698_), .B1(new_n500_), .B2(new_n701_), .ZN(G1328gat));
  AND3_X1   g501(.A1(new_n687_), .A2(KEYINPUT110), .A3(new_n673_), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT110), .B1(new_n687_), .B2(new_n673_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n691_), .B1(new_n705_), .B2(new_n671_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n694_), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n552_), .B(new_n696_), .C1(new_n706_), .C2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(G36gat), .ZN(new_n709_));
  INV_X1    g508(.A(G36gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n699_), .A2(new_n710_), .A3(new_n552_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT45), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n699_), .A2(KEYINPUT45), .A3(new_n710_), .A4(new_n552_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n709_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT112), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT46), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n715_), .B1(new_n708_), .B2(G36gat), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT46), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n720_), .A2(KEYINPUT112), .A3(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n719_), .A2(new_n722_), .ZN(G1329gat));
  NAND4_X1  g522(.A1(new_n695_), .A2(G43gat), .A3(new_n516_), .A4(new_n696_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n700_), .A2(new_n515_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(G43gat), .B2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n726_), .B(new_n727_), .ZN(G1330gat));
  NAND3_X1  g527(.A1(new_n699_), .A2(new_n238_), .A3(new_n573_), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n695_), .A2(new_n573_), .A3(new_n696_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(new_n730_), .B2(new_n238_), .ZN(G1331gat));
  NOR2_X1   g530(.A1(new_n605_), .A2(new_n624_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n632_), .A2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(G57gat), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n734_), .A2(new_n735_), .A3(new_n500_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n576_), .A2(new_n732_), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n737_), .A2(KEYINPUT114), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(KEYINPUT114), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n738_), .A2(new_n499_), .A3(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n736_), .B1(new_n740_), .B2(new_n735_), .ZN(G1332gat));
  OAI21_X1  g540(.A(G64gat), .B1(new_n734_), .B2(new_n419_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT48), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n419_), .A2(G64gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(new_n737_), .B2(new_n744_), .ZN(G1333gat));
  INV_X1    g544(.A(G71gat), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n746_), .B1(new_n733_), .B2(new_n516_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(KEYINPUT115), .B(KEYINPUT49), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n747_), .A2(new_n748_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n516_), .A2(new_n746_), .ZN(new_n751_));
  OAI22_X1  g550(.A1(new_n749_), .A2(new_n750_), .B1(new_n737_), .B2(new_n751_), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n752_), .B(KEYINPUT116), .Z(G1334gat));
  OAI21_X1  g552(.A(G78gat), .B1(new_n734_), .B2(new_n549_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT50), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n549_), .A2(G78gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n755_), .B1(new_n737_), .B2(new_n756_), .ZN(G1335gat));
  NAND2_X1  g556(.A1(new_n732_), .A2(new_n690_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n705_), .B2(new_n671_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n759_), .A2(G85gat), .A3(new_n499_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n575_), .A2(new_n630_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n758_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n225_), .B1(new_n763_), .B2(new_n500_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n760_), .A2(new_n764_), .ZN(G1336gat));
  INV_X1    g564(.A(new_n763_), .ZN(new_n766_));
  AOI21_X1  g565(.A(G92gat), .B1(new_n766_), .B2(new_n552_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n419_), .A2(new_n226_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n759_), .B2(new_n768_), .ZN(G1337gat));
  AOI21_X1  g568(.A(new_n207_), .B1(new_n759_), .B2(new_n516_), .ZN(new_n770_));
  AND2_X1   g569(.A1(KEYINPUT117), .A2(KEYINPUT51), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n766_), .A2(new_n221_), .A3(new_n516_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n770_), .A2(new_n771_), .A3(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(KEYINPUT117), .A2(KEYINPUT51), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n773_), .B(new_n774_), .ZN(G1338gat));
  NAND3_X1  g574(.A1(new_n766_), .A2(new_n208_), .A3(new_n573_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n689_), .A2(new_n573_), .A3(new_n762_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n777_), .A2(new_n778_), .A3(G106gat), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n777_), .B2(G106gat), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n776_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g581(.A1(new_n281_), .A2(new_n605_), .A3(new_n625_), .A4(new_n309_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT54), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n783_), .B(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT120), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n584_), .A2(new_n586_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n586_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n581_), .A2(new_n788_), .A3(new_n583_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n787_), .A2(KEYINPUT55), .A3(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n595_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT55), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n584_), .A2(new_n792_), .A3(new_n586_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n790_), .A2(new_n791_), .A3(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT56), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT118), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n790_), .A2(KEYINPUT56), .A3(new_n791_), .A4(new_n793_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n796_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n794_), .A2(KEYINPUT118), .A3(new_n795_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n799_), .A2(new_n624_), .A3(new_n596_), .A4(new_n800_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n610_), .A2(new_n616_), .A3(new_n612_), .A4(new_n613_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n615_), .A2(new_n611_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n621_), .A3(new_n803_), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n622_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(new_n601_), .A3(new_n599_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n801_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n630_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT57), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n786_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n807_), .A2(KEYINPUT120), .A3(KEYINPUT57), .A4(new_n630_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n796_), .A2(new_n798_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n805_), .A2(new_n813_), .A3(new_n596_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT58), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n805_), .A2(new_n813_), .A3(KEYINPUT58), .A4(new_n596_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n281_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(KEYINPUT119), .A3(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n816_), .A2(new_n280_), .A3(new_n273_), .A4(new_n817_), .ZN(new_n822_));
  AOI22_X1  g621(.A1(new_n821_), .A2(new_n822_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n812_), .A2(new_n820_), .A3(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n785_), .B1(new_n824_), .B2(new_n690_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n419_), .A2(new_n549_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n826_), .A2(new_n500_), .A3(new_n515_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT59), .B1(new_n825_), .B2(new_n828_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n828_), .A2(KEYINPUT59), .ZN(new_n830_));
  AOI22_X1  g629(.A1(new_n810_), .A2(new_n811_), .B1(new_n819_), .B2(new_n818_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n808_), .A2(new_n809_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n309_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n830_), .B1(new_n833_), .B2(new_n785_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n829_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n836_));
  OAI21_X1  g635(.A(G113gat), .B1(new_n625_), .B2(new_n836_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n835_), .B(new_n837_), .C1(new_n836_), .C2(G113gat), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n825_), .A2(new_n828_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n441_), .B1(new_n840_), .B2(new_n625_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n838_), .A2(new_n841_), .ZN(G1340gat));
  OAI21_X1  g641(.A(new_n442_), .B1(new_n605_), .B2(KEYINPUT60), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n839_), .B(new_n843_), .C1(KEYINPUT60), .C2(new_n442_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n835_), .A2(new_n606_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n845_), .B2(new_n442_), .ZN(G1341gat));
  OAI21_X1  g645(.A(new_n438_), .B1(new_n840_), .B2(new_n690_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n829_), .A2(new_n834_), .A3(G127gat), .A4(new_n309_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT122), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT122), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n847_), .A2(new_n848_), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(G1342gat));
  NAND3_X1  g652(.A1(new_n835_), .A2(G134gat), .A3(new_n819_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n439_), .B1(new_n840_), .B2(new_n630_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n854_), .A2(new_n855_), .ZN(G1343gat));
  NOR3_X1   g655(.A1(new_n825_), .A2(new_n549_), .A3(new_n516_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n552_), .A2(new_n500_), .ZN(new_n858_));
  AND3_X1   g657(.A1(new_n857_), .A2(new_n624_), .A3(new_n858_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(new_n432_), .ZN(G1344gat));
  AND2_X1   g659(.A1(new_n857_), .A2(new_n858_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n606_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(G148gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n861_), .A2(new_n433_), .A3(new_n606_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(G1345gat));
  NAND2_X1  g664(.A1(new_n824_), .A2(new_n690_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n785_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n516_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n868_), .A2(new_n573_), .A3(new_n309_), .A4(new_n858_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(KEYINPUT123), .ZN(new_n870_));
  XOR2_X1   g669(.A(KEYINPUT61), .B(G155gat), .Z(new_n871_));
  INV_X1    g670(.A(KEYINPUT123), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n857_), .A2(new_n872_), .A3(new_n309_), .A4(new_n858_), .ZN(new_n873_));
  AND3_X1   g672(.A1(new_n870_), .A2(new_n871_), .A3(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n871_), .B1(new_n870_), .B2(new_n873_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n874_), .A2(new_n875_), .ZN(G1346gat));
  INV_X1    g675(.A(new_n630_), .ZN(new_n877_));
  AOI21_X1  g676(.A(G162gat), .B1(new_n861_), .B2(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n670_), .A2(new_n427_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(KEYINPUT124), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n878_), .B1(new_n861_), .B2(new_n880_), .ZN(G1347gat));
  NOR4_X1   g680(.A1(new_n419_), .A2(new_n515_), .A3(new_n573_), .A4(new_n499_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n624_), .B(new_n882_), .C1(new_n833_), .C2(new_n785_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(G169gat), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT62), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  OR2_X1    g685(.A1(new_n883_), .A2(new_n381_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n883_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n886_), .A2(new_n887_), .A3(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT125), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n886_), .A2(new_n887_), .A3(KEYINPUT125), .A4(new_n888_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1348gat));
  OR2_X1    g692(.A1(new_n833_), .A2(new_n785_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n882_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(G176gat), .B1(new_n896_), .B2(new_n606_), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n825_), .A2(new_n356_), .A3(new_n605_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n897_), .B1(new_n882_), .B2(new_n898_), .ZN(G1349gat));
  NOR3_X1   g698(.A1(new_n895_), .A2(new_n367_), .A3(new_n690_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n354_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n785_), .A2(new_n309_), .A3(new_n882_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n900_), .B1(new_n901_), .B2(new_n902_), .ZN(G1350gat));
  OAI21_X1  g702(.A(G190gat), .B1(new_n895_), .B2(new_n281_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n877_), .B1(new_n368_), .B2(new_n373_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n895_), .B2(new_n905_), .ZN(G1351gat));
  NOR2_X1   g705(.A1(new_n419_), .A2(new_n499_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n857_), .A2(new_n907_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n908_), .A2(new_n625_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(new_n341_), .ZN(G1352gat));
  NOR2_X1   g709(.A1(new_n908_), .A2(new_n605_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(new_n339_), .ZN(G1353gat));
  INV_X1    g711(.A(KEYINPUT63), .ZN(new_n913_));
  INV_X1    g712(.A(G211gat), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n309_), .B1(new_n913_), .B2(new_n914_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(KEYINPUT126), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n857_), .A2(new_n907_), .A3(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n913_), .A2(new_n914_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n917_), .B(new_n918_), .ZN(G1354gat));
  INV_X1    g718(.A(G218gat), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n908_), .A2(new_n920_), .A3(new_n281_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n857_), .A2(new_n877_), .A3(new_n907_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n921_), .B1(new_n920_), .B2(new_n922_), .ZN(G1355gat));
endmodule


