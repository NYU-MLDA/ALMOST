//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n812_, new_n813_, new_n814_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n932_,
    new_n933_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n954_,
    new_n955_, new_n957_, new_n958_, new_n959_, new_n961_, new_n963_,
    new_n964_, new_n965_, new_n967_, new_n968_, new_n969_, new_n970_;
  INV_X1    g000(.A(G169gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT22), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT22), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G169gat), .ZN(new_n205_));
  INV_X1    g004(.A(G176gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n203_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n207_), .B1(new_n202_), .B2(new_n206_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT78), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n202_), .A2(new_n206_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT22), .B(G169gat), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n211_), .B1(new_n212_), .B2(new_n206_), .ZN(new_n213_));
  INV_X1    g012(.A(G183gat), .ZN(new_n214_));
  INV_X1    g013(.A(G190gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT23), .B1(new_n214_), .B2(new_n215_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(G183gat), .A3(G190gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  AOI22_X1  g019(.A1(new_n213_), .A2(KEYINPUT78), .B1(new_n216_), .B2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT24), .B1(new_n202_), .B2(new_n206_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n224_), .B1(new_n225_), .B2(new_n222_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT25), .B(G183gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT76), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT26), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n228_), .B1(new_n229_), .B2(G190gat), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n227_), .A2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n229_), .A2(G190gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n215_), .A2(KEYINPUT26), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT76), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n226_), .B1(new_n231_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT77), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n219_), .A2(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n219_), .A2(new_n236_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n217_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  AOI22_X1  g038(.A1(new_n210_), .A2(new_n221_), .B1(new_n235_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT88), .ZN(new_n241_));
  INV_X1    g040(.A(G211gat), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n242_), .A2(G218gat), .ZN(new_n243_));
  INV_X1    g042(.A(G218gat), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n244_), .A2(G211gat), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n241_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(G211gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n242_), .A2(G218gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n247_), .A2(new_n248_), .A3(KEYINPUT88), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(G204gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(G197gat), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n251_), .A2(G197gat), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT21), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(KEYINPUT87), .B1(new_n251_), .B2(G197gat), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT87), .ZN(new_n257_));
  INV_X1    g056(.A(G197gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n257_), .A2(new_n258_), .A3(G204gat), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n256_), .A2(new_n259_), .A3(new_n252_), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n250_), .B(new_n255_), .C1(KEYINPUT21), .C2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT89), .ZN(new_n262_));
  AND3_X1   g061(.A1(new_n247_), .A2(new_n248_), .A3(KEYINPUT88), .ZN(new_n263_));
  AOI21_X1  g062(.A(KEYINPUT88), .B1(new_n247_), .B2(new_n248_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n262_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n246_), .A2(KEYINPUT89), .A3(new_n249_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n260_), .A2(KEYINPUT21), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT90), .B1(new_n267_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT90), .ZN(new_n271_));
  AOI211_X1 g070(.A(new_n271_), .B(new_n268_), .C1(new_n265_), .C2(new_n266_), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n240_), .B(new_n261_), .C1(new_n270_), .C2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n261_), .ZN(new_n274_));
  NOR3_X1   g073(.A1(new_n263_), .A2(new_n264_), .A3(new_n262_), .ZN(new_n275_));
  AOI21_X1  g074(.A(KEYINPUT89), .B1(new_n246_), .B2(new_n249_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n269_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n271_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n267_), .A2(KEYINPUT90), .A3(new_n269_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n274_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n239_), .A2(new_n216_), .ZN(new_n281_));
  NOR3_X1   g080(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n223_), .B1(G169gat), .B2(G176gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n222_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n282_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n285_), .A2(new_n220_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT26), .B(G190gat), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT92), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT92), .B1(new_n232_), .B2(new_n233_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n289_), .A2(new_n290_), .A3(new_n227_), .ZN(new_n291_));
  AOI22_X1  g090(.A1(new_n281_), .A2(new_n213_), .B1(new_n286_), .B2(new_n291_), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n273_), .B(KEYINPUT20), .C1(new_n280_), .C2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G226gat), .A2(G233gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT19), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n295_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT20), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n261_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n207_), .B(KEYINPUT78), .C1(new_n202_), .C2(new_n206_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n220_), .A2(new_n216_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n213_), .A2(KEYINPUT78), .ZN(new_n303_));
  OAI211_X1 g102(.A(new_n227_), .B(new_n230_), .C1(new_n287_), .C2(new_n228_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n285_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n217_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n219_), .A2(new_n236_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n219_), .A2(new_n236_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n306_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  OAI22_X1  g108(.A1(new_n302_), .A2(new_n303_), .B1(new_n305_), .B2(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n298_), .B1(new_n299_), .B2(new_n310_), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n261_), .B(new_n292_), .C1(new_n270_), .C2(new_n272_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n296_), .A2(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(G8gat), .B(G36gat), .Z(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G64gat), .B(G92gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n314_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n319_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n296_), .A2(new_n321_), .A3(new_n313_), .ZN(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT27), .B1(new_n320_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT99), .ZN(new_n324_));
  XOR2_X1   g123(.A(KEYINPUT96), .B(KEYINPUT20), .Z(new_n325_));
  NAND3_X1  g124(.A1(new_n312_), .A2(KEYINPUT97), .A3(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n299_), .A2(new_n310_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(KEYINPUT97), .B1(new_n312_), .B2(new_n325_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n295_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n293_), .A2(new_n295_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n321_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n322_), .A2(KEYINPUT27), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n324_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT27), .ZN(new_n335_));
  AOI22_X1  g134(.A1(new_n293_), .A2(new_n295_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n335_), .B1(new_n336_), .B2(new_n321_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n293_), .A2(new_n295_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n312_), .A2(new_n325_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT97), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n341_), .A2(new_n327_), .A3(new_n326_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n338_), .B1(new_n342_), .B2(new_n295_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n337_), .B(KEYINPUT99), .C1(new_n343_), .C2(new_n321_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n323_), .B1(new_n334_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G141gat), .A2(G148gat), .ZN(new_n346_));
  NOR2_X1   g145(.A1(G141gat), .A2(G148gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT82), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n346_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n349_), .B1(new_n348_), .B2(new_n347_), .ZN(new_n350_));
  INV_X1    g149(.A(G155gat), .ZN(new_n351_));
  INV_X1    g150(.A(G162gat), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(new_n352_), .A3(KEYINPUT83), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT83), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n354_), .B1(G155gat), .B2(G162gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G155gat), .A2(G162gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT1), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n350_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n346_), .A2(KEYINPUT2), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT2), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n361_), .A2(G141gat), .A3(G148gat), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT3), .ZN(new_n363_));
  AOI22_X1  g162(.A1(new_n360_), .A2(new_n362_), .B1(new_n363_), .B2(new_n347_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT84), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  OAI211_X1 g166(.A(KEYINPUT84), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT85), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n364_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n353_), .A2(new_n355_), .A3(KEYINPUT86), .A4(new_n357_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n353_), .A2(new_n355_), .A3(new_n357_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT86), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n371_), .A2(new_n372_), .A3(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n370_), .B1(new_n364_), .B2(new_n369_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n359_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G127gat), .B(G134gat), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G113gat), .B(G120gat), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n379_), .A2(new_n381_), .ZN(new_n384_));
  AOI21_X1  g183(.A(KEYINPUT79), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT79), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n386_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n378_), .A2(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n379_), .A2(new_n381_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n384_), .ZN(new_n391_));
  OAI221_X1 g190(.A(new_n359_), .B1(new_n390_), .B2(new_n391_), .C1(new_n376_), .C2(new_n377_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n389_), .A2(new_n392_), .A3(KEYINPUT4), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G225gat), .A2(G233gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT94), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT4), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n378_), .A2(new_n396_), .A3(new_n388_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n393_), .A2(new_n395_), .A3(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n395_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n389_), .A2(new_n392_), .A3(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G1gat), .B(G29gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(G85gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT0), .B(G57gat), .ZN(new_n403_));
  XOR2_X1   g202(.A(new_n402_), .B(new_n403_), .Z(new_n404_));
  AND3_X1   g203(.A1(new_n398_), .A2(new_n400_), .A3(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n404_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT98), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n398_), .A2(new_n400_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n404_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n398_), .A2(new_n400_), .A3(new_n404_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT98), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n410_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n407_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(G228gat), .ZN(new_n415_));
  INV_X1    g214(.A(G233gat), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n378_), .A2(KEYINPUT29), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n299_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n418_), .B1(new_n299_), .B2(new_n419_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G22gat), .B(G50gat), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n424_), .B(KEYINPUT28), .Z(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n426_), .B1(new_n378_), .B2(KEYINPUT29), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n364_), .A2(new_n369_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT85), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n429_), .A2(new_n371_), .A3(new_n372_), .A4(new_n375_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT29), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n430_), .A2(new_n431_), .A3(new_n359_), .A4(new_n425_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n427_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT91), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  XOR2_X1   g234(.A(G78gat), .B(G106gat), .Z(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n427_), .A2(KEYINPUT91), .A3(new_n432_), .A4(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n436_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n423_), .A2(new_n435_), .A3(new_n438_), .A4(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n438_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n422_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n442_), .A2(new_n435_), .A3(new_n420_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n440_), .A2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT31), .B1(new_n385_), .B2(new_n387_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n386_), .B1(new_n391_), .B2(new_n390_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n387_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT31), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n446_), .A2(new_n450_), .A3(KEYINPUT80), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G227gat), .A2(G233gat), .ZN(new_n452_));
  INV_X1    g251(.A(G15gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT30), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n310_), .A2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G71gat), .B(G99gat), .ZN(new_n458_));
  INV_X1    g257(.A(G43gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n221_), .A2(new_n210_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n239_), .A2(new_n285_), .A3(new_n304_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(new_n463_), .A3(new_n455_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n457_), .A2(new_n461_), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n461_), .B1(new_n457_), .B2(new_n464_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n451_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT81), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT80), .ZN(new_n470_));
  NOR3_X1   g269(.A1(new_n385_), .A2(KEYINPUT31), .A3(new_n387_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n449_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n470_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(new_n451_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n310_), .A2(new_n456_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n455_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n460_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n474_), .A2(new_n477_), .A3(new_n465_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n468_), .A2(new_n469_), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n469_), .B1(new_n468_), .B2(new_n478_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n445_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n468_), .A2(new_n478_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n440_), .A2(new_n444_), .A3(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n414_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT33), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n411_), .A2(new_n486_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n398_), .A2(KEYINPUT33), .A3(new_n400_), .A4(new_n404_), .ZN(new_n488_));
  AND2_X1   g287(.A1(new_n389_), .A2(new_n392_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n404_), .B1(new_n489_), .B2(new_n395_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT95), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n393_), .A2(new_n399_), .A3(new_n397_), .ZN(new_n492_));
  AND3_X1   g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n491_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n487_), .B(new_n488_), .C1(new_n493_), .C2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n320_), .A2(new_n322_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n321_), .A2(KEYINPUT32), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  OAI22_X1  g297(.A1(new_n405_), .A2(new_n406_), .B1(new_n314_), .B2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n497_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n500_));
  OAI22_X1  g299(.A1(new_n495_), .A2(new_n496_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n481_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n502_), .A2(new_n445_), .ZN(new_n503_));
  AOI22_X1  g302(.A1(new_n345_), .A2(new_n485_), .B1(new_n501_), .B2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G29gat), .B(G36gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G43gat), .B(G50gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT15), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G15gat), .B(G22gat), .ZN(new_n509_));
  INV_X1    g308(.A(G1gat), .ZN(new_n510_));
  INV_X1    g309(.A(G8gat), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT14), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n509_), .A2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G1gat), .B(G8gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n508_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n515_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(new_n507_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G229gat), .A2(G233gat), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n516_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n507_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n515_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n518_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n519_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n520_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G113gat), .B(G141gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G169gat), .B(G197gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n527_), .B(new_n528_), .Z(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n526_), .A2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n520_), .A2(new_n525_), .A3(new_n529_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(KEYINPUT75), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT75), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n526_), .A2(new_n534_), .A3(new_n530_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n504_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT8), .ZN(new_n538_));
  OR3_X1    g337(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT6), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT66), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT66), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT6), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G99gat), .A2(G106gat), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n543_), .A2(new_n545_), .A3(G99gat), .A4(G106gat), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n541_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(G85gat), .B(G92gat), .Z(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n538_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n539_), .A2(new_n540_), .ZN(new_n554_));
  AND4_X1   g353(.A1(G99gat), .A2(new_n543_), .A3(new_n545_), .A4(G106gat), .ZN(new_n555_));
  AOI22_X1  g354(.A1(new_n543_), .A2(new_n545_), .B1(G99gat), .B2(G106gat), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n554_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n557_), .A2(KEYINPUT8), .A3(new_n551_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n548_), .A2(new_n549_), .ZN(new_n559_));
  INV_X1    g358(.A(G85gat), .ZN(new_n560_));
  INV_X1    g359(.A(G92gat), .ZN(new_n561_));
  NOR3_X1   g360(.A1(new_n560_), .A2(new_n561_), .A3(KEYINPUT9), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n562_), .B1(new_n551_), .B2(KEYINPUT9), .ZN(new_n563_));
  AND2_X1   g362(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n564_));
  NOR2_X1   g363(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT64), .B(G106gat), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT65), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n566_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n568_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n559_), .B(new_n563_), .C1(new_n569_), .C2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n553_), .A2(new_n558_), .A3(new_n571_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n572_), .A2(new_n508_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G232gat), .A2(G233gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(KEYINPUT69), .B(KEYINPUT35), .Z(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n578_), .B1(new_n572_), .B2(new_n521_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n573_), .A2(new_n579_), .ZN(new_n580_));
  OAI211_X1 g379(.A(KEYINPUT70), .B(new_n578_), .C1(new_n572_), .C2(new_n521_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n576_), .A2(new_n577_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n580_), .A2(new_n583_), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n581_), .B(new_n582_), .C1(new_n573_), .C2(new_n579_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G190gat), .B(G218gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G134gat), .B(G162gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n589_), .B(KEYINPUT36), .Z(new_n590_));
  XOR2_X1   g389(.A(new_n590_), .B(KEYINPUT71), .Z(new_n591_));
  OAI21_X1  g390(.A(KEYINPUT73), .B1(new_n586_), .B2(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n589_), .A2(KEYINPUT36), .ZN(new_n593_));
  AND3_X1   g392(.A1(new_n584_), .A2(new_n585_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT37), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n591_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT73), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n592_), .A2(new_n595_), .A3(new_n596_), .A4(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(KEYINPUT37), .B1(new_n594_), .B2(new_n597_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT72), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT72), .ZN(new_n603_));
  OAI211_X1 g402(.A(new_n603_), .B(KEYINPUT37), .C1(new_n594_), .C2(new_n597_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n600_), .A2(new_n602_), .A3(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT17), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G127gat), .B(G155gat), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n607_), .B(KEYINPUT16), .Z(new_n608_));
  XNOR2_X1  g407(.A(G183gat), .B(G211gat), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n607_), .B(KEYINPUT16), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(new_n609_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n606_), .B1(new_n611_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT74), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n517_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n613_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n612_), .A2(new_n609_), .ZN(new_n618_));
  OAI21_X1  g417(.A(KEYINPUT17), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n619_), .A2(KEYINPUT74), .A3(new_n515_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n616_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(G231gat), .A2(G233gat), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n616_), .A2(new_n620_), .A3(G231gat), .A4(G233gat), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G57gat), .B(G64gat), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(KEYINPUT11), .ZN(new_n627_));
  XOR2_X1   g426(.A(G71gat), .B(G78gat), .Z(new_n628_));
  NOR2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n627_), .A2(new_n628_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n626_), .A2(KEYINPUT11), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n630_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n625_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n623_), .A2(new_n633_), .A3(new_n624_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n613_), .A2(new_n611_), .A3(new_n606_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n635_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n605_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n572_), .A2(new_n634_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n633_), .A2(new_n553_), .A3(new_n558_), .A4(new_n571_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(KEYINPUT12), .A3(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT12), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n572_), .A2(new_n643_), .A3(new_n634_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(G230gat), .A2(G233gat), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n646_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(G120gat), .B(G148gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT5), .ZN(new_n651_));
  XNOR2_X1  g450(.A(G176gat), .B(G204gat), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n651_), .B(new_n652_), .Z(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n647_), .A2(new_n649_), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n646_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n656_), .B1(new_n642_), .B2(new_n644_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n653_), .B1(new_n657_), .B2(new_n648_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT13), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n659_), .A2(KEYINPUT67), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n655_), .A2(new_n658_), .A3(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(KEYINPUT67), .B(KEYINPUT13), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n663_), .B1(new_n655_), .B2(new_n658_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n639_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n537_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n414_), .ZN(new_n668_));
  NOR3_X1   g467(.A1(new_n667_), .A2(G1gat), .A3(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n592_), .A2(new_n595_), .A3(new_n599_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n504_), .A2(new_n673_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n533_), .A2(new_n535_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n675_), .B1(new_n662_), .B2(new_n664_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT101), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT101), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n678_), .B(new_n675_), .C1(new_n662_), .C2(new_n664_), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n677_), .A2(new_n638_), .A3(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n674_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(new_n414_), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n683_), .A2(KEYINPUT102), .A3(G1gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(KEYINPUT102), .B1(new_n683_), .B2(G1gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n671_), .B1(new_n684_), .B2(new_n685_), .ZN(G1324gat));
  INV_X1    g485(.A(new_n667_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n345_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(new_n511_), .A3(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n682_), .A2(new_n688_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT39), .ZN(new_n691_));
  AND4_X1   g490(.A1(KEYINPUT103), .A2(new_n690_), .A3(new_n691_), .A4(G8gat), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n511_), .B1(new_n693_), .B2(KEYINPUT39), .ZN(new_n694_));
  AOI22_X1  g493(.A1(new_n690_), .A2(new_n694_), .B1(KEYINPUT103), .B2(new_n691_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n689_), .B1(new_n692_), .B2(new_n695_), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g496(.A(G15gat), .B1(new_n681_), .B2(new_n481_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT41), .Z(new_n699_));
  NAND3_X1  g498(.A1(new_n687_), .A2(new_n453_), .A3(new_n502_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1326gat));
  INV_X1    g500(.A(new_n445_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G22gat), .B1(new_n681_), .B2(new_n702_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT42), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n702_), .A2(G22gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n704_), .B1(new_n667_), .B2(new_n705_), .ZN(G1327gat));
  INV_X1    g505(.A(new_n638_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n673_), .A2(new_n707_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n708_), .A2(new_n665_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n537_), .A2(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(G29gat), .B1(new_n710_), .B2(new_n414_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n677_), .A2(new_n707_), .A3(new_n679_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT104), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT104), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n677_), .A2(new_n715_), .A3(new_n707_), .A4(new_n679_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n345_), .A2(new_n485_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n501_), .A2(new_n503_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n720_));
  INV_X1    g519(.A(new_n605_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n719_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(KEYINPUT43), .B1(new_n504_), .B2(new_n605_), .ZN(new_n723_));
  AOI221_X4 g522(.A(new_n712_), .B1(new_n714_), .B2(new_n716_), .C1(new_n722_), .C2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n723_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n714_), .A2(new_n716_), .ZN(new_n726_));
  AOI21_X1  g525(.A(KEYINPUT44), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n724_), .A2(new_n727_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n414_), .A2(G29gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n711_), .B1(new_n728_), .B2(new_n729_), .ZN(G1328gat));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n731_));
  INV_X1    g530(.A(G36gat), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n537_), .A2(new_n732_), .A3(new_n688_), .A4(new_n709_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n733_), .B(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n720_), .B1(new_n719_), .B2(new_n721_), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n504_), .A2(KEYINPUT43), .A3(new_n605_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n726_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(new_n712_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n725_), .A2(KEYINPUT44), .A3(new_n726_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(new_n688_), .A3(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n735_), .B1(new_n741_), .B2(G36gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n731_), .B1(new_n742_), .B2(KEYINPUT105), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT105), .ZN(new_n744_));
  AOI211_X1 g543(.A(new_n744_), .B(new_n735_), .C1(new_n741_), .C2(G36gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(KEYINPUT106), .B1(new_n743_), .B2(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n732_), .B1(new_n728_), .B2(new_n688_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n744_), .B1(new_n747_), .B2(new_n735_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT106), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n742_), .A2(KEYINPUT105), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n748_), .A2(new_n749_), .A3(new_n731_), .A4(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n742_), .A2(KEYINPUT46), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n746_), .A2(new_n751_), .A3(new_n752_), .ZN(G1329gat));
  AOI21_X1  g552(.A(new_n459_), .B1(new_n468_), .B2(new_n478_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n728_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT107), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n728_), .A2(KEYINPUT107), .A3(new_n754_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n710_), .A2(new_n502_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(new_n459_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n757_), .A2(new_n758_), .A3(new_n760_), .ZN(new_n761_));
  XOR2_X1   g560(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n762_));
  XNOR2_X1  g561(.A(new_n761_), .B(new_n762_), .ZN(G1330gat));
  NAND2_X1  g562(.A1(new_n728_), .A2(new_n445_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(G50gat), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n702_), .A2(G50gat), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT109), .Z(new_n767_));
  NAND2_X1  g566(.A1(new_n710_), .A2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n765_), .A2(new_n768_), .ZN(G1331gat));
  NOR2_X1   g568(.A1(new_n504_), .A2(new_n675_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n664_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n655_), .A2(new_n658_), .A3(new_n661_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n639_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n770_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(G57gat), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n776_), .A2(new_n777_), .A3(new_n414_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n638_), .A2(new_n536_), .ZN(new_n779_));
  NOR4_X1   g578(.A1(new_n504_), .A2(new_n673_), .A3(new_n773_), .A4(new_n779_), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n780_), .A2(new_n414_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n778_), .B1(new_n781_), .B2(new_n777_), .ZN(G1332gat));
  INV_X1    g581(.A(G64gat), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(new_n780_), .B2(new_n688_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n784_), .B(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n688_), .A2(new_n783_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT111), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n786_), .B1(new_n775_), .B2(new_n788_), .ZN(G1333gat));
  INV_X1    g588(.A(G71gat), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n790_), .B1(new_n780_), .B2(new_n502_), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT49), .Z(new_n792_));
  NAND3_X1  g591(.A1(new_n776_), .A2(new_n790_), .A3(new_n502_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(G1334gat));
  INV_X1    g593(.A(G78gat), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n780_), .B2(new_n445_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT113), .ZN(new_n797_));
  XOR2_X1   g596(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n798_));
  XNOR2_X1  g597(.A(new_n797_), .B(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n445_), .A2(new_n795_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n799_), .B1(new_n775_), .B2(new_n800_), .ZN(G1335gat));
  NAND4_X1  g600(.A1(new_n725_), .A2(new_n707_), .A3(new_n665_), .A4(new_n536_), .ZN(new_n802_));
  OAI21_X1  g601(.A(G85gat), .B1(new_n802_), .B2(new_n668_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n708_), .A2(new_n773_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n770_), .A2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n806_), .A2(new_n560_), .A3(new_n414_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n803_), .A2(new_n807_), .ZN(G1336gat));
  OAI21_X1  g607(.A(G92gat), .B1(new_n802_), .B2(new_n345_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n806_), .A2(new_n561_), .A3(new_n688_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(G1337gat));
  OAI21_X1  g610(.A(G99gat), .B1(new_n802_), .B2(new_n481_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n806_), .A2(new_n566_), .A3(new_n483_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(KEYINPUT51), .ZN(G1338gat));
  AND3_X1   g614(.A1(new_n806_), .A2(new_n567_), .A3(new_n445_), .ZN(new_n816_));
  OAI21_X1  g615(.A(G106gat), .B1(new_n802_), .B2(new_n702_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT52), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n819_), .B(G106gat), .C1(new_n802_), .C2(new_n702_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n816_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n822_));
  XOR2_X1   g621(.A(new_n821_), .B(new_n822_), .Z(G1339gat));
  INV_X1    g622(.A(new_n484_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n345_), .A2(new_n414_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n665_), .B2(new_n779_), .ZN(new_n828_));
  AND2_X1   g627(.A1(new_n638_), .A2(new_n536_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n773_), .A2(new_n829_), .A3(KEYINPUT115), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n605_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT54), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n831_), .A2(new_n834_), .A3(new_n605_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT58), .ZN(new_n837_));
  INV_X1    g636(.A(new_n532_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n523_), .A2(new_n519_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT116), .B1(new_n839_), .B2(new_n530_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n519_), .B1(new_n517_), .B2(new_n507_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n840_), .B1(new_n516_), .B2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n839_), .A2(KEYINPUT116), .A3(new_n530_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n838_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n844_), .A2(new_n655_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n642_), .A2(new_n656_), .A3(new_n644_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n647_), .A2(KEYINPUT55), .A3(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT55), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n654_), .B1(new_n657_), .B2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n847_), .A2(KEYINPUT56), .A3(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT56), .B1(new_n847_), .B2(new_n849_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n845_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n605_), .B1(new_n837_), .B2(new_n853_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n845_), .B(KEYINPUT58), .C1(new_n852_), .C2(new_n851_), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n655_), .B(new_n675_), .C1(new_n851_), .C2(new_n852_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n655_), .A2(new_n658_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n844_), .A2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n673_), .B1(new_n856_), .B2(new_n858_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  AOI22_X1  g660(.A1(new_n854_), .A2(new_n855_), .B1(new_n859_), .B2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n856_), .A2(new_n858_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n672_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n860_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n638_), .B1(new_n862_), .B2(new_n865_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n824_), .B(new_n826_), .C1(new_n836_), .C2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(G113gat), .B1(new_n868_), .B2(new_n675_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT59), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n867_), .A2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n859_), .A2(new_n861_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n853_), .A2(new_n837_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n873_), .A2(new_n721_), .A3(new_n855_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n865_), .A2(new_n872_), .A3(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n707_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n833_), .A2(new_n835_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n825_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n878_), .A2(KEYINPUT59), .A3(new_n824_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n871_), .A2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n675_), .A2(G113gat), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(KEYINPUT118), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n869_), .B1(new_n880_), .B2(new_n882_), .ZN(G1340gat));
  INV_X1    g682(.A(KEYINPUT60), .ZN(new_n884_));
  AOI21_X1  g683(.A(G120gat), .B1(new_n665_), .B2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(KEYINPUT119), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n887_), .B1(new_n884_), .B2(G120gat), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n868_), .B(new_n886_), .C1(new_n885_), .C2(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n773_), .B1(new_n871_), .B2(new_n879_), .ZN(new_n890_));
  INV_X1    g689(.A(G120gat), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n889_), .B1(new_n890_), .B2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(KEYINPUT120), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT120), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n894_), .B(new_n889_), .C1(new_n890_), .C2(new_n891_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n893_), .A2(new_n895_), .ZN(G1341gat));
  INV_X1    g695(.A(G127gat), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n868_), .A2(new_n897_), .A3(new_n638_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n707_), .B1(new_n871_), .B2(new_n879_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(new_n897_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  OAI211_X1 g701(.A(KEYINPUT121), .B(new_n898_), .C1(new_n899_), .C2(new_n897_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1342gat));
  INV_X1    g703(.A(G134gat), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n868_), .A2(new_n905_), .A3(new_n673_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n605_), .B1(new_n871_), .B2(new_n879_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n907_), .B2(new_n905_), .ZN(G1343gat));
  AOI211_X1 g707(.A(new_n482_), .B(new_n825_), .C1(new_n876_), .C2(new_n877_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(new_n675_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n665_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(KEYINPUT122), .B(G148gat), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n912_), .B(new_n913_), .ZN(G1345gat));
  XNOR2_X1  g713(.A(KEYINPUT61), .B(G155gat), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n482_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n878_), .A2(new_n917_), .A3(new_n638_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(KEYINPUT123), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT123), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n909_), .A2(new_n920_), .A3(new_n638_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT124), .ZN(new_n922_));
  AND3_X1   g721(.A1(new_n919_), .A2(new_n921_), .A3(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n922_), .B1(new_n919_), .B2(new_n921_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n916_), .B1(new_n923_), .B2(new_n924_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n918_), .A2(KEYINPUT123), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n920_), .B1(new_n909_), .B2(new_n638_), .ZN(new_n927_));
  OAI21_X1  g726(.A(KEYINPUT124), .B1(new_n926_), .B2(new_n927_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n919_), .A2(new_n921_), .A3(new_n922_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n928_), .A2(new_n915_), .A3(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n925_), .A2(new_n930_), .ZN(G1346gat));
  INV_X1    g730(.A(new_n909_), .ZN(new_n932_));
  OAI21_X1  g731(.A(G162gat), .B1(new_n932_), .B2(new_n605_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n909_), .A2(new_n352_), .A3(new_n673_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(G1347gat));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n345_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n937_));
  NOR3_X1   g736(.A1(new_n414_), .A2(new_n445_), .A3(new_n481_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n937_), .A2(new_n938_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n939_), .A2(new_n536_), .ZN(new_n940_));
  OAI21_X1  g739(.A(new_n936_), .B1(new_n940_), .B2(new_n202_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n212_), .ZN(new_n942_));
  OAI211_X1 g741(.A(KEYINPUT62), .B(G169gat), .C1(new_n939_), .C2(new_n536_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n941_), .A2(new_n942_), .A3(new_n943_), .ZN(G1348gat));
  NOR2_X1   g743(.A1(new_n939_), .A2(new_n773_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(new_n206_), .ZN(G1349gat));
  NOR2_X1   g745(.A1(new_n939_), .A2(new_n707_), .ZN(new_n947_));
  INV_X1    g746(.A(new_n227_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n947_), .A2(new_n948_), .ZN(new_n949_));
  OR2_X1    g748(.A1(new_n949_), .A2(KEYINPUT125), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n949_), .A2(KEYINPUT125), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n947_), .A2(G183gat), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n950_), .B1(new_n951_), .B2(new_n952_), .ZN(G1350gat));
  OAI21_X1  g752(.A(G190gat), .B1(new_n939_), .B2(new_n605_), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n673_), .A2(new_n290_), .A3(new_n289_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n954_), .B1(new_n939_), .B2(new_n955_), .ZN(G1351gat));
  NOR2_X1   g755(.A1(new_n482_), .A2(new_n414_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n937_), .A2(new_n957_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n958_), .A2(new_n536_), .ZN(new_n959_));
  XNOR2_X1  g758(.A(new_n959_), .B(new_n258_), .ZN(G1352gat));
  NOR2_X1   g759(.A1(new_n958_), .A2(new_n773_), .ZN(new_n961_));
  XNOR2_X1  g760(.A(new_n961_), .B(new_n251_), .ZN(G1353gat));
  NOR2_X1   g761(.A1(new_n958_), .A2(new_n707_), .ZN(new_n963_));
  NOR3_X1   g762(.A1(new_n963_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n964_));
  XOR2_X1   g763(.A(KEYINPUT63), .B(G211gat), .Z(new_n965_));
  AOI21_X1  g764(.A(new_n964_), .B1(new_n963_), .B2(new_n965_), .ZN(G1354gat));
  INV_X1    g765(.A(new_n958_), .ZN(new_n967_));
  AOI21_X1  g766(.A(G218gat), .B1(new_n967_), .B2(new_n673_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n721_), .A2(G218gat), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n969_), .B(KEYINPUT126), .ZN(new_n970_));
  AOI21_X1  g769(.A(new_n968_), .B1(new_n967_), .B2(new_n970_), .ZN(G1355gat));
endmodule


