//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 1 0 1 1 1 1 1 1 0 0 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n912_, new_n913_, new_n915_, new_n916_, new_n917_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_;
  INV_X1    g000(.A(KEYINPUT38), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n203_), .B(KEYINPUT94), .Z(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT19), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT22), .B(G169gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT95), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G176gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT79), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT82), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n215_), .B1(new_n216_), .B2(KEYINPUT23), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT81), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n216_), .B(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n217_), .B1(new_n219_), .B2(KEYINPUT23), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n216_), .B(KEYINPUT81), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT23), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(new_n215_), .A3(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n220_), .A2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G183gat), .A2(G190gat), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n211_), .B(new_n214_), .C1(new_n224_), .C2(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n227_), .B1(new_n221_), .B2(KEYINPUT23), .ZN(new_n228_));
  NOR3_X1   g027(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n229_), .B1(new_n231_), .B2(new_n212_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT26), .B(G190gat), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  XOR2_X1   g033(.A(KEYINPUT25), .B(G183gat), .Z(new_n235_));
  OAI211_X1 g034(.A(new_n228_), .B(new_n232_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n226_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G211gat), .B(G218gat), .ZN(new_n238_));
  XOR2_X1   g037(.A(G197gat), .B(G204gat), .Z(new_n239_));
  OAI21_X1  g038(.A(new_n238_), .B1(new_n239_), .B2(KEYINPUT21), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(KEYINPUT21), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT20), .B1(new_n237_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n224_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n214_), .A2(new_n231_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT78), .ZN(new_n247_));
  INV_X1    g046(.A(G183gat), .ZN(new_n248_));
  OR3_X1    g047(.A1(new_n247_), .A2(new_n248_), .A3(KEYINPUT25), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT25), .B1(new_n247_), .B2(new_n248_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(new_n233_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n246_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT80), .ZN(new_n253_));
  INV_X1    g052(.A(new_n229_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT80), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n246_), .A2(new_n251_), .A3(new_n255_), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n245_), .A2(new_n253_), .A3(new_n254_), .A4(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n228_), .B1(G183gat), .B2(G190gat), .ZN(new_n258_));
  INV_X1    g057(.A(G169gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT22), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n259_), .B1(new_n260_), .B2(KEYINPUT83), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT84), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n261_), .B1(new_n262_), .B2(KEYINPUT22), .ZN(new_n263_));
  NOR4_X1   g062(.A1(new_n260_), .A2(new_n259_), .A3(KEYINPUT83), .A4(KEYINPUT84), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n210_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n258_), .A2(new_n214_), .A3(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n242_), .B1(new_n257_), .B2(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n206_), .B1(new_n244_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n237_), .A2(new_n243_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n257_), .A2(new_n266_), .A3(new_n242_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n269_), .A2(new_n270_), .A3(KEYINPUT20), .A4(new_n205_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(G8gat), .B(G36gat), .Z(new_n273_));
  XNOR2_X1  g072(.A(G64gat), .B(G92gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n272_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n277_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n268_), .A2(new_n279_), .A3(new_n271_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n278_), .A2(KEYINPUT97), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT97), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n272_), .A2(new_n282_), .A3(new_n277_), .ZN(new_n283_));
  XOR2_X1   g082(.A(KEYINPUT103), .B(KEYINPUT27), .Z(new_n284_));
  NAND3_X1  g083(.A1(new_n281_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n205_), .B1(new_n244_), .B2(new_n267_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n269_), .A2(KEYINPUT20), .A3(new_n270_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n286_), .B1(new_n287_), .B2(new_n205_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n279_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n289_), .A2(KEYINPUT27), .A3(new_n278_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n285_), .A2(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(G78gat), .B(G106gat), .Z(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT89), .ZN(new_n294_));
  INV_X1    g093(.A(G228gat), .ZN(new_n295_));
  INV_X1    g094(.A(G233gat), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT90), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(G141gat), .A2(G148gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT3), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G141gat), .A2(G148gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT2), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  AND2_X1   g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306_));
  NOR2_X1   g105(.A1(G155gat), .A2(G162gat), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT1), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n301_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n306_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n311_));
  AOI22_X1  g110(.A1(new_n305_), .A2(new_n308_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT29), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n294_), .B(new_n300_), .C1(new_n312_), .C2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n305_), .A2(new_n308_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n310_), .A2(new_n311_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n317_), .A2(KEYINPUT90), .A3(KEYINPUT29), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n242_), .B1(new_n314_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(KEYINPUT89), .B1(new_n317_), .B2(KEYINPUT29), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(new_n243_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n297_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n293_), .B1(new_n320_), .B2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n297_), .B1(new_n321_), .B2(new_n243_), .ZN(new_n326_));
  NOR3_X1   g125(.A1(new_n326_), .A2(new_n319_), .A3(new_n292_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G22gat), .B(G50gat), .ZN(new_n329_));
  OR3_X1    g128(.A1(new_n317_), .A2(KEYINPUT29), .A3(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n329_), .B1(new_n317_), .B2(KEYINPUT29), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n331_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT91), .B1(new_n328_), .B2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n292_), .B1(new_n326_), .B2(new_n319_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT92), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n337_), .B1(new_n327_), .B2(new_n338_), .ZN(new_n339_));
  OAI211_X1 g138(.A(KEYINPUT92), .B(new_n292_), .C1(new_n326_), .C2(new_n319_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(new_n335_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT91), .ZN(new_n342_));
  OAI221_X1 g141(.A(new_n342_), .B1(new_n333_), .B2(new_n334_), .C1(new_n325_), .C2(new_n327_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n336_), .A2(new_n341_), .A3(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT93), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT93), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n336_), .A2(new_n341_), .A3(new_n346_), .A4(new_n343_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n291_), .B1(new_n345_), .B2(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT86), .B(G113gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(G120gat), .ZN(new_n350_));
  XOR2_X1   g149(.A(G127gat), .B(G134gat), .Z(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(G120gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n349_), .B(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n351_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n352_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(new_n317_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n312_), .A2(new_n352_), .A3(new_n356_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n358_), .A2(KEYINPUT4), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G225gat), .A2(G233gat), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT4), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n357_), .A2(new_n363_), .A3(new_n317_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n360_), .A2(new_n362_), .A3(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT98), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n358_), .A2(new_n359_), .A3(new_n361_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n360_), .A2(KEYINPUT98), .A3(new_n362_), .A4(new_n364_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  XOR2_X1   g169(.A(G1gat), .B(G29gat), .Z(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT100), .ZN(new_n372_));
  XOR2_X1   g171(.A(G57gat), .B(G85gat), .Z(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n370_), .A2(new_n377_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .A4(new_n376_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n345_), .A2(new_n347_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n281_), .A2(new_n283_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n379_), .B(KEYINPUT33), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n358_), .A2(new_n359_), .A3(new_n362_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n360_), .A2(new_n361_), .A3(new_n364_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n377_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n384_), .A2(new_n385_), .A3(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n277_), .A2(KEYINPUT32), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT101), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n272_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT102), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n288_), .A2(KEYINPUT32), .A3(new_n277_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n272_), .A2(KEYINPUT102), .A3(new_n391_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n380_), .A2(new_n394_), .A3(new_n395_), .A4(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n389_), .A2(new_n397_), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n348_), .A2(new_n381_), .B1(new_n383_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT30), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n257_), .A2(new_n400_), .A3(new_n266_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n400_), .B1(new_n257_), .B2(new_n266_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n404_), .A2(KEYINPUT85), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n357_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n352_), .B(new_n356_), .C1(new_n404_), .C2(KEYINPUT85), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n257_), .A2(new_n266_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT30), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n410_), .A2(KEYINPUT85), .A3(new_n401_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT31), .ZN(new_n412_));
  XOR2_X1   g211(.A(G71gat), .B(G99gat), .Z(new_n413_));
  XNOR2_X1  g212(.A(G15gat), .B(G43gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G227gat), .A2(G233gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  AND3_X1   g216(.A1(new_n411_), .A2(new_n412_), .A3(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n412_), .B1(new_n411_), .B2(new_n417_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n408_), .A2(new_n420_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n406_), .B(new_n407_), .C1(new_n418_), .C2(new_n419_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n421_), .A2(KEYINPUT87), .A3(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT87), .B1(new_n421_), .B2(new_n422_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT104), .B1(new_n399_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n383_), .A2(new_n398_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n285_), .A2(new_n290_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n382_), .A2(new_n428_), .A3(new_n381_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT104), .ZN(new_n431_));
  INV_X1    g230(.A(new_n425_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n382_), .A2(new_n291_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n421_), .A2(new_n422_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n435_), .A2(new_n380_), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n426_), .A2(new_n433_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT67), .ZN(new_n438_));
  INV_X1    g237(.A(G99gat), .ZN(new_n439_));
  INV_X1    g238(.A(G106gat), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n438_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT7), .ZN(new_n442_));
  AND3_X1   g241(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n443_));
  AOI21_X1  g242(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT7), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n438_), .A2(new_n446_), .A3(new_n439_), .A4(new_n440_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n442_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(G92gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(G85gat), .ZN(new_n450_));
  INV_X1    g249(.A(G85gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(G92gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n448_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT8), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT8), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n448_), .A2(new_n456_), .A3(new_n453_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  NOR3_X1   g257(.A1(new_n449_), .A2(KEYINPUT65), .A3(KEYINPUT9), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT65), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n460_), .A2(G92gat), .ZN(new_n461_));
  OAI21_X1  g260(.A(G85gat), .B1(new_n459_), .B2(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n451_), .A2(G92gat), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n449_), .A2(G85gat), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT9), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT66), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n462_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT9), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n460_), .A2(new_n468_), .A3(G92gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n449_), .A2(KEYINPUT65), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n451_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n468_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT66), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n467_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT10), .B(G99gat), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n445_), .B1(G106gat), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(KEYINPUT69), .B1(new_n474_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT69), .ZN(new_n479_));
  AOI211_X1 g278(.A(new_n479_), .B(new_n476_), .C1(new_n467_), .C2(new_n473_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n458_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(G57gat), .ZN(new_n482_));
  INV_X1    g281(.A(G64gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT11), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G57gat), .A2(G64gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n484_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G71gat), .A2(G78gat), .ZN(new_n488_));
  INV_X1    g287(.A(G71gat), .ZN(new_n489_));
  INV_X1    g288(.A(G78gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n487_), .A2(new_n488_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT68), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n485_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT68), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n487_), .A2(new_n495_), .A3(new_n488_), .A4(new_n491_), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n493_), .A2(new_n494_), .A3(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n494_), .B1(new_n493_), .B2(new_n496_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT12), .ZN(new_n499_));
  NOR3_X1   g298(.A1(new_n497_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n481_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G230gat), .A2(G233gat), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n502_), .B(KEYINPUT64), .Z(new_n503_));
  INV_X1    g302(.A(new_n498_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n493_), .A2(new_n494_), .A3(new_n496_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  AOI22_X1  g305(.A1(new_n455_), .A2(new_n457_), .B1(new_n474_), .B2(new_n477_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n499_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n507_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n501_), .A2(new_n503_), .A3(new_n508_), .A4(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT70), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n497_), .A2(new_n498_), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n467_), .A2(new_n473_), .ZN(new_n513_));
  AND3_X1   g312(.A1(new_n448_), .A2(new_n456_), .A3(new_n453_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n456_), .B1(new_n448_), .B2(new_n453_), .ZN(new_n515_));
  OAI22_X1  g314(.A1(new_n513_), .A2(new_n476_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT12), .B1(new_n512_), .B2(new_n516_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n512_), .A2(new_n516_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT70), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n519_), .A2(new_n520_), .A3(new_n503_), .A4(new_n501_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n511_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n503_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n506_), .A2(new_n507_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n523_), .B1(new_n524_), .B2(new_n518_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n522_), .A2(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(G120gat), .B(G148gat), .Z(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(G204gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT5), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(new_n210_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n526_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n522_), .A2(new_n525_), .A3(new_n530_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT71), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT13), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n534_), .A2(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n534_), .B1(new_n537_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G1gat), .B(G8gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT76), .ZN(new_n543_));
  OR2_X1    g342(.A1(G15gat), .A2(G22gat), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G15gat), .A2(G22gat), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G1gat), .A2(G8gat), .ZN(new_n546_));
  AOI22_X1  g345(.A1(new_n544_), .A2(new_n545_), .B1(KEYINPUT14), .B2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n543_), .B(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G29gat), .B(G36gat), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n549_), .A2(G43gat), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(G43gat), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(G50gat), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(G50gat), .B1(new_n550_), .B2(new_n551_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n548_), .B(new_n555_), .Z(new_n556_));
  NAND3_X1  g355(.A1(new_n556_), .A2(G229gat), .A3(G233gat), .ZN(new_n557_));
  OR3_X1    g356(.A1(new_n548_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT15), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n559_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n549_), .B(G43gat), .ZN(new_n561_));
  INV_X1    g360(.A(G50gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n563_), .A2(KEYINPUT15), .A3(new_n552_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n560_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(new_n548_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G229gat), .A2(G233gat), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n558_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n557_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G113gat), .B(G141gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(new_n259_), .ZN(new_n571_));
  INV_X1    g370(.A(G197gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n569_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n573_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n557_), .A2(new_n568_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n541_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT37), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G232gat), .A2(G233gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT34), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT35), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT72), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT74), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n581_), .A2(KEYINPUT35), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(new_n507_), .B2(new_n555_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT73), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n481_), .A2(new_n587_), .A3(new_n565_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n587_), .B1(new_n481_), .B2(new_n565_), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n584_), .B(new_n586_), .C1(new_n588_), .C2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n583_), .A2(KEYINPUT74), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(G134gat), .ZN(new_n594_));
  INV_X1    g393(.A(G162gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT36), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n514_), .A2(new_n515_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n479_), .B1(new_n513_), .B2(new_n476_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n474_), .A2(KEYINPUT69), .A3(new_n477_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n599_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NOR3_X1   g401(.A1(new_n553_), .A2(new_n559_), .A3(new_n554_), .ZN(new_n603_));
  AOI21_X1  g402(.A(KEYINPUT15), .B1(new_n563_), .B2(new_n552_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(KEYINPUT73), .B1(new_n602_), .B2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n481_), .A2(new_n587_), .A3(new_n565_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n591_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n608_), .A2(new_n609_), .A3(new_n584_), .A4(new_n586_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n592_), .A2(new_n598_), .A3(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n592_), .A2(KEYINPUT75), .A3(new_n610_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n596_), .A2(new_n597_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n611_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n612_), .B1(new_n613_), .B2(new_n611_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n579_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n592_), .A2(new_n610_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n613_), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n617_), .B(KEYINPUT75), .C1(new_n618_), .C2(new_n598_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n611_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(KEYINPUT37), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n616_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G231gat), .A2(G233gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n548_), .B(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(new_n506_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT16), .B(G183gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(G211gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G127gat), .B(G155gat), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n627_), .B(new_n628_), .Z(new_n629_));
  INV_X1    g428(.A(KEYINPUT17), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n629_), .A2(new_n630_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n625_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n633_), .B1(new_n631_), .B2(new_n625_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT77), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n622_), .A2(new_n635_), .ZN(new_n636_));
  NOR4_X1   g435(.A1(new_n437_), .A2(G1gat), .A3(new_n578_), .A4(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT105), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n637_), .A2(new_n638_), .A3(new_n380_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n638_), .B1(new_n637_), .B2(new_n380_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n202_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n641_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n643_), .A2(KEYINPUT38), .A3(new_n639_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n434_), .A2(new_n436_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n431_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n646_));
  AOI211_X1 g445(.A(KEYINPUT104), .B(new_n425_), .C1(new_n427_), .C2(new_n429_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n645_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n578_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n619_), .A2(new_n620_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n648_), .A2(new_n649_), .A3(new_n635_), .A4(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(G1gat), .B1(new_n652_), .B2(new_n381_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n642_), .A2(new_n644_), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT106), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n642_), .A2(new_n644_), .A3(KEYINPUT106), .A4(new_n653_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1324gat));
  XNOR2_X1  g457(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT39), .ZN(new_n661_));
  OAI211_X1 g460(.A(new_n661_), .B(G8gat), .C1(new_n652_), .C2(new_n428_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT108), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n426_), .A2(new_n433_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n650_), .B1(new_n665_), .B2(new_n645_), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n666_), .A2(new_n649_), .A3(new_n635_), .A4(new_n291_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n667_), .A2(KEYINPUT108), .A3(new_n661_), .A4(G8gat), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n664_), .A2(new_n668_), .ZN(new_n669_));
  AOI211_X1 g468(.A(KEYINPUT107), .B(new_n661_), .C1(new_n667_), .C2(G8gat), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT107), .ZN(new_n671_));
  OAI21_X1  g470(.A(G8gat), .B1(new_n652_), .B2(new_n428_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n672_), .B2(KEYINPUT39), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n669_), .A2(new_n670_), .A3(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n437_), .A2(new_n636_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(new_n649_), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n676_), .A2(G8gat), .A3(new_n428_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n660_), .B1(new_n674_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n677_), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n670_), .A2(new_n673_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n659_), .B(new_n679_), .C1(new_n680_), .C2(new_n669_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n678_), .A2(new_n681_), .ZN(G1325gat));
  OAI21_X1  g481(.A(G15gat), .B1(new_n652_), .B2(new_n432_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT41), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n683_), .B(new_n684_), .ZN(new_n685_));
  OR3_X1    g484(.A1(new_n676_), .A2(G15gat), .A3(new_n432_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT110), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(G1326gat));
  XNOR2_X1  g488(.A(new_n382_), .B(KEYINPUT111), .ZN(new_n690_));
  OAI21_X1  g489(.A(G22gat), .B1(new_n652_), .B2(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT42), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n690_), .A2(G22gat), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n692_), .B1(new_n676_), .B2(new_n693_), .ZN(G1327gat));
  NAND2_X1  g493(.A1(new_n648_), .A2(new_n650_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n578_), .A2(new_n635_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G29gat), .B1(new_n698_), .B2(new_n380_), .ZN(new_n699_));
  OAI21_X1  g498(.A(KEYINPUT43), .B1(new_n437_), .B2(new_n622_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n701_));
  INV_X1    g500(.A(new_n622_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n648_), .A2(new_n701_), .A3(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n700_), .A2(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT44), .B1(new_n704_), .B2(new_n696_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706_));
  AOI211_X1 g505(.A(new_n706_), .B(new_n697_), .C1(new_n700_), .C2(new_n703_), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n705_), .A2(new_n707_), .A3(new_n381_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n699_), .B1(new_n708_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g508(.A(KEYINPUT112), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n710_), .A2(KEYINPUT46), .ZN(new_n711_));
  INV_X1    g510(.A(G36gat), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n705_), .A2(new_n707_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(new_n291_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n698_), .A2(new_n712_), .A3(new_n291_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT45), .Z(new_n716_));
  OAI21_X1  g515(.A(new_n711_), .B1(new_n714_), .B2(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n715_), .B(KEYINPUT45), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n705_), .A2(new_n707_), .A3(new_n428_), .ZN(new_n719_));
  OAI221_X1 g518(.A(new_n718_), .B1(new_n710_), .B2(KEYINPUT46), .C1(new_n719_), .C2(new_n712_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n717_), .A2(new_n720_), .ZN(G1329gat));
  INV_X1    g520(.A(new_n705_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n704_), .A2(KEYINPUT44), .A3(new_n696_), .ZN(new_n723_));
  INV_X1    g522(.A(new_n435_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n724_), .A2(G43gat), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n722_), .A2(new_n723_), .A3(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(G43gat), .B1(new_n698_), .B2(new_n425_), .ZN(new_n727_));
  OAI21_X1  g526(.A(KEYINPUT47), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n713_), .B2(new_n725_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT47), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n728_), .A2(new_n731_), .ZN(G1330gat));
  NAND3_X1  g531(.A1(new_n722_), .A2(new_n382_), .A3(new_n723_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT113), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n713_), .A2(KEYINPUT113), .A3(new_n382_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(new_n736_), .A3(G50gat), .ZN(new_n737_));
  INV_X1    g536(.A(new_n690_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n698_), .A2(new_n562_), .A3(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(G1331gat));
  NOR2_X1   g539(.A1(new_n541_), .A2(new_n577_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n648_), .A2(new_n635_), .A3(new_n651_), .A4(new_n741_), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n742_), .A2(new_n482_), .A3(new_n381_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n675_), .A2(new_n741_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n380_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n743_), .B1(new_n745_), .B2(new_n482_), .ZN(G1332gat));
  OAI21_X1  g545(.A(G64gat), .B1(new_n742_), .B2(new_n428_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT114), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT114), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n749_), .B(G64gat), .C1(new_n742_), .C2(new_n428_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT48), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n744_), .A2(new_n483_), .A3(new_n291_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n748_), .A2(KEYINPUT48), .A3(new_n750_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n753_), .A2(new_n754_), .A3(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT115), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n753_), .A2(KEYINPUT115), .A3(new_n754_), .A4(new_n755_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(G1333gat));
  OAI21_X1  g559(.A(G71gat), .B1(new_n742_), .B2(new_n432_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT49), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n744_), .A2(new_n489_), .A3(new_n425_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1334gat));
  OAI21_X1  g563(.A(G78gat), .B1(new_n742_), .B2(new_n690_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT50), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n744_), .A2(new_n490_), .A3(new_n738_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(G1335gat));
  INV_X1    g567(.A(new_n635_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n741_), .A2(new_n769_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n695_), .A2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(G85gat), .B1(new_n771_), .B2(new_n380_), .ZN(new_n772_));
  XOR2_X1   g571(.A(new_n770_), .B(KEYINPUT116), .Z(new_n773_));
  NAND2_X1  g572(.A1(new_n704_), .A2(new_n773_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n774_), .A2(new_n381_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n772_), .B1(new_n775_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g575(.A(G92gat), .B1(new_n771_), .B2(new_n291_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n774_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n460_), .A2(G92gat), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n428_), .B1(new_n470_), .B2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n777_), .B1(new_n778_), .B2(new_n780_), .ZN(G1337gat));
  OAI21_X1  g580(.A(G99gat), .B1(new_n774_), .B2(new_n432_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n475_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n771_), .A2(new_n783_), .A3(new_n724_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g585(.A1(new_n771_), .A2(new_n440_), .A3(new_n382_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n704_), .A2(new_n382_), .A3(new_n773_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n788_), .A2(new_n789_), .A3(G106gat), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n788_), .B2(G106gat), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n787_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT53), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n794_), .B(new_n787_), .C1(new_n790_), .C2(new_n791_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(G1339gat));
  INV_X1    g595(.A(KEYINPUT117), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT55), .B1(new_n511_), .B2(new_n521_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n508_), .A2(new_n509_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n481_), .A2(new_n500_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n523_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(new_n510_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n531_), .B1(new_n798_), .B2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT56), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n556_), .A2(new_n567_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n558_), .A2(new_n566_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n806_), .B(new_n573_), .C1(new_n567_), .C2(new_n807_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n808_), .A2(new_n576_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT56), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n810_), .B(new_n531_), .C1(new_n798_), .C2(new_n803_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n805_), .A2(new_n533_), .A3(new_n809_), .A4(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT58), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n797_), .B1(new_n814_), .B2(new_n622_), .ZN(new_n815_));
  OR2_X1    g614(.A1(new_n812_), .A2(new_n813_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n812_), .A2(new_n813_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n817_), .A2(KEYINPUT117), .A3(new_n621_), .A4(new_n616_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n815_), .A2(new_n816_), .A3(new_n818_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n805_), .A2(new_n577_), .A3(new_n533_), .A4(new_n811_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n534_), .A2(new_n809_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n650_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT57), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n822_), .B(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n819_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n769_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n827_));
  INV_X1    g626(.A(new_n577_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n622_), .A2(new_n541_), .A3(new_n828_), .A4(new_n635_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n829_), .B(KEYINPUT54), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n826_), .A2(new_n827_), .A3(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n635_), .B1(new_n819_), .B2(new_n824_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n829_), .B(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT118), .B1(new_n832_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n831_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n434_), .A2(new_n380_), .A3(new_n724_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(G113gat), .B1(new_n838_), .B2(new_n577_), .ZN(new_n839_));
  OAI21_X1  g638(.A(KEYINPUT59), .B1(new_n836_), .B2(new_n837_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n826_), .A2(new_n830_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT59), .ZN(new_n842_));
  INV_X1    g641(.A(new_n837_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n841_), .A2(new_n842_), .A3(new_n843_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n840_), .A2(new_n844_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n845_), .A2(new_n577_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n839_), .B1(new_n846_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g646(.A(new_n541_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n840_), .A2(new_n848_), .A3(new_n844_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT119), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT119), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n840_), .A2(new_n851_), .A3(new_n848_), .A4(new_n844_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n850_), .A2(G120gat), .A3(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n353_), .B1(new_n541_), .B2(KEYINPUT60), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n838_), .B(new_n854_), .C1(KEYINPUT60), .C2(new_n353_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n853_), .A2(new_n855_), .ZN(G1341gat));
  AOI21_X1  g655(.A(G127gat), .B1(new_n838_), .B2(new_n635_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n845_), .A2(new_n635_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g658(.A(G134gat), .B1(new_n838_), .B2(new_n650_), .ZN(new_n860_));
  XOR2_X1   g659(.A(KEYINPUT120), .B(G134gat), .Z(new_n861_));
  NOR2_X1   g660(.A1(new_n622_), .A2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n860_), .B1(new_n845_), .B2(new_n862_), .ZN(G1343gat));
  NOR2_X1   g662(.A1(new_n425_), .A2(new_n383_), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n831_), .A2(new_n835_), .A3(new_n428_), .A4(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT121), .B1(new_n865_), .B2(new_n381_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n865_), .A2(KEYINPUT121), .A3(new_n381_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n577_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(G141gat), .ZN(new_n870_));
  INV_X1    g669(.A(G141gat), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n871_), .B(new_n577_), .C1(new_n867_), .C2(new_n868_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n872_), .ZN(G1344gat));
  OAI21_X1  g672(.A(new_n848_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(G148gat), .ZN(new_n875_));
  INV_X1    g674(.A(G148gat), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n876_), .B(new_n848_), .C1(new_n867_), .C2(new_n868_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n877_), .ZN(G1345gat));
  OAI21_X1  g677(.A(new_n635_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(KEYINPUT61), .B(G155gat), .ZN(new_n880_));
  XOR2_X1   g679(.A(new_n880_), .B(KEYINPUT122), .Z(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n881_), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n635_), .B(new_n883_), .C1(new_n867_), .C2(new_n868_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n882_), .A2(new_n884_), .ZN(G1346gat));
  OAI21_X1  g684(.A(new_n650_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n865_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n887_), .A2(new_n888_), .A3(new_n380_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n595_), .B1(new_n889_), .B2(new_n866_), .ZN(new_n890_));
  AOI22_X1  g689(.A1(new_n886_), .A2(new_n595_), .B1(new_n890_), .B2(new_n702_), .ZN(G1347gat));
  NOR2_X1   g690(.A1(new_n428_), .A2(new_n380_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n425_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n841_), .A2(new_n690_), .A3(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(G169gat), .B1(new_n895_), .B2(new_n828_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(KEYINPUT62), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n577_), .A2(new_n209_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(KEYINPUT123), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n897_), .B1(new_n895_), .B2(new_n899_), .ZN(G1348gat));
  INV_X1    g699(.A(KEYINPUT124), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n827_), .B1(new_n826_), .B2(new_n830_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n832_), .A2(new_n834_), .A3(KEYINPUT118), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n904_), .A2(new_n383_), .A3(new_n894_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n905_), .A2(new_n210_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n901_), .B1(new_n906_), .B2(new_n848_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n895_), .ZN(new_n908_));
  AOI21_X1  g707(.A(G176gat), .B1(new_n908_), .B2(new_n848_), .ZN(new_n909_));
  NOR4_X1   g708(.A1(new_n905_), .A2(KEYINPUT124), .A3(new_n210_), .A4(new_n541_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n907_), .A2(new_n909_), .A3(new_n910_), .ZN(G1349gat));
  AND3_X1   g710(.A1(new_n908_), .A2(new_n635_), .A3(new_n235_), .ZN(new_n912_));
  OR2_X1    g711(.A1(new_n905_), .A2(new_n769_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n248_), .ZN(G1350gat));
  OAI21_X1  g713(.A(G190gat), .B1(new_n895_), .B2(new_n622_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n650_), .A2(new_n233_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n895_), .B2(new_n916_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(KEYINPUT125), .ZN(G1351gat));
  INV_X1    g717(.A(KEYINPUT126), .ZN(new_n919_));
  NAND4_X1  g718(.A1(new_n904_), .A2(new_n919_), .A3(new_n864_), .A4(new_n892_), .ZN(new_n920_));
  NAND4_X1  g719(.A1(new_n831_), .A2(new_n835_), .A3(new_n864_), .A4(new_n892_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(KEYINPUT126), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n828_), .B1(new_n920_), .B2(new_n922_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(new_n572_), .ZN(G1352gat));
  NAND2_X1  g723(.A1(new_n920_), .A2(new_n922_), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n925_), .A2(G204gat), .A3(new_n848_), .ZN(new_n926_));
  AOI21_X1  g725(.A(G204gat), .B1(new_n925_), .B2(new_n848_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n926_), .A2(new_n927_), .ZN(G1353gat));
  NAND2_X1  g727(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n929_));
  AND2_X1   g728(.A1(new_n921_), .A2(KEYINPUT126), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n921_), .A2(KEYINPUT126), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n635_), .B(new_n929_), .C1(new_n930_), .C2(new_n931_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(KEYINPUT127), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n932_), .A2(new_n935_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n929_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n937_), .B1(new_n920_), .B2(new_n922_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n934_), .B1(new_n938_), .B2(new_n635_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n936_), .A2(new_n939_), .ZN(G1354gat));
  AOI21_X1  g739(.A(G218gat), .B1(new_n925_), .B2(new_n650_), .ZN(new_n941_));
  AND2_X1   g740(.A1(new_n925_), .A2(G218gat), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n941_), .B1(new_n702_), .B2(new_n942_), .ZN(G1355gat));
endmodule


