//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 0 0 0 0 0 1 1 0 0 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 0 1 1 1 1 0 1 1 1 0 1 0 1 0 1 0 1 0 0 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n875_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n917_, new_n919_, new_n920_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n932_;
  XOR2_X1   g000(.A(G1gat), .B(G8gat), .Z(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G15gat), .B(G22gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT76), .ZN(new_n205_));
  INV_X1    g004(.A(G1gat), .ZN(new_n206_));
  INV_X1    g005(.A(G8gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT14), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n204_), .A2(new_n205_), .A3(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n205_), .B1(new_n204_), .B2(new_n208_), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n203_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G29gat), .B(G36gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G43gat), .B(G50gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(G15gat), .B(G22gat), .Z(new_n216_));
  INV_X1    g015(.A(KEYINPUT14), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n217_), .B1(G1gat), .B2(G8gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT76), .B1(new_n216_), .B2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n219_), .A2(new_n202_), .A3(new_n209_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n212_), .A2(new_n215_), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G229gat), .A2(G233gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n215_), .B(KEYINPUT15), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NOR3_X1   g023(.A1(new_n210_), .A2(new_n203_), .A3(new_n211_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n202_), .B1(new_n219_), .B2(new_n209_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n221_), .B(new_n222_), .C1(new_n224_), .C2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n215_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n229_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(new_n221_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n222_), .ZN(new_n232_));
  AOI21_X1  g031(.A(KEYINPUT78), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT78), .ZN(new_n234_));
  AOI211_X1 g033(.A(new_n234_), .B(new_n222_), .C1(new_n230_), .C2(new_n221_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n228_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G113gat), .B(G141gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT79), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G169gat), .B(G197gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n236_), .A2(new_n241_), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n228_), .B(new_n240_), .C1(new_n233_), .C2(new_n235_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT80), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT96), .B(G106gat), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G22gat), .B(G50gat), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G155gat), .A2(G162gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT1), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT1), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n252_), .A2(G155gat), .A3(G162gat), .ZN(new_n253_));
  OR2_X1    g052(.A1(G155gat), .A2(G162gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n251_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(G141gat), .B(G148gat), .Z(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT89), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n255_), .A2(new_n256_), .A3(KEYINPUT89), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT29), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n254_), .A2(new_n250_), .ZN(new_n263_));
  AOI21_X1  g062(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT90), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(G141gat), .A2(G148gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT3), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n263_), .B1(new_n266_), .B2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n261_), .A2(new_n262_), .A3(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT28), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n264_), .B(KEYINPUT90), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n269_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  AOI22_X1  g077(.A1(new_n259_), .A2(new_n260_), .B1(new_n278_), .B2(new_n263_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT28), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n279_), .A2(new_n280_), .A3(new_n262_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G228gat), .A2(G233gat), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT95), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n275_), .A2(new_n281_), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n284_), .B1(new_n275_), .B2(new_n281_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n249_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n275_), .A2(new_n281_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n289_), .A2(new_n283_), .A3(new_n282_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n290_), .A2(new_n248_), .A3(new_n285_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G197gat), .B(G204gat), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n292_), .A2(KEYINPUT94), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT21), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n294_), .B1(new_n292_), .B2(KEYINPUT94), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G211gat), .B(G218gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT93), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G197gat), .B(G204gat), .Z(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT21), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT91), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT93), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n297_), .B(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(KEYINPUT92), .B(KEYINPUT21), .Z(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(new_n292_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n299_), .B1(new_n303_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n261_), .A2(new_n273_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT29), .ZN(new_n311_));
  NAND3_X1  g110(.A1(KEYINPUT95), .A2(G228gat), .A3(G233gat), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n309_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(G78gat), .ZN(new_n314_));
  INV_X1    g113(.A(G78gat), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n309_), .A2(new_n311_), .A3(new_n315_), .A4(new_n312_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  AND3_X1   g116(.A1(new_n288_), .A2(new_n291_), .A3(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n317_), .B1(new_n288_), .B2(new_n291_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n247_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n288_), .A2(new_n291_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n317_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n288_), .A2(new_n291_), .A3(new_n317_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(new_n246_), .A3(new_n324_), .ZN(new_n325_));
  AND2_X1   g124(.A1(new_n320_), .A2(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(G1gat), .B(G29gat), .Z(new_n327_));
  XNOR2_X1  g126(.A(G57gat), .B(G85gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT84), .ZN(new_n332_));
  XOR2_X1   g131(.A(G127gat), .B(G134gat), .Z(new_n333_));
  INV_X1    g132(.A(KEYINPUT83), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G127gat), .B(G134gat), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n336_), .A2(KEYINPUT83), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G113gat), .B(G120gat), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NOR3_X1   g138(.A1(new_n335_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n333_), .A2(new_n334_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n336_), .A2(KEYINPUT83), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n338_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n332_), .B1(new_n340_), .B2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n339_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n341_), .A2(new_n342_), .A3(new_n338_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(KEYINPUT84), .A3(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n279_), .B1(new_n344_), .B2(new_n347_), .ZN(new_n348_));
  NOR3_X1   g147(.A1(new_n310_), .A2(new_n340_), .A3(new_n343_), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT4), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n344_), .A2(new_n347_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(new_n310_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT4), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n350_), .A2(new_n354_), .A3(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n279_), .A2(new_n346_), .A3(new_n345_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n352_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n355_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n331_), .B1(new_n357_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n356_), .B1(new_n350_), .B2(new_n354_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n331_), .B1(new_n359_), .B2(new_n355_), .ZN(new_n364_));
  OAI21_X1  g163(.A(KEYINPUT33), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n362_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G226gat), .A2(G233gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT19), .ZN(new_n368_));
  INV_X1    g167(.A(new_n308_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n301_), .B(KEYINPUT91), .ZN(new_n370_));
  AOI22_X1  g169(.A1(new_n369_), .A2(new_n370_), .B1(new_n298_), .B2(new_n296_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT25), .B(G183gat), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT97), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n372_), .A2(new_n373_), .ZN(new_n375_));
  XOR2_X1   g174(.A(KEYINPUT26), .B(G190gat), .Z(new_n376_));
  OR3_X1    g175(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT24), .ZN(new_n378_));
  INV_X1    g177(.A(G169gat), .ZN(new_n379_));
  INV_X1    g178(.A(G176gat), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n378_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G183gat), .A2(G190gat), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT23), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n381_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n379_), .A2(new_n380_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G169gat), .A2(G176gat), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n387_), .A2(KEYINPUT24), .A3(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n386_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n388_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT22), .B(G169gat), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n392_), .B1(new_n393_), .B2(new_n380_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n384_), .A2(new_n385_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n395_), .B1(G183gat), .B2(G190gat), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n377_), .A2(new_n391_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT20), .B1(new_n371_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(G190gat), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n372_), .B1(KEYINPUT26), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(KEYINPUT81), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT81), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(G190gat), .ZN(new_n403_));
  AND3_X1   g202(.A1(new_n401_), .A2(new_n403_), .A3(KEYINPUT26), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n386_), .B(new_n389_), .C1(new_n400_), .C2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(G183gat), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n401_), .A2(new_n403_), .A3(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n395_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n394_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT82), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n405_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n410_), .B1(new_n405_), .B2(new_n409_), .ZN(new_n413_));
  NOR3_X1   g212(.A1(new_n309_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n368_), .B1(new_n398_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT20), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n416_), .B1(new_n371_), .B2(new_n397_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n368_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n309_), .B1(new_n413_), .B2(new_n412_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n417_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  XOR2_X1   g219(.A(G8gat), .B(G36gat), .Z(new_n421_));
  XNOR2_X1  g220(.A(G64gat), .B(G92gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n415_), .A2(new_n420_), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n426_), .B1(new_n415_), .B2(new_n420_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n361_), .A2(KEYINPUT100), .A3(KEYINPUT33), .ZN(new_n431_));
  AOI21_X1  g230(.A(KEYINPUT100), .B1(new_n361_), .B2(KEYINPUT33), .ZN(new_n432_));
  OAI211_X1 g231(.A(new_n366_), .B(new_n430_), .C1(new_n431_), .C2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n357_), .A2(new_n331_), .A3(new_n360_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n362_), .A2(new_n434_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n426_), .A2(KEYINPUT32), .ZN(new_n436_));
  NOR3_X1   g235(.A1(new_n398_), .A2(new_n414_), .A3(new_n368_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n418_), .B1(new_n417_), .B2(new_n419_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n436_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n415_), .A2(new_n420_), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n435_), .B(new_n439_), .C1(new_n440_), .C2(new_n436_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n326_), .A2(new_n433_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT31), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n351_), .B(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G71gat), .B(G99gat), .ZN(new_n445_));
  INV_X1    g244(.A(G43gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n447_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n405_), .A2(new_n409_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT82), .ZN(new_n450_));
  INV_X1    g249(.A(new_n447_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n450_), .A2(new_n411_), .A3(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G227gat), .A2(G233gat), .ZN(new_n453_));
  INV_X1    g252(.A(G15gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT30), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n448_), .A2(new_n452_), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n456_), .B1(new_n448_), .B2(new_n452_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n444_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT85), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  OAI211_X1 g261(.A(KEYINPUT85), .B(new_n444_), .C1(new_n458_), .C2(new_n459_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n448_), .A2(new_n452_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n456_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n351_), .B(KEYINPUT31), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n467_), .A2(new_n468_), .A3(new_n457_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT86), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n467_), .A2(new_n468_), .A3(KEYINPUT86), .A4(new_n457_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n464_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT87), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT87), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n464_), .A2(new_n473_), .A3(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n475_), .A2(KEYINPUT88), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT88), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n464_), .A2(new_n476_), .A3(new_n473_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n476_), .B1(new_n464_), .B2(new_n473_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n479_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n425_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n483_), .A2(KEYINPUT27), .A3(new_n427_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n484_), .B1(new_n430_), .B2(KEYINPUT27), .ZN(new_n485_));
  NOR3_X1   g284(.A1(new_n318_), .A2(new_n319_), .A3(new_n247_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n246_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n487_));
  OAI22_X1  g286(.A1(new_n485_), .A2(new_n435_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n442_), .A2(new_n478_), .A3(new_n482_), .A4(new_n488_), .ZN(new_n489_));
  NOR3_X1   g288(.A1(new_n485_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n435_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n475_), .A2(new_n477_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n245_), .B1(new_n489_), .B2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G120gat), .B(G148gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT5), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G176gat), .B(G204gat), .ZN(new_n497_));
  XOR2_X1   g296(.A(new_n496_), .B(new_n497_), .Z(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G57gat), .B(G64gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT11), .ZN(new_n501_));
  XOR2_X1   g300(.A(G71gat), .B(G78gat), .Z(new_n502_));
  OR2_X1    g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n500_), .A2(KEYINPUT11), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n501_), .A2(new_n502_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n503_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(G85gat), .A2(G92gat), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT65), .B1(G85gat), .B2(G92gat), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT9), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n507_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n510_), .B1(new_n509_), .B2(new_n508_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G99gat), .A2(G106gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT6), .ZN(new_n513_));
  OR2_X1    g312(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n514_), .A2(KEYINPUT64), .A3(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT64), .B1(new_n514_), .B2(new_n515_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n511_), .B(new_n513_), .C1(new_n518_), .C2(G106gat), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT8), .ZN(new_n520_));
  INV_X1    g319(.A(new_n512_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT67), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n522_), .A2(KEYINPUT6), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT6), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n524_), .A2(KEYINPUT67), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n521_), .B1(new_n523_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT66), .ZN(new_n527_));
  INV_X1    g326(.A(G99gat), .ZN(new_n528_));
  INV_X1    g327(.A(G106gat), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n527_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(KEYINPUT7), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT7), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n527_), .A2(new_n532_), .A3(new_n528_), .A4(new_n529_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n524_), .A2(KEYINPUT67), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n522_), .A2(KEYINPUT6), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n535_), .A3(new_n512_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n526_), .A2(new_n531_), .A3(new_n533_), .A4(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(G85gat), .B(G92gat), .Z(new_n538_));
  AOI21_X1  g337(.A(new_n520_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n520_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n531_), .A2(new_n533_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n540_), .B1(new_n541_), .B2(new_n513_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n506_), .B(new_n519_), .C1(new_n539_), .C2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G230gat), .A2(G233gat), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n519_), .B1(new_n539_), .B2(new_n542_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT12), .ZN(new_n547_));
  INV_X1    g346(.A(new_n506_), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n546_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n547_), .B1(new_n546_), .B2(new_n548_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n545_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n546_), .A2(new_n548_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(new_n543_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n544_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n551_), .A2(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n499_), .B1(new_n556_), .B2(KEYINPUT68), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n557_), .B1(KEYINPUT68), .B2(new_n556_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT69), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n559_), .B1(new_n556_), .B2(new_n498_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n551_), .A2(KEYINPUT69), .A3(new_n555_), .A4(new_n499_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n558_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n566_), .B1(new_n564_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n506_), .B(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(new_n227_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT77), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G127gat), .B(G155gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT16), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G183gat), .B(G211gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT17), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n573_), .B(new_n578_), .ZN(new_n579_));
  OR3_X1    g378(.A1(new_n571_), .A2(KEYINPUT17), .A3(new_n577_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G190gat), .B(G218gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G134gat), .B(G162gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT74), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT35), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G232gat), .A2(G233gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT34), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  AOI22_X1  g390(.A1(new_n546_), .A2(new_n223_), .B1(new_n588_), .B2(new_n591_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n215_), .B(new_n519_), .C1(new_n539_), .C2(new_n542_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT71), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n593_), .A2(new_n594_), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n587_), .B(new_n592_), .C1(new_n595_), .C2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(KEYINPUT72), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n593_), .B(new_n594_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT72), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n599_), .A2(new_n600_), .A3(new_n592_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n591_), .A2(new_n588_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n598_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n602_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n599_), .A2(new_n592_), .ZN(new_n605_));
  OAI211_X1 g404(.A(KEYINPUT72), .B(new_n604_), .C1(new_n605_), .C2(KEYINPUT74), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n586_), .B1(new_n603_), .B2(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(KEYINPUT73), .B1(new_n603_), .B2(new_n606_), .ZN(new_n608_));
  OAI22_X1  g407(.A1(KEYINPUT36), .A2(new_n607_), .B1(new_n608_), .B2(new_n585_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n603_), .A2(new_n606_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT73), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT36), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n612_), .A2(new_n613_), .A3(new_n586_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n609_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(KEYINPUT75), .B(KEYINPUT37), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n609_), .A2(new_n614_), .A3(new_n616_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n582_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n494_), .A2(new_n568_), .A3(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(new_n206_), .A3(new_n435_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT103), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n623_), .A2(KEYINPUT38), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n623_), .A2(KEYINPUT38), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n622_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT101), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n489_), .A2(new_n493_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n615_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n627_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  AOI211_X1 g429(.A(KEYINPUT101), .B(new_n615_), .C1(new_n489_), .C2(new_n493_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n568_), .A2(new_n581_), .A3(new_n244_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(KEYINPUT102), .B1(new_n632_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n632_), .A2(KEYINPUT102), .A3(new_n634_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n491_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  OAI221_X1 g437(.A(new_n626_), .B1(new_n624_), .B2(new_n622_), .C1(new_n638_), .C2(new_n206_), .ZN(G1324gat));
  NAND3_X1  g438(.A1(new_n621_), .A2(new_n207_), .A3(new_n485_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n485_), .B(new_n634_), .C1(new_n630_), .C2(new_n631_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT104), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n641_), .A2(new_n642_), .A3(G8gat), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n642_), .B1(new_n641_), .B2(G8gat), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n644_), .A2(new_n645_), .A3(KEYINPUT39), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT39), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n641_), .A2(G8gat), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT104), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n647_), .B1(new_n649_), .B2(new_n643_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n640_), .B1(new_n646_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT40), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  OAI211_X1 g452(.A(KEYINPUT40), .B(new_n640_), .C1(new_n646_), .C2(new_n650_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1325gat));
  NAND2_X1  g454(.A1(new_n482_), .A2(new_n478_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n621_), .A2(new_n454_), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n637_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n656_), .B1(new_n658_), .B2(new_n635_), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n659_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(KEYINPUT41), .B1(new_n659_), .B2(G15gat), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n657_), .B1(new_n660_), .B2(new_n661_), .ZN(G1326gat));
  INV_X1    g461(.A(G22gat), .ZN(new_n663_));
  INV_X1    g462(.A(new_n326_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n621_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n664_), .B1(new_n658_), .B2(new_n635_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT42), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n666_), .A2(new_n667_), .A3(G22gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n667_), .B1(new_n666_), .B2(G22gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n665_), .B1(new_n668_), .B2(new_n669_), .ZN(G1327gat));
  INV_X1    g469(.A(new_n568_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n615_), .A2(new_n582_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n494_), .A2(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(G29gat), .B1(new_n674_), .B2(new_n435_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n619_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n616_), .B1(new_n609_), .B2(new_n614_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n628_), .A2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT43), .ZN(new_n680_));
  INV_X1    g479(.A(new_n244_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n671_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(new_n582_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n680_), .A2(KEYINPUT44), .A3(new_n684_), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n685_), .A2(G29gat), .A3(new_n435_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n679_), .B(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n687_), .B1(new_n689_), .B2(new_n683_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n675_), .B1(new_n686_), .B2(new_n690_), .ZN(G1328gat));
  NAND3_X1  g490(.A1(new_n690_), .A2(new_n485_), .A3(new_n685_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(G36gat), .ZN(new_n693_));
  INV_X1    g492(.A(G36gat), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n485_), .A2(KEYINPUT105), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n485_), .A2(KEYINPUT105), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n674_), .A2(new_n694_), .A3(new_n697_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT45), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n693_), .A2(new_n699_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n693_), .B(new_n699_), .C1(KEYINPUT106), .C2(KEYINPUT46), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1329gat));
  NAND4_X1  g503(.A1(new_n690_), .A2(new_n685_), .A3(G43gat), .A4(new_n492_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n674_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n656_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n446_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n705_), .A2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n709_), .B(new_n710_), .ZN(G1330gat));
  AOI21_X1  g510(.A(G50gat), .B1(new_n674_), .B2(new_n664_), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n685_), .A2(G50gat), .A3(new_n664_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(new_n690_), .ZN(G1331gat));
  AND4_X1   g513(.A1(new_n632_), .A2(new_n581_), .A3(new_n671_), .A4(new_n245_), .ZN(new_n715_));
  INV_X1    g514(.A(G57gat), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n491_), .A2(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n244_), .B1(new_n489_), .B2(new_n493_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n718_), .A2(new_n671_), .A3(new_n620_), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n719_), .A2(KEYINPUT108), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(KEYINPUT108), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n720_), .A2(new_n435_), .A3(new_n721_), .ZN(new_n722_));
  AOI22_X1  g521(.A1(new_n715_), .A2(new_n717_), .B1(new_n722_), .B2(new_n716_), .ZN(G1332gat));
  INV_X1    g522(.A(new_n697_), .ZN(new_n724_));
  OR3_X1    g523(.A1(new_n719_), .A2(G64gat), .A3(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n715_), .A2(new_n697_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(G64gat), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n727_), .A2(KEYINPUT48), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n727_), .A2(KEYINPUT48), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(G1333gat));
  OR3_X1    g529(.A1(new_n719_), .A2(G71gat), .A3(new_n707_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n715_), .A2(new_n656_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(G71gat), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n733_), .A2(KEYINPUT49), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n733_), .A2(KEYINPUT49), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n731_), .B1(new_n734_), .B2(new_n735_), .ZN(G1334gat));
  NAND2_X1  g535(.A1(new_n715_), .A2(new_n664_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(G78gat), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n738_), .A2(KEYINPUT50), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(KEYINPUT50), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n664_), .A2(new_n315_), .ZN(new_n741_));
  OAI22_X1  g540(.A1(new_n739_), .A2(new_n740_), .B1(new_n719_), .B2(new_n741_), .ZN(G1335gat));
  NAND4_X1  g541(.A1(new_n718_), .A2(new_n615_), .A3(new_n582_), .A4(new_n671_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(G85gat), .B1(new_n744_), .B2(new_n435_), .ZN(new_n745_));
  NOR3_X1   g544(.A1(new_n568_), .A2(new_n581_), .A3(new_n244_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n680_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n435_), .A2(G85gat), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT109), .Z(new_n749_));
  AOI21_X1  g548(.A(new_n745_), .B1(new_n747_), .B2(new_n749_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT110), .Z(G1336gat));
  AOI21_X1  g550(.A(G92gat), .B1(new_n744_), .B2(new_n485_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n697_), .A2(G92gat), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT111), .Z(new_n754_));
  AOI21_X1  g553(.A(new_n752_), .B1(new_n747_), .B2(new_n754_), .ZN(G1337gat));
  AOI211_X1 g554(.A(new_n518_), .B(new_n743_), .C1(new_n475_), .C2(new_n477_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n747_), .A2(new_n656_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n757_), .B2(G99gat), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n758_), .B(new_n759_), .ZN(G1338gat));
  NAND3_X1  g559(.A1(new_n744_), .A2(new_n529_), .A3(new_n664_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n680_), .A2(new_n664_), .A3(new_n746_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n762_), .A2(new_n763_), .A3(G106gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n762_), .B2(G106gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n761_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n761_), .B(new_n767_), .C1(new_n764_), .C2(new_n765_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(G1339gat));
  OAI211_X1 g570(.A(new_n545_), .B(KEYINPUT55), .C1(new_n549_), .C2(new_n550_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n552_), .A2(KEYINPUT12), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n546_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n777_), .A2(KEYINPUT113), .A3(KEYINPUT55), .A4(new_n545_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT55), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n551_), .A2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n543_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n554_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n774_), .A2(new_n778_), .A3(new_n780_), .A4(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT56), .B1(new_n783_), .B2(new_n498_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n783_), .A2(KEYINPUT56), .A3(new_n498_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n562_), .A2(new_n244_), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n221_), .B(new_n232_), .C1(new_n224_), .C2(new_n227_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n240_), .B1(new_n231_), .B2(new_n222_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n243_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT114), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT114), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n243_), .A2(new_n791_), .A3(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  AOI22_X1  g595(.A1(new_n787_), .A2(new_n788_), .B1(new_n563_), .B2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT57), .ZN(new_n798_));
  OR3_X1    g597(.A1(new_n797_), .A2(new_n798_), .A3(new_n615_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT116), .ZN(new_n800_));
  AOI22_X1  g599(.A1(new_n793_), .A2(new_n795_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n783_), .A2(KEYINPUT56), .A3(new_n498_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n800_), .B(new_n801_), .C1(new_n802_), .C2(new_n784_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT58), .B1(new_n803_), .B2(KEYINPUT117), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT116), .B1(KEYINPUT117), .B2(KEYINPUT58), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n805_), .B1(new_n787_), .B2(new_n801_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n619_), .B(new_n618_), .C1(new_n804_), .C2(new_n806_), .ZN(new_n807_));
  XOR2_X1   g606(.A(KEYINPUT115), .B(KEYINPUT57), .Z(new_n808_));
  OAI21_X1  g607(.A(new_n808_), .B1(new_n797_), .B2(new_n615_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n799_), .A2(new_n807_), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n581_), .B1(new_n810_), .B2(KEYINPUT118), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n799_), .A2(new_n807_), .A3(new_n812_), .A4(new_n809_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n581_), .B(new_n568_), .C1(new_n676_), .C2(new_n677_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n245_), .ZN(new_n815_));
  OAI21_X1  g614(.A(KEYINPUT54), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n620_), .A2(new_n817_), .A3(new_n568_), .A4(new_n245_), .ZN(new_n818_));
  AOI22_X1  g617(.A1(new_n811_), .A2(new_n813_), .B1(new_n816_), .B2(new_n818_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n490_), .A2(new_n492_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n435_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT59), .B1(new_n819_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n807_), .A2(new_n809_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n807_), .A2(KEYINPUT119), .A3(new_n809_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(new_n799_), .A3(new_n826_), .ZN(new_n827_));
  AOI22_X1  g626(.A1(new_n827_), .A2(new_n582_), .B1(new_n816_), .B2(new_n818_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n821_), .A2(KEYINPUT59), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n822_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(G113gat), .B1(new_n831_), .B2(new_n245_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n819_), .A2(new_n821_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  OR2_X1    g633(.A1(new_n681_), .A2(G113gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n832_), .B1(new_n834_), .B2(new_n835_), .ZN(G1340gat));
  INV_X1    g635(.A(G120gat), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n816_), .A2(new_n818_), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n807_), .A2(KEYINPUT119), .A3(new_n809_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT119), .B1(new_n807_), .B2(new_n809_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n799_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n839_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n838_), .B1(new_n842_), .B2(new_n581_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n568_), .B1(new_n843_), .B2(new_n829_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n837_), .B1(new_n844_), .B2(new_n822_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n837_), .B1(new_n568_), .B2(KEYINPUT60), .ZN(new_n846_));
  OR2_X1    g645(.A1(new_n837_), .A2(KEYINPUT60), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n833_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(KEYINPUT120), .B1(new_n845_), .B2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n671_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT59), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n810_), .A2(KEYINPUT118), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n852_), .A2(new_n582_), .A3(new_n813_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n838_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n821_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n851_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(G120gat), .B1(new_n850_), .B2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n833_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n857_), .A2(new_n858_), .A3(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n849_), .A2(new_n860_), .ZN(G1341gat));
  OAI21_X1  g660(.A(G127gat), .B1(new_n831_), .B2(new_n582_), .ZN(new_n862_));
  OR2_X1    g661(.A1(new_n582_), .A2(G127gat), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n834_), .B2(new_n863_), .ZN(G1342gat));
  INV_X1    g663(.A(new_n678_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(KEYINPUT121), .B(G134gat), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n831_), .A2(new_n865_), .A3(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(G134gat), .B1(new_n833_), .B2(new_n615_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(G1343gat));
  NAND4_X1  g668(.A1(new_n724_), .A2(new_n707_), .A3(new_n435_), .A4(new_n664_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(KEYINPUT122), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n819_), .A2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n244_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g673(.A1(new_n872_), .A2(new_n671_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g675(.A1(new_n872_), .A2(new_n581_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(KEYINPUT61), .B(G155gat), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1346gat));
  AOI21_X1  g678(.A(G162gat), .B1(new_n872_), .B2(new_n615_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n678_), .A2(G162gat), .ZN(new_n881_));
  XOR2_X1   g680(.A(new_n881_), .B(KEYINPUT123), .Z(new_n882_));
  AOI21_X1  g681(.A(new_n880_), .B1(new_n872_), .B2(new_n882_), .ZN(G1347gat));
  INV_X1    g682(.A(KEYINPUT124), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n379_), .B1(new_n884_), .B2(KEYINPUT62), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n724_), .A2(new_n435_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n656_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n843_), .A2(new_n326_), .A3(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n885_), .B1(new_n889_), .B2(new_n681_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT62), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n890_), .A2(KEYINPUT124), .A3(new_n891_), .ZN(new_n892_));
  OAI221_X1 g691(.A(new_n885_), .B1(new_n884_), .B2(KEYINPUT62), .C1(new_n889_), .C2(new_n681_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n889_), .A2(new_n681_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n393_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n892_), .A2(new_n893_), .A3(new_n895_), .ZN(G1348gat));
  OR2_X1    g695(.A1(new_n889_), .A2(new_n568_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n819_), .A2(new_n664_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n887_), .A2(new_n380_), .A3(new_n568_), .ZN(new_n899_));
  AOI22_X1  g698(.A1(new_n897_), .A2(new_n380_), .B1(new_n898_), .B2(new_n899_), .ZN(G1349gat));
  OAI21_X1  g699(.A(new_n581_), .B1(new_n375_), .B2(new_n374_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n889_), .A2(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n887_), .A2(new_n582_), .ZN(new_n903_));
  AOI21_X1  g702(.A(G183gat), .B1(new_n898_), .B2(new_n903_), .ZN(new_n904_));
  OAI21_X1  g703(.A(KEYINPUT125), .B1(new_n902_), .B2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n854_), .A2(new_n326_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n903_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n406_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT125), .ZN(new_n909_));
  OAI211_X1 g708(.A(new_n908_), .B(new_n909_), .C1(new_n889_), .C2(new_n901_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n905_), .A2(new_n910_), .ZN(G1350gat));
  OAI21_X1  g710(.A(G190gat), .B1(new_n889_), .B2(new_n865_), .ZN(new_n912_));
  OR2_X1    g711(.A1(new_n629_), .A2(new_n376_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n889_), .B2(new_n913_), .ZN(G1351gat));
  NAND3_X1  g713(.A1(new_n886_), .A2(new_n707_), .A3(new_n664_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n819_), .A2(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n244_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g717(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n919_));
  XNOR2_X1  g718(.A(KEYINPUT126), .B(G204gat), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n916_), .A2(new_n671_), .ZN(new_n921_));
  MUX2_X1   g720(.A(new_n919_), .B(new_n920_), .S(new_n921_), .Z(G1353gat));
  INV_X1    g721(.A(KEYINPUT63), .ZN(new_n923_));
  INV_X1    g722(.A(G211gat), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n581_), .B1(new_n923_), .B2(new_n924_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(KEYINPUT127), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n916_), .A2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n923_), .A2(new_n924_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n927_), .B(new_n928_), .ZN(G1354gat));
  INV_X1    g728(.A(G218gat), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n916_), .A2(new_n930_), .A3(new_n615_), .ZN(new_n931_));
  NOR3_X1   g730(.A1(new_n819_), .A2(new_n865_), .A3(new_n915_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n932_), .B2(new_n930_), .ZN(G1355gat));
endmodule


