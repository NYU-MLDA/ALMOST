//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 1 1 0 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n809_, new_n810_, new_n811_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n824_, new_n825_, new_n826_, new_n827_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n853_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n945_, new_n946_, new_n947_,
    new_n949_, new_n951_, new_n952_, new_n954_, new_n955_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n979_, new_n980_, new_n982_, new_n983_, new_n985_,
    new_n986_, new_n987_, new_n989_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_,
    new_n1001_, new_n1002_, new_n1003_, new_n1004_;
  XNOR2_X1  g000(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G226gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT21), .ZN(new_n205_));
  INV_X1    g004(.A(G204gat), .ZN(new_n206_));
  INV_X1    g005(.A(G197gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT93), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT93), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G197gat), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n206_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G197gat), .A2(G204gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n205_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G218gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(G211gat), .ZN(new_n215_));
  INV_X1    g014(.A(G211gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(G218gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n208_), .A2(new_n210_), .A3(new_n206_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n205_), .B1(G197gat), .B2(G204gat), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n218_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n208_), .A2(new_n210_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n212_), .B1(new_n222_), .B2(G204gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n205_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n224_));
  AOI22_X1  g023(.A1(new_n213_), .A2(new_n221_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT23), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(G183gat), .A3(G190gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT83), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n226_), .A2(KEYINPUT83), .A3(G183gat), .A4(G190gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231_));
  AND3_X1   g030(.A1(new_n231_), .A2(KEYINPUT82), .A3(KEYINPUT23), .ZN(new_n232_));
  AOI21_X1  g031(.A(KEYINPUT82), .B1(new_n231_), .B2(KEYINPUT23), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n229_), .B(new_n230_), .C1(new_n232_), .C2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(G183gat), .ZN(new_n235_));
  INV_X1    g034(.A(G190gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n234_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT100), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT100), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n234_), .A2(new_n240_), .A3(new_n237_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT22), .B(G169gat), .ZN(new_n242_));
  INV_X1    g041(.A(G176gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G169gat), .A2(G176gat), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT81), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n244_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n239_), .A2(new_n241_), .A3(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(G169gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(new_n243_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n252_), .A2(KEYINPUT24), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n231_), .A2(KEYINPUT23), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n253_), .B1(new_n254_), .B2(new_n227_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n245_), .A2(KEYINPUT24), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n256_), .A2(KEYINPUT99), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n252_), .B1(new_n256_), .B2(KEYINPUT99), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT25), .B(G183gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT98), .ZN(new_n260_));
  XOR2_X1   g059(.A(KEYINPUT26), .B(G190gat), .Z(new_n261_));
  OAI221_X1 g060(.A(new_n255_), .B1(new_n257_), .B2(new_n258_), .C1(new_n260_), .C2(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n225_), .B1(new_n250_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n252_), .A2(KEYINPUT24), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n253_), .B1(new_n247_), .B2(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n236_), .A2(KEYINPUT26), .ZN(new_n267_));
  AOI22_X1  g066(.A1(new_n267_), .A2(KEYINPUT80), .B1(KEYINPUT25), .B2(new_n235_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT80), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n269_), .B1(new_n236_), .B2(KEYINPUT26), .ZN(new_n270_));
  OR2_X1    g069(.A1(KEYINPUT79), .A2(G190gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(KEYINPUT79), .A2(G190gat), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(KEYINPUT26), .A3(new_n272_), .ZN(new_n273_));
  OR2_X1    g072(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n274_));
  NAND2_X1  g073(.A1(KEYINPUT78), .A2(KEYINPUT25), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n274_), .A2(G183gat), .A3(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n268_), .A2(new_n270_), .A3(new_n273_), .A4(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n266_), .A2(new_n277_), .A3(new_n234_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT84), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n279_), .B1(new_n251_), .B2(KEYINPUT22), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n243_), .B(new_n280_), .C1(new_n242_), .C2(new_n279_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n271_), .A2(new_n235_), .A3(new_n272_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n254_), .A2(new_n227_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n281_), .A2(new_n247_), .A3(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n278_), .A2(new_n225_), .A3(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT20), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n204_), .B1(new_n263_), .B2(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(G8gat), .B(G36gat), .Z(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT18), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G64gat), .B(G92gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n250_), .A2(new_n262_), .A3(new_n225_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT20), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n278_), .A2(new_n285_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n213_), .A2(new_n221_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n223_), .A2(new_n224_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n294_), .B1(new_n295_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n204_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n293_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n288_), .A2(new_n292_), .A3(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT27), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n293_), .A2(new_n299_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n204_), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n234_), .A2(new_n240_), .A3(new_n237_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n240_), .B1(new_n234_), .B2(new_n237_), .ZN(new_n307_));
  NOR3_X1   g106(.A1(new_n306_), .A2(new_n307_), .A3(new_n248_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT98), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n259_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n259_), .A2(new_n309_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n261_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n255_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n257_), .A2(new_n258_), .ZN(new_n314_));
  NOR3_X1   g113(.A1(new_n312_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n298_), .B1(new_n308_), .B2(new_n315_), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n286_), .A2(KEYINPUT20), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n316_), .A2(new_n317_), .A3(new_n300_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n292_), .B1(new_n305_), .B2(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n303_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n292_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n300_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n293_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n321_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(KEYINPUT27), .B1(new_n324_), .B2(new_n302_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n320_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G78gat), .B(G106gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT94), .ZN(new_n329_));
  INV_X1    g128(.A(G228gat), .ZN(new_n330_));
  INV_X1    g129(.A(G233gat), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n225_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(G155gat), .ZN(new_n335_));
  INV_X1    g134(.A(G162gat), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(new_n336_), .A3(KEYINPUT88), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT88), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n338_), .B1(G155gat), .B2(G162gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G155gat), .A2(G162gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n337_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT3), .ZN(new_n343_));
  INV_X1    g142(.A(G141gat), .ZN(new_n344_));
  INV_X1    g143(.A(G148gat), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n343_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT89), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(G141gat), .A2(G148gat), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n349_), .A2(KEYINPUT89), .A3(new_n343_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G141gat), .A2(G148gat), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT90), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT2), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n352_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n356_));
  AOI21_X1  g155(.A(KEYINPUT90), .B1(G141gat), .B2(G148gat), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n355_), .B(new_n356_), .C1(new_n354_), .C2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n342_), .B1(new_n351_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n340_), .A2(KEYINPUT1), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT1), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n361_), .A2(G155gat), .A3(G162gat), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n360_), .A2(new_n337_), .A3(new_n339_), .A4(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n352_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n364_), .A2(new_n349_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n359_), .A2(KEYINPUT91), .A3(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(KEYINPUT91), .B1(new_n359_), .B2(new_n366_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n334_), .B1(new_n369_), .B2(KEYINPUT29), .ZN(new_n370_));
  INV_X1    g169(.A(new_n349_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(KEYINPUT90), .A2(KEYINPUT2), .ZN(new_n372_));
  AOI22_X1  g171(.A1(new_n371_), .A2(KEYINPUT3), .B1(new_n372_), .B2(new_n352_), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT2), .B1(new_n364_), .B2(KEYINPUT90), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n373_), .A2(new_n348_), .A3(new_n374_), .A4(new_n350_), .ZN(new_n375_));
  AOI22_X1  g174(.A1(new_n375_), .A2(new_n342_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT29), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n298_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n378_), .A2(new_n332_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n329_), .B1(new_n370_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT95), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT91), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n355_), .A2(new_n356_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n357_), .A2(new_n354_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NOR4_X1   g184(.A1(new_n347_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n386_));
  AOI21_X1  g185(.A(KEYINPUT89), .B1(new_n349_), .B2(new_n343_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n341_), .B1(new_n385_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n366_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n382_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n359_), .A2(KEYINPUT91), .A3(new_n366_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(KEYINPUT29), .A3(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(new_n333_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n329_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n378_), .A2(new_n332_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n380_), .A2(new_n381_), .A3(new_n397_), .ZN(new_n398_));
  OAI211_X1 g197(.A(KEYINPUT95), .B(new_n329_), .C1(new_n370_), .C2(new_n379_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G22gat), .B(G50gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT28), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n401_), .B1(new_n369_), .B2(KEYINPUT29), .ZN(new_n402_));
  INV_X1    g201(.A(new_n401_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n377_), .B(new_n403_), .C1(new_n367_), .C2(new_n368_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT92), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n402_), .A2(KEYINPUT92), .A3(new_n404_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n398_), .A2(new_n399_), .A3(new_n407_), .A4(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT96), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n395_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n410_), .B1(new_n413_), .B2(new_n405_), .ZN(new_n414_));
  AND4_X1   g213(.A1(new_n410_), .A2(new_n380_), .A3(new_n405_), .A4(new_n397_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n409_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G113gat), .B(G120gat), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G127gat), .B(G134gat), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT87), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n419_), .A2(new_n420_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n418_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n423_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(new_n421_), .A3(new_n417_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n391_), .A2(new_n392_), .A3(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n376_), .A2(new_n426_), .A3(new_n424_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G225gat), .A2(G233gat), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n428_), .A2(KEYINPUT4), .A3(new_n429_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT4), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n391_), .A2(new_n433_), .A3(new_n392_), .A4(new_n427_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n430_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n431_), .B1(new_n432_), .B2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G1gat), .B(G29gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(G85gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT0), .B(G57gat), .ZN(new_n440_));
  XOR2_X1   g239(.A(new_n439_), .B(new_n440_), .Z(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n437_), .A2(new_n442_), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n431_), .B(new_n441_), .C1(new_n432_), .C2(new_n436_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G227gat), .A2(G233gat), .ZN(new_n447_));
  XOR2_X1   g246(.A(new_n447_), .B(G71gat), .Z(new_n448_));
  INV_X1    g247(.A(G99gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(KEYINPUT85), .B(KEYINPUT30), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n448_), .B(G99gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n451_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(new_n427_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G15gat), .B(G43gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT86), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n295_), .A2(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n295_), .A2(new_n459_), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT31), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  OR3_X1    g261(.A1(new_n460_), .A2(new_n461_), .A3(KEYINPUT31), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n457_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n457_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n446_), .A2(new_n466_), .ZN(new_n467_));
  NOR3_X1   g266(.A1(new_n327_), .A2(new_n416_), .A3(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n416_), .A2(new_n326_), .A3(new_n446_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n324_), .A2(new_n302_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT33), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n444_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n428_), .A2(new_n429_), .A3(KEYINPUT4), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n474_), .A2(new_n435_), .A3(new_n434_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n442_), .A2(new_n472_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n475_), .A2(new_n431_), .A3(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n428_), .A2(new_n429_), .A3(new_n435_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n434_), .A2(new_n430_), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n442_), .B(new_n478_), .C1(new_n432_), .C2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n473_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n305_), .A2(new_n318_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n292_), .A2(KEYINPUT32), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT101), .B1(new_n483_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT101), .ZN(new_n487_));
  AOI211_X1 g286(.A(new_n487_), .B(new_n484_), .C1(new_n305_), .C2(new_n318_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n288_), .A2(new_n301_), .A3(new_n484_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n491_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n492_));
  AOI22_X1  g291(.A1(new_n471_), .A2(new_n482_), .B1(new_n489_), .B2(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n469_), .B1(new_n493_), .B2(new_n416_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n466_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n468_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G113gat), .B(G141gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G169gat), .B(G197gat), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n497_), .B(new_n498_), .Z(new_n499_));
  XNOR2_X1  g298(.A(G29gat), .B(G36gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT69), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G43gat), .B(G50gat), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n500_), .A2(KEYINPUT69), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n500_), .A2(KEYINPUT69), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(new_n506_), .A3(new_n502_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n504_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G15gat), .B(G22gat), .ZN(new_n509_));
  INV_X1    g308(.A(G1gat), .ZN(new_n510_));
  INV_X1    g309(.A(G8gat), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT14), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n509_), .A2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G1gat), .B(G8gat), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n513_), .B(new_n514_), .Z(new_n515_));
  NAND2_X1  g314(.A1(new_n508_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G229gat), .A2(G233gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n504_), .A2(KEYINPUT15), .A3(new_n507_), .ZN(new_n519_));
  AOI21_X1  g318(.A(KEYINPUT15), .B1(new_n504_), .B2(new_n507_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n515_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n521_), .A2(KEYINPUT77), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT15), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n508_), .A2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n504_), .A2(KEYINPUT15), .A3(new_n507_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n525_), .A2(new_n522_), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT77), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n518_), .B1(new_n523_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n522_), .A2(new_n504_), .A3(new_n507_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n516_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT76), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n517_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n532_), .A2(KEYINPUT76), .A3(new_n516_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n499_), .B1(new_n531_), .B2(new_n538_), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n499_), .ZN(new_n541_));
  NOR3_X1   g340(.A1(new_n540_), .A2(new_n530_), .A3(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n539_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n496_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT102), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n544_), .A2(KEYINPUT102), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT37), .ZN(new_n549_));
  AND2_X1   g348(.A1(G85gat), .A2(G92gat), .ZN(new_n550_));
  NOR2_X1   g349(.A1(G85gat), .A2(G92gat), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(G99gat), .A2(G106gat), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT7), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G99gat), .A2(G106gat), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT6), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n552_), .B1(new_n555_), .B2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT8), .ZN(new_n560_));
  XOR2_X1   g359(.A(KEYINPUT10), .B(G99gat), .Z(new_n561_));
  INV_X1    g360(.A(G106gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n552_), .A2(KEYINPUT9), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n556_), .B(KEYINPUT6), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT9), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n550_), .A2(new_n566_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n563_), .A2(new_n564_), .A3(new_n565_), .A4(new_n567_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n560_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT35), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G232gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT34), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  AOI22_X1  g372(.A1(new_n569_), .A2(new_n508_), .B1(new_n570_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT66), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n568_), .A2(new_n575_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n565_), .A2(new_n567_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n577_), .A2(KEYINPUT66), .A3(new_n563_), .A4(new_n564_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n559_), .A2(KEYINPUT8), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n559_), .A2(KEYINPUT8), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n576_), .B(new_n578_), .C1(new_n579_), .C2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n581_), .A2(new_n526_), .A3(new_n525_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n582_), .A2(KEYINPUT70), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT70), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n584_), .B1(new_n521_), .B2(new_n581_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n574_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n573_), .A2(new_n570_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n582_), .A2(KEYINPUT70), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n521_), .A2(new_n584_), .A3(new_n581_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n587_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n591_), .A2(new_n592_), .A3(new_n574_), .ZN(new_n593_));
  XOR2_X1   g392(.A(G190gat), .B(G218gat), .Z(new_n594_));
  XNOR2_X1  g393(.A(G134gat), .B(G162gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT36), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT71), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n588_), .A2(new_n593_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT72), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n549_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n596_), .B(KEYINPUT36), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n591_), .A2(new_n592_), .A3(new_n574_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n592_), .B1(new_n591_), .B2(new_n574_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n603_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(new_n600_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n602_), .A2(new_n607_), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n606_), .B(new_n600_), .C1(new_n601_), .C2(new_n549_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G57gat), .B(G64gat), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT64), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(KEYINPUT11), .ZN(new_n614_));
  XOR2_X1   g413(.A(G71gat), .B(G78gat), .Z(new_n615_));
  OR2_X1    g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G231gat), .A2(G233gat), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n611_), .B(KEYINPUT64), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT11), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n614_), .A2(new_n621_), .A3(new_n615_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n616_), .A2(new_n618_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n618_), .B1(new_n616_), .B2(new_n622_), .ZN(new_n625_));
  OAI21_X1  g424(.A(KEYINPUT73), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n616_), .A2(new_n622_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n617_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT73), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(new_n629_), .A3(new_n623_), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n626_), .A2(new_n630_), .A3(new_n515_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n515_), .B1(new_n626_), .B2(new_n630_), .ZN(new_n632_));
  OAI21_X1  g431(.A(KEYINPUT74), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n626_), .A2(new_n630_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(new_n522_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT74), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n626_), .A2(new_n630_), .A3(new_n515_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n635_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  XOR2_X1   g437(.A(G127gat), .B(G155gat), .Z(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT16), .ZN(new_n640_));
  XNOR2_X1  g439(.A(G183gat), .B(G211gat), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT17), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n633_), .A2(new_n638_), .A3(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n642_), .B(KEYINPUT17), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n646_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT75), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  OAI211_X1 g448(.A(KEYINPUT75), .B(new_n646_), .C1(new_n631_), .C2(new_n632_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n645_), .A2(new_n649_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT65), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n614_), .A2(new_n615_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n614_), .A2(new_n615_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n653_), .B1(new_n654_), .B2(new_n621_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n560_), .A2(new_n568_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n652_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n569_), .A2(KEYINPUT65), .A3(new_n627_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n655_), .A2(new_n656_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n657_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(G230gat), .A2(G233gat), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT12), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n664_), .B1(new_n569_), .B2(new_n627_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n662_), .B1(new_n569_), .B2(new_n627_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n655_), .A2(KEYINPUT12), .A3(new_n581_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n665_), .A2(new_n666_), .A3(new_n667_), .ZN(new_n668_));
  XOR2_X1   g467(.A(G120gat), .B(G148gat), .Z(new_n669_));
  XNOR2_X1  g468(.A(G176gat), .B(G204gat), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n671_), .B(new_n672_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n663_), .A2(new_n668_), .A3(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n663_), .B2(new_n668_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(KEYINPUT68), .A2(KEYINPUT13), .ZN(new_n676_));
  NAND2_X1  g475(.A1(KEYINPUT68), .A2(KEYINPUT13), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  OAI22_X1  g477(.A1(new_n674_), .A2(new_n675_), .B1(new_n676_), .B2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n663_), .A2(new_n668_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n673_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n663_), .A2(new_n668_), .A3(new_n673_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(new_n683_), .A3(new_n677_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n679_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n610_), .A2(new_n651_), .A3(new_n686_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n548_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n446_), .A2(G1gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n688_), .A2(new_n689_), .A3(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n548_), .A2(new_n687_), .A3(new_n690_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(KEYINPUT103), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(new_n694_));
  XOR2_X1   g493(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n695_));
  OAI21_X1  g494(.A(KEYINPUT105), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n697_));
  INV_X1    g496(.A(new_n695_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n691_), .A2(new_n697_), .A3(new_n693_), .A4(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n696_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n651_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n543_), .B1(new_n679_), .B2(new_n684_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT106), .ZN(new_n704_));
  INV_X1    g503(.A(new_n607_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n496_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n510_), .B1(new_n708_), .B2(new_n445_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n700_), .A2(new_n710_), .ZN(G1324gat));
  NAND3_X1  g510(.A1(new_n688_), .A2(new_n511_), .A3(new_n327_), .ZN(new_n712_));
  OAI21_X1  g511(.A(G8gat), .B1(new_n707_), .B2(new_n326_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT39), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n715_), .B(new_n716_), .Z(G1325gat));
  OAI21_X1  g516(.A(G15gat), .B1(new_n707_), .B2(new_n495_), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT41), .Z(new_n719_));
  INV_X1    g518(.A(G15gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n688_), .A2(new_n720_), .A3(new_n466_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(G1326gat));
  INV_X1    g521(.A(G22gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n688_), .A2(new_n723_), .A3(new_n416_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n380_), .A2(new_n405_), .A3(new_n397_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT96), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n413_), .A2(new_n410_), .A3(new_n405_), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n407_), .A2(new_n399_), .A3(new_n408_), .ZN(new_n728_));
  AOI22_X1  g527(.A1(new_n726_), .A2(new_n727_), .B1(new_n728_), .B2(new_n398_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G22gat), .B1(new_n707_), .B2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT42), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n724_), .A2(new_n731_), .ZN(G1327gat));
  NAND2_X1  g531(.A1(new_n651_), .A2(new_n705_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n733_), .A2(new_n686_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n548_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(G29gat), .B1(new_n736_), .B2(new_n445_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT108), .ZN(new_n738_));
  INV_X1    g537(.A(new_n543_), .ZN(new_n739_));
  AND4_X1   g538(.A1(new_n738_), .A2(new_n685_), .A3(new_n739_), .A4(new_n651_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n738_), .B1(new_n702_), .B2(new_n651_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n608_), .A2(new_n609_), .ZN(new_n743_));
  OAI21_X1  g542(.A(KEYINPUT43), .B1(new_n496_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT43), .ZN(new_n745_));
  INV_X1    g544(.A(new_n444_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n441_), .B1(new_n475_), .B2(new_n431_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n490_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n263_), .A2(new_n287_), .A3(new_n204_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n300_), .B1(new_n293_), .B2(new_n299_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n485_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(new_n487_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n483_), .A2(KEYINPUT101), .A3(new_n485_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n748_), .A2(new_n754_), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n473_), .A2(new_n470_), .A3(new_n481_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n729_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n466_), .B1(new_n757_), .B2(new_n469_), .ZN(new_n758_));
  OAI211_X1 g557(.A(new_n610_), .B(new_n745_), .C1(new_n758_), .C2(new_n468_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n742_), .B1(new_n744_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT109), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n740_), .A2(new_n741_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n468_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n477_), .B(new_n480_), .C1(new_n746_), .C2(KEYINPUT33), .ZN(new_n765_));
  OAI22_X1  g564(.A1(new_n765_), .A2(new_n470_), .B1(new_n748_), .B2(new_n754_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n727_), .A2(new_n726_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n445_), .B1(new_n767_), .B2(new_n409_), .ZN(new_n768_));
  AOI22_X1  g567(.A1(new_n766_), .A2(new_n729_), .B1(new_n768_), .B2(new_n326_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n764_), .B1(new_n769_), .B2(new_n466_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n745_), .B1(new_n770_), .B2(new_n610_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n759_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n763_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT44), .B1(new_n773_), .B2(KEYINPUT109), .ZN(new_n774_));
  OAI211_X1 g573(.A(KEYINPUT44), .B(new_n763_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT110), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT110), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n760_), .A2(new_n777_), .A3(KEYINPUT44), .ZN(new_n778_));
  AOI22_X1  g577(.A1(new_n762_), .A2(new_n774_), .B1(new_n776_), .B2(new_n778_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n445_), .A2(G29gat), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n737_), .B1(new_n779_), .B2(new_n780_), .ZN(G1328gat));
  INV_X1    g580(.A(KEYINPUT112), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT46), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n782_), .A2(KEYINPUT46), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n326_), .A2(G36gat), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n734_), .B(new_n785_), .C1(new_n546_), .C2(new_n547_), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n786_), .A2(KEYINPUT45), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(KEYINPUT45), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n784_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n776_), .A2(new_n778_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n773_), .A2(KEYINPUT109), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT44), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n792_), .A3(new_n762_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n790_), .A2(new_n793_), .A3(KEYINPUT111), .A4(new_n327_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(G36gat), .ZN(new_n795_));
  AOI21_X1  g594(.A(KEYINPUT111), .B1(new_n779_), .B2(new_n327_), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n783_), .B(new_n789_), .C1(new_n795_), .C2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT111), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n775_), .A2(KEYINPUT110), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n777_), .B1(new_n760_), .B2(KEYINPUT44), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n792_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n802_));
  AOI211_X1 g601(.A(KEYINPUT109), .B(new_n742_), .C1(new_n744_), .C2(new_n759_), .ZN(new_n803_));
  OAI22_X1  g602(.A1(new_n800_), .A2(new_n801_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n799_), .B1(new_n804_), .B2(new_n326_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(G36gat), .A3(new_n794_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n783_), .B1(new_n806_), .B2(new_n789_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n798_), .A2(new_n807_), .ZN(G1329gat));
  NAND3_X1  g607(.A1(new_n779_), .A2(G43gat), .A3(new_n466_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n735_), .A2(new_n495_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(G43gat), .B2(new_n810_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g611(.A1(new_n735_), .A2(G50gat), .A3(new_n729_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n779_), .A2(KEYINPUT113), .A3(new_n416_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(G50gat), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT113), .B1(new_n779_), .B2(new_n416_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n813_), .B1(new_n815_), .B2(new_n816_), .ZN(G1331gat));
  NAND4_X1  g616(.A1(new_n706_), .A2(new_n543_), .A3(new_n701_), .A4(new_n686_), .ZN(new_n818_));
  OAI21_X1  g617(.A(G57gat), .B1(new_n818_), .B2(new_n446_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n496_), .A2(new_n739_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n820_), .A2(new_n743_), .A3(new_n701_), .A4(new_n686_), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n446_), .A2(G57gat), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n819_), .B1(new_n821_), .B2(new_n822_), .ZN(G1332gat));
  OAI21_X1  g622(.A(G64gat), .B1(new_n818_), .B2(new_n326_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(KEYINPUT48), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n326_), .A2(G64gat), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(KEYINPUT114), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n825_), .B1(new_n821_), .B2(new_n827_), .ZN(G1333gat));
  OAI21_X1  g627(.A(G71gat), .B1(new_n818_), .B2(new_n495_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n829_), .B(KEYINPUT49), .ZN(new_n830_));
  OR2_X1    g629(.A1(new_n495_), .A2(G71gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n821_), .B2(new_n831_), .ZN(G1334gat));
  OAI21_X1  g631(.A(G78gat), .B1(new_n818_), .B2(new_n729_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(KEYINPUT50), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n729_), .A2(G78gat), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(KEYINPUT115), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n834_), .B1(new_n821_), .B2(new_n836_), .ZN(G1335gat));
  NOR2_X1   g636(.A1(new_n733_), .A2(new_n685_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n820_), .A2(new_n838_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n839_), .A2(G85gat), .A3(new_n446_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n686_), .A2(new_n543_), .A3(new_n651_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n841_), .B1(new_n744_), .B2(new_n759_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n445_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n840_), .B1(G85gat), .B2(new_n843_), .ZN(new_n844_));
  XOR2_X1   g643(.A(new_n844_), .B(KEYINPUT116), .Z(G1336gat));
  INV_X1    g644(.A(new_n839_), .ZN(new_n846_));
  INV_X1    g645(.A(G92gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(new_n847_), .A3(new_n327_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n842_), .A2(new_n327_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(new_n847_), .ZN(G1337gat));
  AOI21_X1  g649(.A(new_n449_), .B1(new_n842_), .B2(new_n466_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n466_), .A2(new_n561_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n851_), .B1(new_n846_), .B2(new_n852_), .ZN(new_n853_));
  XOR2_X1   g652(.A(new_n853_), .B(KEYINPUT51), .Z(G1338gat));
  AOI21_X1  g653(.A(new_n562_), .B1(new_n842_), .B2(new_n416_), .ZN(new_n855_));
  XOR2_X1   g654(.A(new_n855_), .B(KEYINPUT52), .Z(new_n856_));
  NAND3_X1  g655(.A1(new_n846_), .A2(new_n562_), .A3(new_n416_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g658(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n705_), .A2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n674_), .A2(new_n675_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n540_), .A2(new_n530_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n499_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n535_), .A2(new_n517_), .A3(new_n537_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n866_), .A2(new_n541_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n523_), .A2(new_n529_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n868_), .A2(new_n536_), .A3(new_n516_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n867_), .A2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n865_), .A2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n862_), .B1(new_n863_), .B2(new_n871_), .ZN(new_n872_));
  AOI22_X1  g671(.A1(new_n864_), .A2(new_n499_), .B1(new_n867_), .B2(new_n869_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n873_), .B(KEYINPUT118), .C1(new_n675_), .C2(new_n674_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n872_), .A2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n683_), .B1(new_n539_), .B2(new_n542_), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n665_), .A2(new_n657_), .A3(new_n658_), .A4(new_n667_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n662_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT55), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n668_), .A2(new_n879_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n665_), .A2(new_n666_), .A3(KEYINPUT55), .A4(new_n667_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n878_), .A2(new_n880_), .A3(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n681_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT56), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n882_), .A2(KEYINPUT56), .A3(new_n681_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n876_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n861_), .B1(new_n875_), .B2(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n888_), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n889_));
  NAND2_X1  g688(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n890_), .B(new_n861_), .C1(new_n875_), .C2(new_n887_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n885_), .A2(new_n886_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n871_), .A2(new_n674_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n892_), .A2(KEYINPUT58), .A3(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n893_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT58), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n743_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n897_));
  AOI22_X1  g696(.A1(new_n889_), .A2(new_n891_), .B1(new_n894_), .B2(new_n897_), .ZN(new_n898_));
  OAI21_X1  g697(.A(KEYINPUT122), .B1(new_n898_), .B2(new_n701_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n687_), .A2(new_n543_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n900_), .B(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n895_), .A2(new_n896_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n903_), .A2(new_n610_), .A3(new_n894_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n876_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n892_), .A2(new_n905_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n906_), .A2(new_n872_), .A3(new_n874_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n890_), .B1(new_n907_), .B2(new_n861_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n891_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n904_), .B1(new_n908_), .B2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n910_), .A2(new_n911_), .A3(new_n651_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n899_), .A2(new_n902_), .A3(new_n912_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n327_), .A2(new_n416_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n914_), .A2(new_n445_), .A3(new_n466_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  XOR2_X1   g715(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n917_));
  NAND3_X1  g716(.A1(new_n913_), .A2(new_n916_), .A3(new_n917_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n904_), .B(KEYINPUT119), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n889_), .A2(new_n891_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n701_), .B1(new_n919_), .B2(new_n920_), .ZN(new_n921_));
  XOR2_X1   g720(.A(new_n900_), .B(new_n901_), .Z(new_n922_));
  NOR2_X1   g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n923_), .A2(new_n915_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT59), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n918_), .B1(new_n924_), .B2(new_n925_), .ZN(new_n926_));
  OAI21_X1  g725(.A(G113gat), .B1(new_n926_), .B2(new_n543_), .ZN(new_n927_));
  OR2_X1    g726(.A1(new_n921_), .A2(new_n922_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(new_n916_), .ZN(new_n929_));
  OR2_X1    g728(.A1(new_n543_), .A2(G113gat), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n927_), .B1(new_n929_), .B2(new_n930_), .ZN(G1340gat));
  OAI21_X1  g730(.A(G120gat), .B1(new_n926_), .B2(new_n685_), .ZN(new_n932_));
  INV_X1    g731(.A(G120gat), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n933_), .B1(new_n685_), .B2(KEYINPUT60), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n934_), .B1(KEYINPUT60), .B2(new_n933_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n932_), .B1(new_n929_), .B2(new_n935_), .ZN(G1341gat));
  OAI21_X1  g735(.A(G127gat), .B1(new_n926_), .B2(new_n651_), .ZN(new_n937_));
  OR2_X1    g736(.A1(new_n651_), .A2(G127gat), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n929_), .B2(new_n938_), .ZN(G1342gat));
  AOI21_X1  g738(.A(G134gat), .B1(new_n924_), .B2(new_n705_), .ZN(new_n940_));
  INV_X1    g739(.A(new_n926_), .ZN(new_n941_));
  XOR2_X1   g740(.A(KEYINPUT123), .B(G134gat), .Z(new_n942_));
  NOR2_X1   g741(.A1(new_n743_), .A2(new_n942_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n940_), .B1(new_n941_), .B2(new_n943_), .ZN(G1343gat));
  NOR4_X1   g743(.A1(new_n327_), .A2(new_n729_), .A3(new_n446_), .A4(new_n466_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n928_), .A2(new_n945_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n946_), .A2(new_n543_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(new_n344_), .ZN(G1344gat));
  NOR2_X1   g747(.A1(new_n946_), .A2(new_n685_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n949_), .B(new_n345_), .ZN(G1345gat));
  NOR2_X1   g749(.A1(new_n946_), .A2(new_n651_), .ZN(new_n951_));
  XOR2_X1   g750(.A(KEYINPUT61), .B(G155gat), .Z(new_n952_));
  XNOR2_X1  g751(.A(new_n951_), .B(new_n952_), .ZN(G1346gat));
  OAI21_X1  g752(.A(G162gat), .B1(new_n946_), .B2(new_n743_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n705_), .A2(new_n336_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n954_), .B1(new_n946_), .B2(new_n955_), .ZN(G1347gat));
  NOR2_X1   g755(.A1(new_n467_), .A2(new_n326_), .ZN(new_n957_));
  INV_X1    g756(.A(new_n957_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n958_), .A2(new_n416_), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n913_), .A2(new_n739_), .A3(new_n959_), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n960_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n961_));
  NAND4_X1  g760(.A1(new_n913_), .A2(new_n739_), .A3(new_n242_), .A4(new_n959_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n961_), .A2(new_n962_), .ZN(new_n963_));
  AOI21_X1  g762(.A(KEYINPUT62), .B1(new_n960_), .B2(G169gat), .ZN(new_n964_));
  OAI21_X1  g763(.A(KEYINPUT124), .B1(new_n963_), .B2(new_n964_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n960_), .A2(G169gat), .ZN(new_n966_));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n966_), .A2(new_n967_), .ZN(new_n968_));
  INV_X1    g767(.A(KEYINPUT124), .ZN(new_n969_));
  NAND4_X1  g768(.A1(new_n968_), .A2(new_n969_), .A3(new_n962_), .A4(new_n961_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n965_), .A2(new_n970_), .ZN(G1348gat));
  INV_X1    g770(.A(new_n913_), .ZN(new_n972_));
  INV_X1    g771(.A(new_n959_), .ZN(new_n973_));
  NOR2_X1   g772(.A1(new_n972_), .A2(new_n973_), .ZN(new_n974_));
  AOI21_X1  g773(.A(G176gat), .B1(new_n974_), .B2(new_n686_), .ZN(new_n975_));
  NOR2_X1   g774(.A1(new_n923_), .A2(new_n416_), .ZN(new_n976_));
  NOR3_X1   g775(.A1(new_n958_), .A2(new_n685_), .A3(new_n243_), .ZN(new_n977_));
  AOI21_X1  g776(.A(new_n975_), .B1(new_n976_), .B2(new_n977_), .ZN(G1349gat));
  NAND3_X1  g777(.A1(new_n976_), .A2(new_n701_), .A3(new_n957_), .ZN(new_n979_));
  AND2_X1   g778(.A1(new_n701_), .A2(new_n260_), .ZN(new_n980_));
  AOI22_X1  g779(.A1(new_n979_), .A2(new_n235_), .B1(new_n974_), .B2(new_n980_), .ZN(G1350gat));
  AOI21_X1  g780(.A(new_n236_), .B1(new_n974_), .B2(new_n610_), .ZN(new_n982_));
  NOR4_X1   g781(.A1(new_n972_), .A2(new_n261_), .A3(new_n607_), .A4(new_n973_), .ZN(new_n983_));
  OR2_X1    g782(.A1(new_n982_), .A2(new_n983_), .ZN(G1351gat));
  NAND3_X1  g783(.A1(new_n768_), .A2(new_n327_), .A3(new_n495_), .ZN(new_n985_));
  NOR2_X1   g784(.A1(new_n923_), .A2(new_n985_), .ZN(new_n986_));
  NAND2_X1  g785(.A1(new_n986_), .A2(new_n739_), .ZN(new_n987_));
  XNOR2_X1  g786(.A(new_n987_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g787(.A1(new_n986_), .A2(new_n686_), .ZN(new_n989_));
  XNOR2_X1  g788(.A(new_n989_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g789(.A1(new_n986_), .A2(new_n701_), .ZN(new_n991_));
  XNOR2_X1  g790(.A(KEYINPUT63), .B(G211gat), .ZN(new_n992_));
  NOR2_X1   g791(.A1(new_n991_), .A2(new_n992_), .ZN(new_n993_));
  NOR2_X1   g792(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n994_));
  AOI21_X1  g793(.A(new_n993_), .B1(new_n991_), .B2(new_n994_), .ZN(G1354gat));
  NOR3_X1   g794(.A1(new_n923_), .A2(new_n607_), .A3(new_n985_), .ZN(new_n996_));
  XNOR2_X1  g795(.A(KEYINPUT125), .B(G218gat), .ZN(new_n997_));
  INV_X1    g796(.A(new_n997_), .ZN(new_n998_));
  NOR2_X1   g797(.A1(new_n996_), .A2(new_n998_), .ZN(new_n999_));
  NOR4_X1   g798(.A1(new_n923_), .A2(new_n743_), .A3(new_n985_), .A4(new_n997_), .ZN(new_n1000_));
  OAI21_X1  g799(.A(KEYINPUT126), .B1(new_n999_), .B2(new_n1000_), .ZN(new_n1001_));
  NAND3_X1  g800(.A1(new_n986_), .A2(new_n610_), .A3(new_n998_), .ZN(new_n1002_));
  INV_X1    g801(.A(KEYINPUT126), .ZN(new_n1003_));
  OAI211_X1 g802(.A(new_n1002_), .B(new_n1003_), .C1(new_n996_), .C2(new_n998_), .ZN(new_n1004_));
  NAND2_X1  g803(.A1(new_n1001_), .A2(new_n1004_), .ZN(G1355gat));
endmodule


