//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 0 1 0 0 1 1 0 0 1 1 1 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n776_, new_n777_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n879_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT87), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G211gat), .B(G218gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT88), .ZN(new_n206_));
  OAI211_X1 g005(.A(KEYINPUT21), .B(new_n204_), .C1(new_n205_), .C2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT21), .ZN(new_n208_));
  INV_X1    g007(.A(G218gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G211gat), .ZN(new_n210_));
  INV_X1    g009(.A(G211gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G218gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n208_), .B1(new_n213_), .B2(KEYINPUT88), .ZN(new_n214_));
  AND2_X1   g013(.A1(G197gat), .A2(G204gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G197gat), .A2(G204gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n217_), .B1(new_n205_), .B2(KEYINPUT21), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n207_), .B1(new_n214_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT86), .ZN(new_n220_));
  AND3_X1   g019(.A1(KEYINPUT82), .A2(G155gat), .A3(G162gat), .ZN(new_n221_));
  AOI21_X1  g020(.A(KEYINPUT82), .B1(G155gat), .B2(G162gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT1), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT82), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT1), .ZN(new_n227_));
  NAND3_X1  g026(.A1(KEYINPUT82), .A2(G155gat), .A3(G162gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT81), .ZN(new_n230_));
  INV_X1    g029(.A(G155gat), .ZN(new_n231_));
  INV_X1    g030(.A(G162gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT81), .B1(G155gat), .B2(G162gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n223_), .A2(new_n229_), .A3(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(G141gat), .B(G148gat), .Z(new_n237_));
  AND3_X1   g036(.A1(new_n236_), .A2(KEYINPUT83), .A3(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(KEYINPUT83), .B1(new_n236_), .B2(new_n237_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n235_), .B1(new_n222_), .B2(new_n221_), .ZN(new_n241_));
  INV_X1    g040(.A(G141gat), .ZN(new_n242_));
  INV_X1    g041(.A(G148gat), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT2), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT2), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n245_), .A2(G141gat), .A3(G148gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n242_), .A2(new_n243_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n248_), .B1(KEYINPUT84), .B2(KEYINPUT3), .ZN(new_n249_));
  NOR2_X1   g048(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n250_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n247_), .A2(new_n249_), .A3(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT85), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n248_), .B(new_n250_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(KEYINPUT85), .A3(new_n247_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n241_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n220_), .B1(new_n240_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n241_), .ZN(new_n259_));
  AOI21_X1  g058(.A(KEYINPUT85), .B1(new_n255_), .B2(new_n247_), .ZN(new_n260_));
  AND4_X1   g059(.A1(KEYINPUT85), .A2(new_n247_), .A3(new_n249_), .A4(new_n251_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n259_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n262_), .B(KEYINPUT86), .C1(new_n239_), .C2(new_n238_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n258_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT29), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n203_), .B(new_n219_), .C1(new_n264_), .C2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n219_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n262_), .B1(new_n239_), .B2(new_n238_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n267_), .B1(new_n268_), .B2(KEYINPUT29), .ZN(new_n269_));
  NOR3_X1   g068(.A1(new_n269_), .A2(KEYINPUT89), .A3(new_n203_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT89), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n254_), .A2(new_n256_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n236_), .A2(new_n237_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT83), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n236_), .A2(KEYINPUT83), .A3(new_n237_), .ZN(new_n276_));
  AOI22_X1  g075(.A1(new_n272_), .A2(new_n259_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n219_), .B1(new_n277_), .B2(new_n265_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n203_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n271_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n266_), .B1(new_n270_), .B2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G78gat), .B(G106gat), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT90), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G22gat), .B(G50gat), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n284_), .B(KEYINPUT28), .Z(new_n285_));
  AND3_X1   g084(.A1(new_n264_), .A2(new_n265_), .A3(new_n285_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n285_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT89), .B1(new_n269_), .B2(new_n203_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n278_), .A2(new_n271_), .A3(new_n279_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n282_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n292_), .A2(new_n293_), .A3(new_n266_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n293_), .B1(new_n292_), .B2(new_n266_), .ZN(new_n296_));
  OAI22_X1  g095(.A1(new_n283_), .A2(new_n289_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n296_), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n298_), .A2(new_n294_), .A3(new_n288_), .A4(KEYINPUT90), .ZN(new_n299_));
  XOR2_X1   g098(.A(G1gat), .B(G29gat), .Z(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT94), .B(G85gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT0), .B(G57gat), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n302_), .B(new_n303_), .Z(new_n304_));
  XOR2_X1   g103(.A(G113gat), .B(G120gat), .Z(new_n305_));
  XNOR2_X1  g104(.A(G127gat), .B(G134gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n258_), .A2(new_n263_), .A3(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n307_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n277_), .A2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n308_), .A2(KEYINPUT4), .A3(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G225gat), .A2(G233gat), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n311_), .B(new_n313_), .C1(KEYINPUT4), .C2(new_n308_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n308_), .A2(new_n310_), .A3(new_n312_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n304_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  AND3_X1   g115(.A1(new_n308_), .A2(KEYINPUT4), .A3(new_n310_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n313_), .B1(new_n308_), .B2(KEYINPUT4), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n315_), .B(new_n304_), .C1(new_n317_), .C2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n316_), .A2(new_n320_), .ZN(new_n321_));
  AND3_X1   g120(.A1(new_n297_), .A2(new_n299_), .A3(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT20), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G183gat), .A2(G190gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT78), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT78), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n326_), .A2(G183gat), .A3(G190gat), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n325_), .A2(new_n327_), .A3(KEYINPUT23), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT80), .ZN(new_n329_));
  AND2_X1   g128(.A1(G183gat), .A2(G190gat), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT23), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n329_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n328_), .A2(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(G183gat), .A2(G190gat), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n325_), .A2(new_n327_), .A3(new_n329_), .A4(KEYINPUT23), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n333_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT79), .B(G176gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT22), .B(G169gat), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n338_), .A2(new_n339_), .B1(G169gat), .B2(G176gat), .ZN(new_n340_));
  INV_X1    g139(.A(G183gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT25), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT25), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(G183gat), .ZN(new_n344_));
  INV_X1    g143(.A(G190gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT26), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT26), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(G190gat), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n342_), .A2(new_n344_), .A3(new_n346_), .A4(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(G169gat), .A2(G176gat), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G169gat), .A2(G176gat), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(KEYINPUT24), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT24), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n350_), .A2(new_n354_), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n349_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n330_), .A2(new_n331_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n325_), .A2(new_n327_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n357_), .B1(new_n358_), .B2(new_n331_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  AOI22_X1  g159(.A1(new_n337_), .A2(new_n340_), .B1(new_n356_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n323_), .B1(new_n362_), .B2(new_n219_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G226gat), .A2(G233gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT19), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n340_), .B1(new_n359_), .B2(new_n334_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT25), .B(G183gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT26), .B(G190gat), .ZN(new_n369_));
  AOI22_X1  g168(.A1(new_n368_), .A2(new_n369_), .B1(new_n354_), .B2(new_n350_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n370_), .A2(new_n333_), .A3(new_n353_), .A4(new_n336_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n367_), .A2(new_n371_), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n363_), .B(new_n366_), .C1(new_n219_), .C2(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n323_), .B1(new_n361_), .B2(new_n267_), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n372_), .A2(KEYINPUT91), .A3(new_n219_), .ZN(new_n375_));
  AOI21_X1  g174(.A(KEYINPUT91), .B1(new_n372_), .B2(new_n219_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n374_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT92), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n377_), .A2(new_n378_), .A3(new_n365_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n378_), .B1(new_n377_), .B2(new_n365_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n373_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  XOR2_X1   g180(.A(G8gat), .B(G36gat), .Z(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G64gat), .B(G92gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n381_), .A2(new_n387_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n386_), .B(new_n373_), .C1(new_n379_), .C2(new_n380_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT27), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT101), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT100), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n389_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n337_), .A2(new_n340_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n356_), .A2(new_n360_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n267_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT20), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n372_), .A2(new_n219_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT91), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n372_), .A2(KEYINPUT91), .A3(new_n219_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n399_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT92), .B1(new_n404_), .B2(new_n366_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n377_), .A2(new_n378_), .A3(new_n365_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n407_), .A2(KEYINPUT100), .A3(new_n386_), .A4(new_n373_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n395_), .A2(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n219_), .B1(new_n372_), .B2(KEYINPUT98), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n410_), .B1(KEYINPUT98), .B2(new_n372_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n366_), .B1(new_n411_), .B2(new_n363_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n374_), .B(new_n366_), .C1(new_n375_), .C2(new_n376_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  XOR2_X1   g214(.A(new_n386_), .B(KEYINPUT99), .Z(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT27), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n393_), .B1(new_n409_), .B2(new_n418_), .ZN(new_n419_));
  AOI211_X1 g218(.A(KEYINPUT101), .B(new_n417_), .C1(new_n395_), .C2(new_n408_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n322_), .B(new_n392_), .C1(new_n419_), .C2(new_n420_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n386_), .A2(KEYINPUT32), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n381_), .A2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n422_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n425_), .A2(new_n321_), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n314_), .A2(KEYINPUT33), .A3(new_n315_), .A4(new_n304_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n304_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n308_), .A2(new_n310_), .A3(new_n313_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n312_), .B1(new_n308_), .B2(KEYINPUT4), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n428_), .B(new_n429_), .C1(new_n317_), .C2(new_n430_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n427_), .A2(new_n388_), .A3(new_n389_), .A4(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT95), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n319_), .A2(new_n433_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n314_), .A2(KEYINPUT95), .A3(new_n315_), .A4(new_n304_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(KEYINPUT96), .B(KEYINPUT33), .Z(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n432_), .B1(new_n438_), .B2(KEYINPUT97), .ZN(new_n439_));
  INV_X1    g238(.A(new_n437_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n440_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT97), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n426_), .B1(new_n439_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n297_), .A2(new_n299_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n421_), .B1(new_n444_), .B2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G71gat), .B(G99gat), .ZN(new_n448_));
  INV_X1    g247(.A(G43gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n361_), .B(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(new_n307_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G227gat), .A2(G233gat), .ZN(new_n453_));
  XOR2_X1   g252(.A(new_n453_), .B(G15gat), .Z(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT30), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT31), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n452_), .B(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n392_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT102), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT102), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n460_), .B(new_n392_), .C1(new_n419_), .C2(new_n420_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n457_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n445_), .A2(new_n321_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n447_), .A2(new_n457_), .B1(new_n462_), .B2(new_n465_), .ZN(new_n466_));
  XOR2_X1   g265(.A(G57gat), .B(G64gat), .Z(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT71), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT11), .ZN(new_n469_));
  OR2_X1    g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(G71gat), .B(G78gat), .Z(new_n471_));
  OR2_X1    g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n468_), .A2(new_n469_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n470_), .A2(new_n473_), .A3(new_n471_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT76), .B(G15gat), .ZN(new_n476_));
  INV_X1    g275(.A(G22gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(G1gat), .ZN(new_n479_));
  INV_X1    g278(.A(G8gat), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT14), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n478_), .A2(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(G1gat), .B(G8gat), .Z(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n475_), .B(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G231gat), .A2(G233gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G127gat), .B(G155gat), .Z(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G183gat), .B(G211gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  OR2_X1    g291(.A1(new_n492_), .A2(KEYINPUT17), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT72), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n492_), .A2(new_n494_), .A3(KEYINPUT17), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  OR2_X1    g295(.A1(new_n487_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n487_), .A2(new_n495_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G232gat), .A2(G233gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT34), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G99gat), .A2(G106gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT6), .ZN(new_n504_));
  XNOR2_X1  g303(.A(KEYINPUT10), .B(G99gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT65), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT66), .B(G106gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT67), .B(G92gat), .ZN(new_n509_));
  INV_X1    g308(.A(G85gat), .ZN(new_n510_));
  NOR3_X1   g309(.A1(new_n509_), .A2(KEYINPUT9), .A3(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(G85gat), .B(G92gat), .Z(new_n512_));
  AOI21_X1  g311(.A(new_n511_), .B1(KEYINPUT9), .B2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT68), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n513_), .A2(new_n514_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n504_), .B(new_n508_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(G99gat), .ZN(new_n518_));
  INV_X1    g317(.A(G106gat), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(new_n519_), .A3(KEYINPUT69), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n520_), .A2(KEYINPUT7), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(KEYINPUT7), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n521_), .A2(new_n504_), .A3(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(KEYINPUT70), .B1(new_n523_), .B2(new_n512_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT8), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n523_), .A2(KEYINPUT70), .A3(new_n512_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n524_), .A2(new_n525_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n517_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G29gat), .B(G36gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G43gat), .B(G50gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT15), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n530_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n533_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n530_), .A2(new_n537_), .ZN(new_n538_));
  OAI211_X1 g337(.A(KEYINPUT35), .B(new_n502_), .C1(new_n536_), .C2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n538_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n502_), .A2(KEYINPUT35), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n502_), .A2(KEYINPUT35), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n540_), .A2(new_n541_), .A3(new_n535_), .A4(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G190gat), .B(G218gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G134gat), .B(G162gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n546_), .A2(KEYINPUT36), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n539_), .A2(new_n543_), .A3(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT74), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n539_), .A2(new_n543_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n547_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n546_), .A2(KEYINPUT36), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n550_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n549_), .A2(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n548_), .A2(KEYINPUT74), .ZN(new_n555_));
  OAI21_X1  g354(.A(KEYINPUT37), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n553_), .A2(new_n548_), .ZN(new_n557_));
  XOR2_X1   g356(.A(KEYINPUT75), .B(KEYINPUT37), .Z(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n556_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NOR3_X1   g360(.A1(new_n466_), .A2(new_n500_), .A3(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G230gat), .A2(G233gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT64), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT12), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n566_), .A2(KEYINPUT72), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n530_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n475_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n517_), .A2(new_n528_), .A3(new_n566_), .A4(new_n529_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n568_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n530_), .A2(new_n567_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n573_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n565_), .B1(new_n572_), .B2(new_n574_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n530_), .A2(new_n475_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n530_), .A2(new_n475_), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n576_), .A2(new_n577_), .A3(new_n564_), .ZN(new_n578_));
  XOR2_X1   g377(.A(G120gat), .B(G148gat), .Z(new_n579_));
  XNOR2_X1  g378(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G176gat), .B(G204gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n575_), .A2(new_n578_), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n584_), .B1(new_n575_), .B2(new_n578_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n588_), .A2(KEYINPUT13), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(KEYINPUT13), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n484_), .B(new_n533_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n593_), .A2(G229gat), .A3(G233gat), .ZN(new_n594_));
  INV_X1    g393(.A(new_n534_), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n484_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G229gat), .A2(G233gat), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n484_), .A2(new_n533_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n596_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n594_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G113gat), .B(G141gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G169gat), .B(G197gat), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n602_), .B(new_n603_), .Z(new_n604_));
  OR2_X1    g403(.A1(new_n601_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n601_), .A2(new_n604_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n592_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n562_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n321_), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n611_), .A2(KEYINPUT103), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(KEYINPUT103), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n610_), .A2(G1gat), .A3(new_n614_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n615_), .A2(KEYINPUT38), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(KEYINPUT38), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n466_), .A2(new_n557_), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n618_), .A2(new_n609_), .A3(new_n499_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  OAI21_X1  g419(.A(G1gat), .B1(new_n620_), .B2(new_n321_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n616_), .A2(new_n617_), .A3(new_n621_), .ZN(G1324gat));
  INV_X1    g421(.A(new_n462_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n562_), .A2(new_n480_), .A3(new_n609_), .A4(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n480_), .B1(new_n619_), .B2(new_n623_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT39), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n625_), .A2(new_n626_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n624_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT40), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  OAI211_X1 g431(.A(KEYINPUT40), .B(new_n624_), .C1(new_n628_), .C2(new_n629_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(G1325gat));
  OAI21_X1  g433(.A(G15gat), .B1(new_n620_), .B2(new_n457_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n636_), .ZN(new_n638_));
  OR3_X1    g437(.A1(new_n610_), .A2(G15gat), .A3(new_n457_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n637_), .A2(new_n638_), .A3(new_n639_), .ZN(G1326gat));
  XNOR2_X1  g439(.A(new_n445_), .B(KEYINPUT105), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n562_), .A2(new_n477_), .A3(new_n609_), .A4(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n477_), .B1(new_n619_), .B2(new_n642_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT42), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n644_), .A2(new_n645_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n643_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT106), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  OAI211_X1 g450(.A(KEYINPUT106), .B(new_n643_), .C1(new_n647_), .C2(new_n648_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(G1327gat));
  INV_X1    g452(.A(KEYINPUT108), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT107), .ZN(new_n655_));
  OAI21_X1  g454(.A(KEYINPUT43), .B1(new_n560_), .B2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n657_), .B1(new_n466_), .B2(new_n560_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n426_), .ZN(new_n659_));
  AND4_X1   g458(.A1(new_n427_), .A2(new_n388_), .A3(new_n389_), .A4(new_n431_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n660_), .B1(new_n442_), .B2(new_n441_), .ZN(new_n661_));
  AOI211_X1 g460(.A(KEYINPUT97), .B(new_n440_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n659_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(new_n445_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n463_), .B1(new_n664_), .B2(new_n421_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n464_), .B1(new_n459_), .B2(new_n461_), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n656_), .B(new_n561_), .C1(new_n665_), .C2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n658_), .A2(new_n667_), .ZN(new_n668_));
  AOI211_X1 g467(.A(new_n608_), .B(new_n499_), .C1(new_n589_), .C2(new_n590_), .ZN(new_n669_));
  AOI21_X1  g468(.A(KEYINPUT44), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671_));
  INV_X1    g470(.A(new_n669_), .ZN(new_n672_));
  AOI211_X1 g471(.A(new_n671_), .B(new_n672_), .C1(new_n658_), .C2(new_n667_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n670_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n614_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n654_), .B1(new_n676_), .B2(G29gat), .ZN(new_n677_));
  INV_X1    g476(.A(G29gat), .ZN(new_n678_));
  AOI211_X1 g477(.A(KEYINPUT108), .B(new_n678_), .C1(new_n674_), .C2(new_n675_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n557_), .B(new_n669_), .C1(new_n665_), .C2(new_n666_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n611_), .A2(new_n678_), .ZN(new_n681_));
  OAI22_X1  g480(.A1(new_n677_), .A2(new_n679_), .B1(new_n680_), .B2(new_n681_), .ZN(G1328gat));
  INV_X1    g481(.A(KEYINPUT112), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT110), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n462_), .A2(G36gat), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n684_), .B1(new_n680_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n557_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n438_), .A2(KEYINPUT97), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n689_), .A2(new_n443_), .A3(new_n660_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n446_), .B1(new_n690_), .B2(new_n659_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n322_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n692_), .A2(new_n458_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n457_), .B1(new_n691_), .B2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n462_), .A2(new_n465_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n688_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n696_), .A2(KEYINPUT110), .A3(new_n669_), .A4(new_n685_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n687_), .A2(new_n697_), .ZN(new_n698_));
  XOR2_X1   g497(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n687_), .A2(new_n697_), .A3(new_n699_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n667_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n694_), .A2(new_n695_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n656_), .B1(new_n705_), .B2(new_n561_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n669_), .B1(new_n704_), .B2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(new_n671_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n668_), .A2(KEYINPUT44), .A3(new_n669_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(new_n623_), .A3(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n703_), .B1(new_n710_), .B2(G36gat), .ZN(new_n711_));
  XOR2_X1   g510(.A(KEYINPUT111), .B(KEYINPUT46), .Z(new_n712_));
  OAI21_X1  g511(.A(new_n683_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n712_), .ZN(new_n714_));
  INV_X1    g513(.A(G36gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n674_), .B2(new_n623_), .ZN(new_n716_));
  OAI211_X1 g515(.A(KEYINPUT112), .B(new_n714_), .C1(new_n716_), .C2(new_n703_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n711_), .A2(KEYINPUT46), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n713_), .A2(new_n717_), .A3(new_n718_), .ZN(G1329gat));
  NAND3_X1  g518(.A1(new_n674_), .A2(G43gat), .A3(new_n463_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n449_), .B1(new_n680_), .B2(new_n457_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT113), .Z(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT47), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT47), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n720_), .A2(new_n725_), .A3(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1330gat));
  OR3_X1    g526(.A1(new_n680_), .A2(G50gat), .A3(new_n641_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n674_), .A2(KEYINPUT114), .A3(new_n446_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(G50gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(KEYINPUT114), .B1(new_n674_), .B2(new_n446_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n728_), .B1(new_n730_), .B2(new_n731_), .ZN(G1331gat));
  NOR2_X1   g531(.A1(new_n591_), .A2(new_n607_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n562_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(G57gat), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n734_), .A2(new_n735_), .A3(new_n675_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n618_), .A2(new_n499_), .A3(new_n733_), .ZN(new_n737_));
  OAI21_X1  g536(.A(G57gat), .B1(new_n737_), .B2(new_n321_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1332gat));
  INV_X1    g538(.A(G64gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n734_), .A2(new_n740_), .A3(new_n623_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G64gat), .B1(new_n737_), .B2(new_n462_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT116), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n742_), .B(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(KEYINPUT115), .B(KEYINPUT48), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n744_), .A2(new_n745_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n741_), .B1(new_n746_), .B2(new_n747_), .ZN(G1333gat));
  OAI21_X1  g547(.A(G71gat), .B1(new_n737_), .B2(new_n457_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT49), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n457_), .A2(G71gat), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT117), .Z(new_n752_));
  NAND2_X1  g551(.A1(new_n734_), .A2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n750_), .A2(new_n753_), .ZN(G1334gat));
  OAI21_X1  g553(.A(G78gat), .B1(new_n737_), .B2(new_n641_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT50), .ZN(new_n756_));
  INV_X1    g555(.A(G78gat), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n734_), .A2(new_n757_), .A3(new_n642_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT118), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT118), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n756_), .A2(new_n761_), .A3(new_n758_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1335gat));
  INV_X1    g562(.A(KEYINPUT119), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n668_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n733_), .A2(new_n500_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n658_), .A2(KEYINPUT119), .A3(new_n667_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n765_), .A2(new_n767_), .A3(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(G85gat), .B1(new_n769_), .B2(new_n321_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n767_), .A2(new_n696_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n772_), .A2(new_n510_), .A3(new_n675_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n770_), .A2(new_n773_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT120), .ZN(G1336gat));
  NOR3_X1   g574(.A1(new_n769_), .A2(new_n509_), .A3(new_n462_), .ZN(new_n776_));
  AOI21_X1  g575(.A(G92gat), .B1(new_n772_), .B2(new_n623_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(new_n777_), .ZN(G1337gat));
  OAI21_X1  g577(.A(G99gat), .B1(new_n769_), .B2(new_n457_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n772_), .A2(new_n506_), .A3(new_n463_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT51), .ZN(G1338gat));
  AND3_X1   g581(.A1(new_n772_), .A2(new_n507_), .A3(new_n446_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n766_), .A2(new_n445_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n519_), .B1(new_n668_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n786_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n783_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n789_), .B(new_n791_), .ZN(G1339gat));
  NOR3_X1   g591(.A1(new_n623_), .A2(new_n457_), .A3(new_n614_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n586_), .A2(new_n607_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n572_), .A2(new_n565_), .A3(new_n574_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT55), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n572_), .A2(new_n574_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n564_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n798_), .A2(KEYINPUT55), .A3(new_n564_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n583_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n802_), .A2(KEYINPUT56), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n575_), .B1(KEYINPUT55), .B2(new_n796_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n801_), .ZN(new_n805_));
  OAI211_X1 g604(.A(KEYINPUT56), .B(new_n584_), .C1(new_n804_), .C2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n795_), .B1(new_n803_), .B2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n596_), .A2(new_n598_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n809_), .A2(KEYINPUT122), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n809_), .A2(KEYINPUT122), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n810_), .A2(new_n811_), .A3(new_n597_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n604_), .B1(new_n593_), .B2(new_n597_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n606_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n815_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n557_), .B1(new_n808_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT123), .ZN(new_n819_));
  OAI21_X1  g618(.A(KEYINPUT57), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n584_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT56), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n794_), .B1(new_n823_), .B2(new_n806_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n688_), .B1(new_n824_), .B2(new_n816_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(KEYINPUT123), .A3(new_n826_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n820_), .A2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT125), .B1(new_n802_), .B2(KEYINPUT56), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT124), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n806_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT125), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n821_), .A2(new_n832_), .A3(new_n822_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n802_), .A2(KEYINPUT124), .A3(KEYINPUT56), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n829_), .A2(new_n831_), .A3(new_n833_), .A4(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n815_), .A2(new_n585_), .ZN(new_n836_));
  AOI21_X1  g635(.A(KEYINPUT58), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n837_), .A2(new_n560_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n835_), .A2(KEYINPUT58), .A3(new_n836_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n499_), .B1(new_n828_), .B2(new_n840_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n591_), .A2(new_n608_), .A3(new_n499_), .A4(new_n560_), .ZN(new_n842_));
  XOR2_X1   g641(.A(new_n842_), .B(KEYINPUT54), .Z(new_n843_));
  OAI211_X1 g642(.A(new_n445_), .B(new_n793_), .C1(new_n841_), .C2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(G113gat), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n846_), .A3(new_n607_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT59), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT126), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n844_), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n839_), .ZN(new_n851_));
  NOR3_X1   g650(.A1(new_n851_), .A2(new_n837_), .A3(new_n560_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n820_), .A2(new_n827_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n500_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n843_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n446_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n856_), .A2(KEYINPUT126), .A3(KEYINPUT59), .A4(new_n793_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n608_), .B1(new_n850_), .B2(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n847_), .B1(new_n858_), .B2(new_n846_), .ZN(G1340gat));
  INV_X1    g658(.A(G120gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n591_), .B2(KEYINPUT60), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n845_), .B(new_n861_), .C1(KEYINPUT60), .C2(new_n860_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n591_), .B1(new_n850_), .B2(new_n857_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n863_), .B2(new_n860_), .ZN(G1341gat));
  INV_X1    g663(.A(G127gat), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n845_), .A2(new_n865_), .A3(new_n499_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n500_), .B1(new_n850_), .B2(new_n857_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n867_), .B2(new_n865_), .ZN(G1342gat));
  INV_X1    g667(.A(G134gat), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n845_), .A2(new_n869_), .A3(new_n557_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n560_), .B1(new_n850_), .B2(new_n857_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n871_), .B2(new_n869_), .ZN(G1343gat));
  AOI21_X1  g671(.A(new_n463_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n623_), .A2(new_n445_), .A3(new_n614_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n608_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(KEYINPUT127), .B(G141gat), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n876_), .B(new_n877_), .ZN(G1344gat));
  NOR2_X1   g677(.A1(new_n875_), .A2(new_n591_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(new_n243_), .ZN(G1345gat));
  NAND3_X1  g679(.A1(new_n873_), .A2(new_n499_), .A3(new_n874_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(KEYINPUT61), .B(G155gat), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n881_), .B(new_n882_), .ZN(G1346gat));
  OAI21_X1  g682(.A(G162gat), .B1(new_n875_), .B2(new_n560_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n557_), .A2(new_n232_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n875_), .B2(new_n885_), .ZN(G1347gat));
  INV_X1    g685(.A(KEYINPUT62), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n854_), .A2(new_n855_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n623_), .A2(new_n463_), .A3(new_n614_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n889_), .A2(new_n642_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n608_), .ZN(new_n892_));
  INV_X1    g691(.A(G169gat), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n887_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n339_), .ZN(new_n895_));
  OAI211_X1 g694(.A(KEYINPUT62), .B(G169gat), .C1(new_n891_), .C2(new_n608_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n894_), .A2(new_n895_), .A3(new_n896_), .ZN(G1348gat));
  INV_X1    g696(.A(new_n891_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n592_), .ZN(new_n899_));
  AOI211_X1 g698(.A(new_n446_), .B(new_n889_), .C1(new_n854_), .C2(new_n855_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n592_), .A2(G176gat), .ZN(new_n901_));
  AOI22_X1  g700(.A1(new_n899_), .A2(new_n338_), .B1(new_n900_), .B2(new_n901_), .ZN(G1349gat));
  AOI21_X1  g701(.A(G183gat), .B1(new_n900_), .B2(new_n499_), .ZN(new_n903_));
  NOR3_X1   g702(.A1(new_n891_), .A2(new_n368_), .A3(new_n500_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1350gat));
  OAI21_X1  g704(.A(G190gat), .B1(new_n891_), .B2(new_n560_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n557_), .A2(new_n369_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n891_), .B2(new_n907_), .ZN(G1351gat));
  NAND3_X1  g707(.A1(new_n873_), .A2(new_n322_), .A3(new_n623_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n909_), .A2(new_n608_), .ZN(new_n910_));
  INV_X1    g709(.A(G197gat), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n910_), .B(new_n911_), .ZN(G1352gat));
  NOR2_X1   g711(.A1(new_n909_), .A2(new_n591_), .ZN(new_n913_));
  INV_X1    g712(.A(G204gat), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n913_), .B(new_n914_), .ZN(G1353gat));
  XNOR2_X1  g714(.A(KEYINPUT63), .B(G211gat), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n909_), .A2(new_n500_), .A3(new_n916_), .ZN(new_n917_));
  OR2_X1    g716(.A1(new_n909_), .A2(new_n500_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n917_), .B1(new_n918_), .B2(new_n919_), .ZN(G1354gat));
  OAI21_X1  g719(.A(G218gat), .B1(new_n909_), .B2(new_n560_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n557_), .A2(new_n209_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n909_), .B2(new_n922_), .ZN(G1355gat));
endmodule


