//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_, new_n946_,
    new_n948_, new_n949_, new_n951_, new_n952_, new_n953_, new_n954_,
    new_n955_, new_n956_, new_n957_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n969_, new_n970_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n977_, new_n978_, new_n979_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n205_), .A2(KEYINPUT36), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(KEYINPUT36), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT66), .B(KEYINPUT34), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G232gat), .A2(G233gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT35), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n211_), .A2(KEYINPUT35), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT7), .ZN(new_n216_));
  INV_X1    g015(.A(G99gat), .ZN(new_n217_));
  INV_X1    g016(.A(G106gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT6), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n219_), .A2(new_n222_), .A3(new_n223_), .A4(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT8), .ZN(new_n226_));
  INV_X1    g025(.A(G85gat), .ZN(new_n227_));
  INV_X1    g026(.A(G92gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G85gat), .A2(G92gat), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  AND3_X1   g030(.A1(new_n225_), .A2(new_n226_), .A3(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n226_), .B1(new_n225_), .B2(new_n231_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT10), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n234_), .A2(G99gat), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n217_), .A2(KEYINPUT10), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT64), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n217_), .A2(KEYINPUT10), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n234_), .A2(G99gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT64), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n238_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(G106gat), .B1(new_n237_), .B2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n229_), .A2(KEYINPUT9), .A3(new_n230_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n230_), .A2(KEYINPUT9), .ZN(new_n244_));
  NAND4_X1  g043(.A1(new_n243_), .A2(new_n244_), .A3(new_n222_), .A4(new_n223_), .ZN(new_n245_));
  OAI22_X1  g044(.A1(new_n232_), .A2(new_n233_), .B1(new_n242_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G29gat), .B(G36gat), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G43gat), .B(G50gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n250_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(new_n248_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n215_), .B1(new_n247_), .B2(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n214_), .B1(new_n256_), .B2(KEYINPUT68), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT65), .B1(new_n232_), .B2(new_n233_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n225_), .A2(new_n231_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT8), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT65), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n225_), .A2(new_n226_), .A3(new_n231_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n260_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n241_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n240_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n218_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n245_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n258_), .A2(new_n263_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT15), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n254_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n251_), .A2(new_n253_), .A3(KEYINPUT15), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n269_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n256_), .A2(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n257_), .A2(new_n275_), .ZN(new_n276_));
  OAI22_X1  g075(.A1(new_n246_), .A2(new_n254_), .B1(KEYINPUT35), .B2(new_n211_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n277_), .B1(new_n273_), .B2(new_n269_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n212_), .B(KEYINPUT67), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n279_), .B1(new_n277_), .B2(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n207_), .B(new_n208_), .C1(new_n276_), .C2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT69), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n257_), .A2(new_n275_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n278_), .A2(new_n281_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n286_), .A2(new_n287_), .A3(new_n206_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n206_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n289_), .A2(KEYINPUT69), .A3(new_n208_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n285_), .A2(new_n288_), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT37), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n283_), .A2(KEYINPUT37), .A3(new_n288_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G57gat), .B(G64gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT11), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G71gat), .B(G78gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT11), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n296_), .B(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n299_), .B1(new_n301_), .B2(new_n298_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n269_), .A2(KEYINPUT12), .A3(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT12), .B1(new_n246_), .B2(new_n302_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n246_), .A2(new_n302_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G230gat), .A2(G233gat), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n303_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n305_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n246_), .A2(new_n302_), .ZN(new_n310_));
  OAI211_X1 g109(.A(G230gat), .B(G233gat), .C1(new_n309_), .C2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n308_), .A2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT5), .B(G176gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(G204gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G120gat), .B(G148gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n312_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n308_), .A2(new_n311_), .A3(new_n316_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT13), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n318_), .A2(KEYINPUT13), .A3(new_n319_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G15gat), .B(G22gat), .ZN(new_n325_));
  INV_X1    g124(.A(G1gat), .ZN(new_n326_));
  INV_X1    g125(.A(G8gat), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT14), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n325_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G1gat), .B(G8gat), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n330_), .ZN(new_n332_));
  INV_X1    g131(.A(G231gat), .ZN(new_n333_));
  INV_X1    g132(.A(G233gat), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n331_), .A2(new_n332_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n336_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n302_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n339_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n302_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n341_), .A2(new_n342_), .A3(new_n337_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n340_), .A2(new_n343_), .A3(KEYINPUT71), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT17), .ZN(new_n345_));
  XOR2_X1   g144(.A(G183gat), .B(G211gat), .Z(new_n346_));
  XNOR2_X1  g145(.A(G127gat), .B(G155gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT70), .B(KEYINPUT16), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n344_), .A2(new_n345_), .A3(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n344_), .A2(new_n350_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n350_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n354_), .A2(new_n340_), .A3(new_n343_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT17), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n351_), .B1(new_n353_), .B2(new_n356_), .ZN(new_n357_));
  NOR3_X1   g156(.A1(new_n295_), .A2(new_n324_), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT72), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G169gat), .A2(G176gat), .ZN(new_n361_));
  INV_X1    g160(.A(G169gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT22), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT76), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n362_), .A2(KEYINPUT76), .A3(KEYINPUT22), .ZN(new_n366_));
  INV_X1    g165(.A(G176gat), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT22), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(G169gat), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n365_), .A2(new_n366_), .A3(new_n367_), .A4(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT23), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n371_), .B1(G183gat), .B2(G190gat), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(G183gat), .A3(G190gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT77), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT77), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n375_), .A2(new_n371_), .A3(G183gat), .A4(G190gat), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n372_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT75), .B(G190gat), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n378_), .A2(G183gat), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n361_), .B(new_n370_), .C1(new_n377_), .C2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(KEYINPUT25), .B(G183gat), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT26), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(G190gat), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n381_), .B(new_n383_), .C1(new_n378_), .C2(new_n382_), .ZN(new_n384_));
  INV_X1    g183(.A(G183gat), .ZN(new_n385_));
  INV_X1    g184(.A(G190gat), .ZN(new_n386_));
  OAI21_X1  g185(.A(KEYINPUT23), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n373_), .ZN(new_n388_));
  NOR3_X1   g187(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n389_), .B1(new_n391_), .B2(new_n361_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n384_), .A2(new_n388_), .A3(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n380_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(G197gat), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n395_), .A2(G204gat), .ZN(new_n396_));
  INV_X1    g195(.A(G204gat), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n397_), .A2(G197gat), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT21), .B1(new_n396_), .B2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G211gat), .B(G218gat), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT84), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n401_), .A2(new_n397_), .A3(G197gat), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT84), .B1(new_n395_), .B2(G204gat), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n402_), .B1(new_n403_), .B2(new_n396_), .ZN(new_n404_));
  XOR2_X1   g203(.A(KEYINPUT85), .B(KEYINPUT21), .Z(new_n405_));
  OAI211_X1 g204(.A(new_n399_), .B(new_n400_), .C1(new_n404_), .C2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n400_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n404_), .A2(new_n407_), .A3(KEYINPUT21), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n406_), .A2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT20), .B1(new_n394_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT86), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G226gat), .A2(G233gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT19), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n387_), .A2(new_n373_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(G183gat), .A2(G190gat), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT89), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT88), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n363_), .A2(new_n369_), .A3(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n419_), .B1(new_n363_), .B2(new_n369_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n367_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT89), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n388_), .B(new_n423_), .C1(G183gat), .C2(G190gat), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n418_), .A2(new_n422_), .A3(new_n361_), .A4(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n377_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n386_), .A2(KEYINPUT26), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n383_), .A2(new_n427_), .A3(KEYINPUT87), .ZN(new_n428_));
  AOI21_X1  g227(.A(KEYINPUT87), .B1(new_n383_), .B2(new_n427_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n381_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n426_), .A2(new_n430_), .A3(new_n392_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n425_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n409_), .ZN(new_n433_));
  OAI211_X1 g232(.A(KEYINPUT86), .B(KEYINPUT20), .C1(new_n394_), .C2(new_n409_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n412_), .A2(new_n415_), .A3(new_n433_), .A4(new_n434_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n406_), .A2(new_n408_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(new_n425_), .A3(new_n431_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n394_), .A2(new_n409_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(KEYINPUT20), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n414_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n435_), .A2(KEYINPUT94), .A3(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G8gat), .B(G36gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(G92gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT18), .B(G64gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  XOR2_X1   g244(.A(new_n445_), .B(KEYINPUT95), .Z(new_n446_));
  OAI211_X1 g245(.A(new_n441_), .B(new_n446_), .C1(KEYINPUT94), .C2(new_n435_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n437_), .A2(new_n438_), .A3(KEYINPUT20), .A4(new_n415_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT90), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n412_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n414_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n445_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n449_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n447_), .A2(KEYINPUT27), .A3(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n451_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT90), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n448_), .B(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n445_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(KEYINPUT27), .B1(new_n458_), .B2(new_n453_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n454_), .A2(new_n459_), .ZN(new_n460_));
  OR3_X1    g259(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT2), .ZN(new_n462_));
  INV_X1    g261(.A(G141gat), .ZN(new_n463_));
  INV_X1    g262(.A(G148gat), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n462_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n461_), .A2(new_n465_), .A3(new_n466_), .A4(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT78), .ZN(new_n469_));
  INV_X1    g268(.A(G155gat), .ZN(new_n470_));
  INV_X1    g269(.A(G162gat), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n469_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT78), .B1(G155gat), .B2(G162gat), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G155gat), .A2(G162gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n468_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(G141gat), .B(G148gat), .Z(new_n478_));
  NAND2_X1  g277(.A1(new_n475_), .A2(KEYINPUT1), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT79), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT79), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n475_), .A2(new_n481_), .A3(KEYINPUT1), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n472_), .B(new_n473_), .C1(KEYINPUT1), .C2(new_n475_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n478_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT80), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT80), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n487_), .B(new_n478_), .C1(new_n483_), .C2(new_n484_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n477_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT29), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n409_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT83), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT83), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n493_), .B(new_n409_), .C1(new_n489_), .C2(new_n490_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT82), .B(KEYINPUT28), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT81), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n497_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n492_), .A2(new_n494_), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G78gat), .B(G106gat), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(G228gat), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n504_), .A2(new_n334_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n489_), .A2(new_n490_), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n506_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n503_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n486_), .A2(new_n488_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(new_n476_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n505_), .B1(new_n512_), .B2(KEYINPUT29), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n513_), .A2(new_n502_), .A3(new_n507_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G22gat), .B(G50gat), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n510_), .A2(new_n514_), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n516_), .B1(new_n510_), .B2(new_n514_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n501_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NOR3_X1   g319(.A1(new_n508_), .A2(new_n503_), .A3(new_n509_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n502_), .B1(new_n513_), .B2(new_n507_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n515_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n523_), .A2(new_n500_), .A3(new_n517_), .A4(new_n498_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n520_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(G15gat), .B(G43gat), .Z(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT31), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n394_), .B(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G127gat), .B(G134gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G113gat), .B(G120gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(G71gat), .ZN(new_n534_));
  AND2_X1   g333(.A1(G227gat), .A2(G233gat), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n534_), .A2(new_n535_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT30), .B(G99gat), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n537_), .A2(new_n538_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n540_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n530_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n543_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n545_), .A2(new_n529_), .A3(new_n541_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(KEYINPUT92), .B(KEYINPUT0), .Z(new_n548_));
  XNOR2_X1  g347(.A(G1gat), .B(G29gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G57gat), .B(G85gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT91), .ZN(new_n553_));
  INV_X1    g352(.A(new_n533_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n512_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT4), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n556_), .B1(new_n489_), .B2(new_n533_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G225gat), .A2(G233gat), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n512_), .A2(new_n553_), .A3(new_n556_), .A4(new_n554_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n558_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n512_), .A2(new_n554_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n489_), .A2(new_n533_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n563_), .A2(new_n559_), .A3(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n552_), .B1(new_n562_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n562_), .A2(new_n565_), .A3(new_n552_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n547_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n460_), .A2(KEYINPUT96), .A3(new_n526_), .A4(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT96), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT27), .ZN(new_n573_));
  INV_X1    g372(.A(new_n453_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n452_), .B1(new_n449_), .B2(new_n451_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n573_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n447_), .A2(KEYINPUT27), .A3(new_n453_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n562_), .A2(new_n565_), .A3(new_n552_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n579_), .A2(new_n566_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n580_), .A2(new_n520_), .A3(new_n524_), .A4(new_n547_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n572_), .B1(new_n578_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n571_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n547_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n525_), .A2(new_n580_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n586_), .A2(new_n578_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n568_), .A2(KEYINPUT33), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT33), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n562_), .A2(new_n589_), .A3(new_n565_), .A4(new_n552_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  AND3_X1   g390(.A1(new_n563_), .A2(KEYINPUT93), .A3(new_n564_), .ZN(new_n592_));
  AOI21_X1  g391(.A(KEYINPUT93), .B1(new_n563_), .B2(new_n564_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n560_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n552_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n558_), .A2(new_n559_), .A3(new_n561_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n594_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n591_), .A2(new_n453_), .A3(new_n458_), .A4(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n452_), .A2(KEYINPUT32), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n449_), .A2(new_n451_), .A3(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n441_), .B1(KEYINPUT94), .B2(new_n435_), .ZN(new_n601_));
  OAI221_X1 g400(.A(new_n600_), .B1(new_n601_), .B2(new_n599_), .C1(new_n566_), .C2(new_n579_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n525_), .B1(new_n598_), .B2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n585_), .B1(new_n587_), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n584_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n331_), .A2(new_n332_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n273_), .A2(KEYINPUT73), .A3(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G229gat), .A2(G233gat), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT73), .ZN(new_n609_));
  INV_X1    g408(.A(new_n606_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n609_), .B1(new_n610_), .B2(new_n255_), .ZN(new_n611_));
  AOI22_X1  g410(.A1(new_n271_), .A2(new_n272_), .B1(new_n332_), .B2(new_n331_), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n607_), .B(new_n608_), .C1(new_n611_), .C2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n606_), .B(new_n254_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n608_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n613_), .A2(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(G113gat), .B(G141gat), .Z(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT74), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G169gat), .B(G197gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n617_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n613_), .A2(new_n616_), .A3(new_n621_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n626_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n360_), .A2(new_n605_), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n580_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(new_n326_), .A3(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT38), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT98), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n324_), .A2(new_n626_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n351_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n356_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n634_), .B1(new_n352_), .B2(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT97), .B1(new_n605_), .B2(new_n291_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT97), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n285_), .A2(new_n288_), .A3(new_n290_), .ZN(new_n639_));
  AOI211_X1 g438(.A(new_n638_), .B(new_n639_), .C1(new_n584_), .C2(new_n604_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n633_), .B(new_n636_), .C1(new_n637_), .C2(new_n640_), .ZN(new_n641_));
  OAI211_X1 g440(.A(new_n632_), .B(G1gat), .C1(new_n641_), .C2(new_n580_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n598_), .A2(new_n602_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(new_n526_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n460_), .A2(new_n580_), .A3(new_n525_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n583_), .B1(new_n647_), .B2(new_n585_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n638_), .B1(new_n648_), .B2(new_n639_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n605_), .A2(KEYINPUT97), .A3(new_n291_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n651_), .A2(new_n629_), .A3(new_n633_), .A4(new_n636_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n632_), .B1(new_n652_), .B2(G1gat), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n631_), .B1(new_n643_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT99), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  OAI211_X1 g455(.A(KEYINPUT99), .B(new_n631_), .C1(new_n643_), .C2(new_n653_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1324gat));
  OAI21_X1  g457(.A(G8gat), .B1(new_n641_), .B2(new_n460_), .ZN(new_n659_));
  XOR2_X1   g458(.A(KEYINPUT100), .B(KEYINPUT39), .Z(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n628_), .A2(new_n327_), .A3(new_n578_), .ZN(new_n663_));
  OAI211_X1 g462(.A(G8gat), .B(new_n660_), .C1(new_n641_), .C2(new_n460_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n662_), .A2(new_n663_), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT40), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n662_), .A2(KEYINPUT40), .A3(new_n663_), .A4(new_n664_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1325gat));
  INV_X1    g468(.A(G15gat), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n628_), .A2(new_n670_), .A3(new_n547_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n357_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n672_), .A2(new_n633_), .A3(new_n547_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(KEYINPUT101), .B(KEYINPUT41), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(G15gat), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n674_), .B1(new_n673_), .B2(G15gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n671_), .B1(new_n676_), .B2(new_n677_), .ZN(G1326gat));
  INV_X1    g477(.A(G22gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n628_), .A2(new_n679_), .A3(new_n525_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n672_), .A2(new_n633_), .A3(new_n525_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT42), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n681_), .A2(new_n682_), .A3(G22gat), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n682_), .B1(new_n681_), .B2(G22gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n680_), .B1(new_n684_), .B2(new_n685_), .ZN(G1327gat));
  NAND2_X1  g485(.A1(KEYINPUT102), .A2(KEYINPUT43), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(KEYINPUT102), .A2(KEYINPUT43), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n295_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n690_), .B1(new_n648_), .B2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n633_), .A2(new_n357_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n547_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n295_), .B(new_n688_), .C1(new_n695_), .C2(new_n583_), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n692_), .A2(KEYINPUT44), .A3(new_n694_), .A4(new_n696_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n697_), .A2(G29gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n691_), .B1(new_n584_), .B2(new_n604_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n690_), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n696_), .B(new_n694_), .C1(new_n699_), .C2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT103), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n701_), .A2(new_n702_), .A3(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n702_), .B1(new_n701_), .B2(new_n703_), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n698_), .B(new_n629_), .C1(new_n705_), .C2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(G29gat), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n648_), .A2(new_n291_), .A3(new_n693_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n708_), .B1(new_n710_), .B2(new_n580_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n707_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT104), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT104), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n707_), .A2(new_n714_), .A3(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1328gat));
  INV_X1    g515(.A(G36gat), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n460_), .B(KEYINPUT105), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n709_), .A2(new_n717_), .A3(new_n718_), .ZN(new_n719_));
  XOR2_X1   g518(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n720_));
  XNOR2_X1  g519(.A(new_n719_), .B(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n697_), .A2(new_n578_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n701_), .A2(new_n703_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT103), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n722_), .B1(new_n724_), .B2(new_n704_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n721_), .B1(new_n725_), .B2(new_n717_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT46), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  OAI211_X1 g527(.A(KEYINPUT46), .B(new_n721_), .C1(new_n725_), .C2(new_n717_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1329gat));
  AND2_X1   g529(.A1(new_n697_), .A2(G43gat), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n731_), .B(new_n547_), .C1(new_n705_), .C2(new_n706_), .ZN(new_n732_));
  INV_X1    g531(.A(G43gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n733_), .B1(new_n710_), .B2(new_n585_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT47), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT47), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n732_), .A2(new_n737_), .A3(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1330gat));
  INV_X1    g538(.A(G50gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n709_), .A2(new_n740_), .A3(new_n525_), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n525_), .B(new_n697_), .C1(new_n705_), .C2(new_n706_), .ZN(new_n742_));
  AOI21_X1  g541(.A(KEYINPUT107), .B1(new_n742_), .B2(G50gat), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n697_), .A2(new_n525_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n744_), .B1(new_n724_), .B2(new_n704_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n745_), .A2(new_n746_), .A3(new_n740_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n741_), .B1(new_n743_), .B2(new_n747_), .ZN(G1331gat));
  INV_X1    g547(.A(new_n324_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n749_), .A2(new_n625_), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n672_), .A2(G57gat), .A3(new_n629_), .A4(new_n750_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n751_), .A2(KEYINPUT109), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n751_), .A2(KEYINPUT109), .ZN(new_n753_));
  INV_X1    g552(.A(new_n750_), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n754_), .A2(new_n357_), .A3(new_n295_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n605_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT108), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n629_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n757_), .B2(new_n756_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n759_), .A2(G57gat), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n752_), .A2(new_n753_), .A3(new_n760_), .ZN(G1332gat));
  INV_X1    g560(.A(new_n718_), .ZN(new_n762_));
  OR3_X1    g561(.A1(new_n756_), .A2(G64gat), .A3(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n651_), .A2(new_n636_), .A3(new_n750_), .ZN(new_n764_));
  OAI21_X1  g563(.A(G64gat), .B1(new_n764_), .B2(new_n762_), .ZN(new_n765_));
  OR2_X1    g564(.A1(new_n765_), .A2(KEYINPUT48), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n765_), .A2(KEYINPUT48), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n763_), .B1(new_n767_), .B2(new_n768_), .ZN(G1333gat));
  INV_X1    g568(.A(KEYINPUT49), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n672_), .A2(new_n547_), .A3(new_n750_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT110), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n772_), .A3(G71gat), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n772_), .B1(new_n771_), .B2(G71gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n770_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n775_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n777_), .A2(KEYINPUT49), .A3(new_n773_), .ZN(new_n778_));
  OR3_X1    g577(.A1(new_n756_), .A2(G71gat), .A3(new_n585_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n776_), .A2(new_n778_), .A3(new_n779_), .ZN(G1334gat));
  OAI21_X1  g579(.A(G78gat), .B1(new_n764_), .B2(new_n526_), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n781_), .A2(KEYINPUT50), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n781_), .A2(KEYINPUT50), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n526_), .A2(G78gat), .ZN(new_n785_));
  XOR2_X1   g584(.A(new_n785_), .B(KEYINPUT111), .Z(new_n786_));
  OAI22_X1  g585(.A1(new_n783_), .A2(new_n784_), .B1(new_n756_), .B2(new_n786_), .ZN(G1335gat));
  NAND2_X1  g586(.A1(new_n692_), .A2(new_n696_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT112), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n754_), .A2(new_n636_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT112), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n692_), .A2(new_n791_), .A3(new_n696_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n789_), .A2(new_n790_), .A3(new_n792_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n580_), .A2(new_n227_), .ZN(new_n794_));
  XOR2_X1   g593(.A(new_n794_), .B(KEYINPUT113), .Z(new_n795_));
  NOR2_X1   g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n648_), .A2(new_n291_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n790_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(G85gat), .B1(new_n799_), .B2(new_n629_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n796_), .A2(new_n800_), .ZN(G1336gat));
  OAI21_X1  g600(.A(new_n228_), .B1(new_n798_), .B2(new_n460_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n789_), .A2(G92gat), .A3(new_n790_), .A4(new_n792_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n803_), .B2(new_n762_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n804_), .B(new_n805_), .ZN(G1337gat));
  OAI21_X1  g605(.A(G99gat), .B1(new_n793_), .B2(new_n585_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n799_), .B(new_n547_), .C1(new_n265_), .C2(new_n264_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT51), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n807_), .A2(new_n811_), .A3(new_n808_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(G1338gat));
  NAND3_X1  g612(.A1(new_n799_), .A2(new_n218_), .A3(new_n525_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n692_), .A2(new_n525_), .A3(new_n696_), .A4(new_n790_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n815_), .A2(new_n816_), .A3(G106gat), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n816_), .B1(new_n815_), .B2(G106gat), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n814_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR3_X1   g619(.A1(new_n578_), .A2(new_n580_), .A3(new_n585_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n307_), .B1(new_n303_), .B2(new_n306_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n308_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n303_), .A2(new_n306_), .A3(KEYINPUT55), .A4(new_n307_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n316_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT56), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n319_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  AOI211_X1 g627(.A(KEYINPUT56), .B(new_n316_), .C1(new_n824_), .C2(new_n825_), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n828_), .A2(new_n626_), .A3(new_n829_), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n607_), .B(new_n615_), .C1(new_n611_), .C2(new_n612_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n614_), .A2(new_n608_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n622_), .A3(new_n832_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n624_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n320_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(KEYINPUT117), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n837_));
  INV_X1    g636(.A(new_n319_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n316_), .B1(new_n308_), .B2(new_n311_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n834_), .B(new_n837_), .C1(new_n838_), .C2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n836_), .A2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n291_), .B1(new_n830_), .B2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT118), .ZN(new_n843_));
  XNOR2_X1  g642(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n824_), .A2(new_n825_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n317_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT56), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n826_), .A2(new_n827_), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n847_), .A2(new_n625_), .A3(new_n319_), .A4(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n840_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n837_), .B1(new_n320_), .B2(new_n834_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n849_), .A2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT118), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n854_), .A3(new_n291_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n843_), .A2(new_n844_), .A3(new_n855_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n847_), .A2(new_n319_), .A3(new_n848_), .A4(new_n834_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT58), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n828_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n860_), .A2(KEYINPUT58), .A3(new_n848_), .A4(new_n834_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n859_), .A2(new_n295_), .A3(new_n861_), .ZN(new_n862_));
  OAI211_X1 g661(.A(KEYINPUT57), .B(new_n291_), .C1(new_n830_), .C2(new_n841_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n636_), .B1(new_n856_), .B2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n626_), .A2(new_n636_), .A3(KEYINPUT115), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT115), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n867_), .B1(new_n357_), .B2(new_n625_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(KEYINPUT116), .B1(new_n869_), .B2(new_n324_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT116), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n749_), .A2(new_n871_), .A3(new_n868_), .A4(new_n866_), .ZN(new_n872_));
  AOI211_X1 g671(.A(KEYINPUT54), .B(new_n295_), .C1(new_n870_), .C2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n872_), .A2(new_n870_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(new_n691_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n873_), .A2(new_n876_), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n526_), .B(new_n821_), .C1(new_n865_), .C2(new_n877_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(KEYINPUT59), .ZN(new_n879_));
  INV_X1    g678(.A(G113gat), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n879_), .A2(new_n880_), .A3(new_n626_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT121), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT120), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n878_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n878_), .A2(new_n883_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n626_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n882_), .B1(new_n886_), .B2(G113gat), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n878_), .B(KEYINPUT120), .ZN(new_n888_));
  OAI211_X1 g687(.A(KEYINPUT121), .B(new_n880_), .C1(new_n888_), .C2(new_n626_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n881_), .B1(new_n887_), .B2(new_n889_), .ZN(G1340gat));
  NAND2_X1  g689(.A1(new_n884_), .A2(new_n885_), .ZN(new_n891_));
  INV_X1    g690(.A(G120gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n892_), .B1(new_n749_), .B2(KEYINPUT60), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n891_), .B(new_n893_), .C1(KEYINPUT60), .C2(new_n892_), .ZN(new_n894_));
  OAI21_X1  g693(.A(G120gat), .B1(new_n879_), .B2(new_n749_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1341gat));
  AOI21_X1  g695(.A(G127gat), .B1(new_n891_), .B2(new_n636_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n879_), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n636_), .A2(G127gat), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n897_), .B1(new_n898_), .B2(new_n899_), .ZN(G1342gat));
  INV_X1    g699(.A(G134gat), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n879_), .A2(new_n901_), .A3(new_n691_), .ZN(new_n902_));
  AOI21_X1  g701(.A(G134gat), .B1(new_n891_), .B2(new_n639_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1343gat));
  NAND2_X1  g703(.A1(new_n862_), .A2(new_n863_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n854_), .B1(new_n853_), .B2(new_n291_), .ZN(new_n906_));
  AOI211_X1 g705(.A(KEYINPUT118), .B(new_n639_), .C1(new_n849_), .C2(new_n852_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n905_), .B1(new_n908_), .B2(new_n844_), .ZN(new_n909_));
  OAI22_X1  g708(.A1(new_n909_), .A2(new_n636_), .B1(new_n876_), .B2(new_n873_), .ZN(new_n910_));
  AND2_X1   g709(.A1(new_n910_), .A2(new_n585_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n718_), .A2(new_n580_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n911_), .A2(new_n525_), .A3(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n914_), .A2(new_n463_), .A3(new_n625_), .ZN(new_n915_));
  OAI21_X1  g714(.A(G141gat), .B1(new_n913_), .B2(new_n626_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1344gat));
  XNOR2_X1  g716(.A(KEYINPUT122), .B(G148gat), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n914_), .A2(new_n324_), .A3(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n918_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n920_), .B1(new_n913_), .B2(new_n749_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n919_), .A2(new_n921_), .ZN(G1345gat));
  XNOR2_X1  g721(.A(KEYINPUT61), .B(G155gat), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n923_), .B1(new_n914_), .B2(new_n636_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n923_), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n913_), .A2(new_n357_), .A3(new_n925_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n924_), .A2(new_n926_), .ZN(G1346gat));
  NOR3_X1   g726(.A1(new_n913_), .A2(new_n471_), .A3(new_n691_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n914_), .A2(new_n639_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n928_), .B1(new_n471_), .B2(new_n929_), .ZN(G1347gat));
  NAND2_X1  g729(.A1(new_n910_), .A2(new_n526_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n420_), .A2(new_n421_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n762_), .A2(new_n569_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(new_n625_), .ZN(new_n934_));
  OR3_X1    g733(.A1(new_n931_), .A2(new_n932_), .A3(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n936_));
  OAI211_X1 g735(.A(new_n910_), .B(new_n526_), .C1(KEYINPUT123), .C2(new_n934_), .ZN(new_n937_));
  AND2_X1   g736(.A1(new_n934_), .A2(KEYINPUT123), .ZN(new_n938_));
  OR2_X1    g737(.A1(new_n937_), .A2(new_n938_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n936_), .B1(new_n939_), .B2(G169gat), .ZN(new_n940_));
  OAI211_X1 g739(.A(new_n936_), .B(G169gat), .C1(new_n937_), .C2(new_n938_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n941_), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n935_), .B1(new_n940_), .B2(new_n942_), .ZN(G1348gat));
  OAI211_X1 g742(.A(new_n526_), .B(new_n933_), .C1(new_n865_), .C2(new_n877_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n944_), .A2(new_n749_), .ZN(new_n945_));
  XOR2_X1   g744(.A(KEYINPUT124), .B(G176gat), .Z(new_n946_));
  XNOR2_X1  g745(.A(new_n945_), .B(new_n946_), .ZN(G1349gat));
  NOR2_X1   g746(.A1(new_n944_), .A2(new_n357_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n948_), .A2(new_n381_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n949_), .B1(new_n385_), .B2(new_n948_), .ZN(G1350gat));
  INV_X1    g749(.A(new_n944_), .ZN(new_n951_));
  OAI211_X1 g750(.A(new_n951_), .B(new_n639_), .C1(new_n428_), .C2(new_n429_), .ZN(new_n952_));
  INV_X1    g751(.A(KEYINPUT125), .ZN(new_n953_));
  NAND4_X1  g752(.A1(new_n910_), .A2(new_n526_), .A3(new_n295_), .A4(new_n933_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n953_), .B1(new_n954_), .B2(G190gat), .ZN(new_n955_));
  OAI211_X1 g754(.A(new_n953_), .B(G190gat), .C1(new_n944_), .C2(new_n691_), .ZN(new_n956_));
  INV_X1    g755(.A(new_n956_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n952_), .B1(new_n955_), .B2(new_n957_), .ZN(new_n958_));
  INV_X1    g757(.A(KEYINPUT126), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n958_), .A2(new_n959_), .ZN(new_n960_));
  OAI211_X1 g759(.A(KEYINPUT126), .B(new_n952_), .C1(new_n955_), .C2(new_n957_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n960_), .A2(new_n961_), .ZN(G1351gat));
  INV_X1    g761(.A(new_n586_), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n911_), .A2(new_n963_), .A3(new_n718_), .ZN(new_n964_));
  INV_X1    g763(.A(new_n964_), .ZN(new_n965_));
  AOI21_X1  g764(.A(G197gat), .B1(new_n965_), .B2(new_n625_), .ZN(new_n966_));
  NOR3_X1   g765(.A1(new_n964_), .A2(new_n395_), .A3(new_n626_), .ZN(new_n967_));
  NOR2_X1   g766(.A1(new_n966_), .A2(new_n967_), .ZN(G1352gat));
  AOI21_X1  g767(.A(G204gat), .B1(new_n965_), .B2(new_n324_), .ZN(new_n969_));
  NOR3_X1   g768(.A1(new_n964_), .A2(new_n397_), .A3(new_n749_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(new_n969_), .A2(new_n970_), .ZN(G1353gat));
  XNOR2_X1  g770(.A(KEYINPUT63), .B(G211gat), .ZN(new_n972_));
  NOR3_X1   g771(.A1(new_n964_), .A2(new_n357_), .A3(new_n972_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n965_), .A2(new_n636_), .ZN(new_n974_));
  NOR2_X1   g773(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n975_));
  AOI21_X1  g774(.A(new_n973_), .B1(new_n974_), .B2(new_n975_), .ZN(G1354gat));
  INV_X1    g775(.A(G218gat), .ZN(new_n977_));
  NOR3_X1   g776(.A1(new_n964_), .A2(new_n977_), .A3(new_n691_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n965_), .A2(new_n639_), .ZN(new_n979_));
  AOI21_X1  g778(.A(new_n978_), .B1(new_n977_), .B2(new_n979_), .ZN(G1355gat));
endmodule


