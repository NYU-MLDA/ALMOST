//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 1 0 0 1 0 0 1 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n670_, new_n671_,
    new_n672_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n774_, new_n775_, new_n777_, new_n778_, new_n779_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT0), .B(G57gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G113gat), .B(G120gat), .ZN(new_n206_));
  INV_X1    g005(.A(G134gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(G127gat), .ZN(new_n208_));
  INV_X1    g007(.A(G127gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G134gat), .ZN(new_n210_));
  AND3_X1   g009(.A1(new_n208_), .A2(new_n210_), .A3(KEYINPUT87), .ZN(new_n211_));
  AOI21_X1  g010(.A(KEYINPUT87), .B1(new_n208_), .B2(new_n210_), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n206_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT87), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n209_), .A2(G134gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n207_), .A2(G127gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n208_), .A2(new_n210_), .A3(KEYINPUT87), .ZN(new_n218_));
  XOR2_X1   g017(.A(G113gat), .B(G120gat), .Z(new_n219_));
  NAND3_X1  g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n213_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n222_));
  INV_X1    g021(.A(G141gat), .ZN(new_n223_));
  INV_X1    g022(.A(G148gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G141gat), .A2(G148gat), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT2), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n225_), .A2(new_n228_), .A3(new_n229_), .A4(new_n230_), .ZN(new_n231_));
  OR2_X1    g030(.A1(G155gat), .A2(G162gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G155gat), .A2(G162gat), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(KEYINPUT1), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT1), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n236_), .A2(G155gat), .A3(G162gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n237_), .A3(new_n232_), .ZN(new_n238_));
  XOR2_X1   g037(.A(G141gat), .B(G148gat), .Z(new_n239_));
  AOI22_X1  g038(.A1(new_n231_), .A2(new_n234_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n221_), .A2(KEYINPUT101), .A3(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(KEYINPUT101), .B1(new_n221_), .B2(new_n240_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT100), .ZN(new_n245_));
  AOI21_X1  g044(.A(KEYINPUT88), .B1(new_n213_), .B2(new_n220_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT88), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n211_), .A2(new_n212_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n247_), .B1(new_n248_), .B2(new_n219_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n231_), .A2(new_n234_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n238_), .A2(new_n239_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n245_), .B1(new_n250_), .B2(new_n253_), .ZN(new_n254_));
  NOR4_X1   g053(.A1(new_n246_), .A2(new_n249_), .A3(KEYINPUT100), .A4(new_n240_), .ZN(new_n255_));
  OAI211_X1 g054(.A(KEYINPUT4), .B(new_n244_), .C1(new_n254_), .C2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n221_), .A2(new_n247_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n248_), .A2(new_n219_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT88), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n257_), .A2(new_n253_), .A3(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n260_), .A2(KEYINPUT4), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G225gat), .A2(G233gat), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n256_), .A2(KEYINPUT102), .A3(new_n263_), .ZN(new_n264_));
  OAI211_X1 g063(.A(new_n244_), .B(new_n262_), .C1(new_n254_), .C2(new_n255_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT102), .B1(new_n256_), .B2(new_n263_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n205_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n256_), .A2(new_n263_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT102), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n205_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n271_), .A2(new_n272_), .A3(new_n265_), .A4(new_n264_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n268_), .A2(KEYINPUT104), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT104), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n275_), .B(new_n205_), .C1(new_n266_), .C2(new_n267_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(KEYINPUT92), .B(KEYINPUT21), .Z(new_n278_));
  INV_X1    g077(.A(G197gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT91), .B1(new_n279_), .B2(G204gat), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT91), .ZN(new_n281_));
  INV_X1    g080(.A(G204gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n281_), .A2(new_n282_), .A3(G197gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n279_), .A2(G204gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n278_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT90), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n287_), .B1(new_n282_), .B2(G197gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n279_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n282_), .A2(G197gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT21), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G211gat), .B(G218gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n286_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n284_), .A2(new_n285_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n293_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n295_), .A2(KEYINPUT21), .A3(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n294_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT25), .B(G183gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT26), .B(G190gat), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303_));
  AOI22_X1  g102(.A1(new_n299_), .A2(new_n300_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  OR3_X1    g103(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT82), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT23), .ZN(new_n307_));
  AND3_X1   g106(.A1(KEYINPUT81), .A2(G183gat), .A3(G190gat), .ZN(new_n308_));
  AOI21_X1  g107(.A(KEYINPUT81), .B1(G183gat), .B2(G190gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n307_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT23), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n306_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT81), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n311_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(KEYINPUT81), .A2(G183gat), .A3(G190gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(KEYINPUT82), .B1(new_n317_), .B2(new_n307_), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n304_), .B(new_n305_), .C1(new_n313_), .C2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT84), .ZN(new_n320_));
  INV_X1    g119(.A(G183gat), .ZN(new_n321_));
  INV_X1    g120(.A(G190gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n315_), .A2(KEYINPUT83), .A3(KEYINPUT23), .A4(new_n316_), .ZN(new_n324_));
  NOR3_X1   g123(.A1(new_n308_), .A2(new_n309_), .A3(new_n307_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n307_), .A2(G183gat), .A3(G190gat), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT83), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n323_), .B(new_n324_), .C1(new_n325_), .C2(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(G169gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n319_), .A2(new_n320_), .A3(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n320_), .B1(new_n319_), .B2(new_n332_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n298_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n324_), .B(new_n305_), .C1(new_n325_), .C2(new_n328_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT97), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n327_), .B(new_n326_), .C1(new_n317_), .C2(new_n307_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT97), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n338_), .A2(new_n339_), .A3(new_n324_), .A4(new_n305_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n337_), .A2(new_n340_), .A3(new_n304_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n298_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n323_), .B1(new_n313_), .B2(new_n318_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(new_n331_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n341_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n335_), .A2(KEYINPUT20), .A3(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G226gat), .A2(G233gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n346_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n304_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n351_), .B1(new_n336_), .B2(KEYINPUT97), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n352_), .A2(new_n340_), .B1(new_n343_), .B2(new_n331_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT20), .B1(new_n353_), .B2(new_n342_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n333_), .A2(new_n334_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n342_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n349_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n355_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n350_), .A2(new_n359_), .ZN(new_n360_));
  XOR2_X1   g159(.A(G8gat), .B(G36gat), .Z(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G64gat), .B(G92gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT105), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n360_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT98), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n349_), .B1(new_n345_), .B2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n353_), .A2(KEYINPUT98), .A3(new_n342_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n369_), .A2(KEYINPUT20), .A3(new_n335_), .A4(new_n370_), .ZN(new_n371_));
  NOR3_X1   g170(.A1(new_n333_), .A2(new_n334_), .A3(new_n298_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n349_), .B1(new_n372_), .B2(new_n354_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n371_), .A2(new_n373_), .A3(new_n365_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n367_), .A2(KEYINPUT27), .A3(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G78gat), .B(G106gat), .ZN(new_n376_));
  AOI22_X1  g175(.A1(new_n294_), .A2(new_n297_), .B1(new_n253_), .B2(KEYINPUT29), .ZN(new_n377_));
  AOI21_X1  g176(.A(KEYINPUT93), .B1(new_n294_), .B2(new_n297_), .ZN(new_n378_));
  INV_X1    g177(.A(G233gat), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n379_), .A2(KEYINPUT89), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n379_), .A2(KEYINPUT89), .ZN(new_n381_));
  OAI21_X1  g180(.A(G228gat), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NOR3_X1   g181(.A1(new_n377_), .A2(new_n378_), .A3(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n253_), .A2(KEYINPUT29), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT93), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n298_), .B(new_n384_), .C1(new_n385_), .C2(new_n382_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n376_), .B1(new_n383_), .B2(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n378_), .A2(new_n382_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n377_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n376_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(new_n386_), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT94), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n388_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G22gat), .B(G50gat), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT28), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT29), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n240_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n398_), .B1(new_n240_), .B2(new_n399_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n397_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n402_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n404_), .A2(new_n400_), .A3(new_n396_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n391_), .A2(KEYINPUT94), .A3(new_n386_), .A4(new_n392_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n395_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n406_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n388_), .A2(new_n393_), .A3(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT95), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT95), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n388_), .A2(new_n393_), .A3(new_n409_), .A4(new_n412_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n408_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT27), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n371_), .A2(new_n373_), .A3(new_n365_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n365_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n415_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n375_), .A2(new_n414_), .A3(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT106), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G227gat), .A2(G233gat), .ZN(new_n421_));
  INV_X1    g220(.A(G15gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(G71gat), .ZN(new_n424_));
  INV_X1    g223(.A(G99gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT30), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n356_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n427_), .A2(new_n356_), .ZN(new_n430_));
  NOR3_X1   g229(.A1(new_n429_), .A2(new_n430_), .A3(new_n250_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(KEYINPUT85), .B(G43gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT86), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(KEYINPUT31), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n250_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n432_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n435_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n250_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n430_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n439_), .B1(new_n440_), .B2(new_n428_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n438_), .B1(new_n441_), .B2(new_n431_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n437_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT106), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n375_), .A2(new_n414_), .A3(new_n418_), .A4(new_n444_), .ZN(new_n445_));
  AND4_X1   g244(.A1(new_n277_), .A2(new_n420_), .A3(new_n443_), .A4(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n365_), .A2(KEYINPUT32), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n447_), .B1(new_n350_), .B2(new_n359_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n371_), .A2(new_n373_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n448_), .B1(new_n447_), .B2(new_n450_), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n274_), .A2(new_n276_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n262_), .ZN(new_n453_));
  OAI211_X1 g252(.A(new_n244_), .B(new_n453_), .C1(new_n254_), .C2(new_n255_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(new_n205_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT103), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT103), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n454_), .A2(new_n457_), .A3(new_n205_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n256_), .B(new_n262_), .C1(KEYINPUT4), .C2(new_n260_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n456_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n365_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n449_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n460_), .A2(new_n374_), .A3(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n273_), .A2(KEYINPUT33), .ZN(new_n464_));
  INV_X1    g263(.A(new_n266_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT33), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n465_), .A2(new_n466_), .A3(new_n272_), .A4(new_n271_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n463_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n414_), .B1(new_n452_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n462_), .A2(new_n374_), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n374_), .A2(KEYINPUT27), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n415_), .A2(new_n470_), .B1(new_n471_), .B2(new_n367_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n414_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n277_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n469_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n443_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n446_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G229gat), .A2(G233gat), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G29gat), .B(G36gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G43gat), .B(G50gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n482_), .A2(new_n483_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G1gat), .A2(G8gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT14), .ZN(new_n488_));
  INV_X1    g287(.A(G22gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n422_), .A2(new_n489_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(G15gat), .A2(G22gat), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n488_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n492_), .A2(KEYINPUT75), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(G1gat), .B(G8gat), .Z(new_n495_));
  NAND2_X1  g294(.A1(new_n492_), .A2(KEYINPUT75), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n495_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n486_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n482_), .B(new_n483_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n499_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n501_), .A2(new_n502_), .A3(new_n497_), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n500_), .A2(new_n503_), .A3(KEYINPUT77), .ZN(new_n504_));
  AOI21_X1  g303(.A(KEYINPUT77), .B1(new_n500_), .B2(new_n503_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n479_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n501_), .B(KEYINPUT15), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n502_), .A2(new_n497_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n509_), .A2(new_n503_), .A3(new_n478_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n506_), .A2(new_n510_), .A3(KEYINPUT78), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(KEYINPUT78), .B1(new_n506_), .B2(new_n510_), .ZN(new_n513_));
  XOR2_X1   g312(.A(G113gat), .B(G141gat), .Z(new_n514_));
  XNOR2_X1  g313(.A(G169gat), .B(G197gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT79), .ZN(new_n517_));
  OR3_X1    g316(.A1(new_n512_), .A2(new_n513_), .A3(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n506_), .A2(new_n510_), .A3(new_n516_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT80), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT80), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n506_), .A2(new_n510_), .A3(new_n521_), .A4(new_n516_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n518_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n477_), .A2(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(G120gat), .B(G148gat), .Z(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G176gat), .B(G204gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G230gat), .A2(G233gat), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n533_), .B(KEYINPUT64), .Z(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G99gat), .A2(G106gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(G85gat), .ZN(new_n539_));
  INV_X1    g338(.A(G92gat), .ZN(new_n540_));
  NOR3_X1   g339(.A1(new_n539_), .A2(new_n540_), .A3(KEYINPUT9), .ZN(new_n541_));
  XOR2_X1   g340(.A(G85gat), .B(G92gat), .Z(new_n542_));
  AOI21_X1  g341(.A(new_n541_), .B1(new_n542_), .B2(KEYINPUT9), .ZN(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT10), .B(G99gat), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n538_), .B(new_n543_), .C1(G106gat), .C2(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(G99gat), .A2(G106gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT7), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n538_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT8), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n548_), .A2(new_n549_), .A3(new_n542_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n549_), .B1(new_n548_), .B2(new_n542_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n545_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G57gat), .B(G64gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G71gat), .B(G78gat), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n553_), .A2(new_n554_), .A3(KEYINPUT11), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n553_), .A2(KEYINPUT11), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n556_), .A2(new_n554_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n553_), .A2(KEYINPUT11), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n555_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n552_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n548_), .A2(new_n542_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT8), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n548_), .A2(new_n549_), .A3(new_n542_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n559_), .B1(new_n565_), .B2(new_n545_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n535_), .B1(new_n561_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT66), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  OAI211_X1 g368(.A(KEYINPUT66), .B(new_n535_), .C1(new_n561_), .C2(new_n566_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n552_), .A2(new_n560_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n565_), .A2(new_n559_), .A3(new_n545_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n572_), .A2(new_n573_), .A3(KEYINPUT12), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT12), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n566_), .A2(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n535_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n532_), .B1(new_n571_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT68), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n574_), .A2(new_n576_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(new_n534_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n581_), .A2(new_n569_), .A3(new_n570_), .A4(new_n531_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n578_), .A2(new_n579_), .A3(new_n582_), .ZN(new_n583_));
  OAI211_X1 g382(.A(KEYINPUT68), .B(new_n532_), .C1(new_n571_), .C2(new_n577_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT13), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT69), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n586_), .A2(KEYINPUT69), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n585_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n583_), .A2(KEYINPUT69), .A3(new_n586_), .A4(new_n584_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n507_), .A2(new_n552_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G232gat), .A2(G233gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  XOR2_X1   g395(.A(KEYINPUT71), .B(KEYINPUT35), .Z(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  OAI211_X1 g397(.A(new_n593_), .B(new_n598_), .C1(new_n486_), .C2(new_n552_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n596_), .A2(new_n597_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G190gat), .B(G218gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G134gat), .B(G162gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT36), .Z(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT74), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n601_), .A2(new_n606_), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n604_), .A2(KEYINPUT36), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n601_), .A2(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(KEYINPUT37), .B1(new_n607_), .B2(new_n609_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n601_), .A2(new_n608_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT37), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n601_), .A2(new_n605_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n611_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n610_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT76), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n508_), .B(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(new_n560_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT17), .ZN(new_n621_));
  XOR2_X1   g420(.A(G127gat), .B(G155gat), .Z(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT16), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G183gat), .B(G211gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  OR3_X1    g424(.A1(new_n620_), .A2(new_n621_), .A3(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(KEYINPUT17), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n620_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n615_), .A2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n592_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n526_), .A2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n277_), .B(KEYINPUT107), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  OR3_X1    g434(.A1(new_n633_), .A2(G1gat), .A3(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(KEYINPUT108), .B(KEYINPUT38), .ZN(new_n637_));
  OR2_X1    g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n637_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n591_), .A2(new_n524_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n611_), .A2(new_n613_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NOR4_X1   g441(.A1(new_n640_), .A2(new_n477_), .A3(new_n629_), .A4(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G1gat), .B1(new_n644_), .B2(new_n277_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n638_), .A2(new_n639_), .A3(new_n645_), .ZN(G1324gat));
  INV_X1    g445(.A(KEYINPUT109), .ZN(new_n647_));
  INV_X1    g446(.A(G8gat), .ZN(new_n648_));
  INV_X1    g447(.A(new_n472_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n643_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n647_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n650_), .A2(KEYINPUT110), .A3(new_n651_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n640_), .A2(new_n629_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n477_), .A2(new_n642_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n655_), .A3(new_n649_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(G8gat), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(KEYINPUT109), .A3(KEYINPUT39), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT110), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n659_), .B1(new_n657_), .B2(KEYINPUT39), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n652_), .A2(new_n653_), .A3(new_n658_), .A4(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n633_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n662_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(KEYINPUT111), .B(KEYINPUT40), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n661_), .A2(new_n663_), .A3(new_n665_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1325gat));
  AOI21_X1  g468(.A(new_n422_), .B1(new_n643_), .B2(new_n443_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT41), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n662_), .A2(new_n422_), .A3(new_n443_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1326gat));
  AOI21_X1  g472(.A(new_n489_), .B1(new_n643_), .B2(new_n473_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT42), .Z(new_n675_));
  NAND3_X1  g474(.A1(new_n662_), .A2(new_n489_), .A3(new_n473_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1327gat));
  NOR2_X1   g476(.A1(new_n630_), .A2(new_n641_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n592_), .A2(new_n679_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n526_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n277_), .ZN(new_n682_));
  AOI21_X1  g481(.A(G29gat), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT112), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n591_), .A2(new_n524_), .A3(new_n629_), .ZN(new_n685_));
  OAI21_X1  g484(.A(KEYINPUT43), .B1(new_n477_), .B2(new_n615_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n467_), .A2(new_n464_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n463_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n274_), .A2(new_n276_), .A3(new_n451_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n473_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  AND3_X1   g490(.A1(new_n277_), .A2(new_n473_), .A3(new_n472_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n476_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n420_), .A2(new_n443_), .A3(new_n277_), .A4(new_n445_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT43), .ZN(new_n696_));
  INV_X1    g495(.A(new_n615_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n695_), .A2(new_n696_), .A3(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n685_), .B1(new_n686_), .B2(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n684_), .B1(new_n699_), .B2(KEYINPUT44), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n696_), .B1(new_n695_), .B2(new_n697_), .ZN(new_n702_));
  AOI211_X1 g501(.A(KEYINPUT43), .B(new_n615_), .C1(new_n693_), .C2(new_n694_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  OAI211_X1 g503(.A(KEYINPUT112), .B(new_n701_), .C1(new_n704_), .C2(new_n685_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n685_), .ZN(new_n706_));
  OAI211_X1 g505(.A(KEYINPUT44), .B(new_n706_), .C1(new_n702_), .C2(new_n703_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT113), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n686_), .A2(new_n698_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT113), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n709_), .A2(new_n710_), .A3(KEYINPUT44), .A4(new_n706_), .ZN(new_n711_));
  AOI22_X1  g510(.A1(new_n700_), .A2(new_n705_), .B1(new_n708_), .B2(new_n711_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n634_), .A2(G29gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n683_), .B1(new_n712_), .B2(new_n713_), .ZN(G1328gat));
  INV_X1    g513(.A(KEYINPUT46), .ZN(new_n715_));
  INV_X1    g514(.A(G36gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n712_), .B2(new_n649_), .ZN(new_n717_));
  XOR2_X1   g516(.A(KEYINPUT114), .B(KEYINPUT45), .Z(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n472_), .A2(G36gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT115), .B1(new_n681_), .B2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n526_), .A2(new_n680_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT115), .ZN(new_n723_));
  INV_X1    g522(.A(new_n720_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n722_), .A2(new_n723_), .A3(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n719_), .B1(new_n721_), .B2(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n681_), .A2(KEYINPUT115), .A3(new_n720_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n723_), .B1(new_n722_), .B2(new_n724_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n727_), .A2(new_n718_), .A3(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n726_), .A2(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n715_), .B1(new_n717_), .B2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n700_), .A2(new_n705_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n708_), .A2(new_n711_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(new_n649_), .A3(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(G36gat), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n726_), .A2(new_n729_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(KEYINPUT46), .A3(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n731_), .A2(new_n737_), .ZN(G1329gat));
  NAND4_X1  g537(.A1(new_n732_), .A2(G43gat), .A3(new_n443_), .A4(new_n733_), .ZN(new_n739_));
  XOR2_X1   g538(.A(KEYINPUT116), .B(G43gat), .Z(new_n740_));
  OAI21_X1  g539(.A(new_n740_), .B1(new_n722_), .B2(new_n476_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT47), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT47), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n739_), .A2(new_n744_), .A3(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1330gat));
  AOI21_X1  g545(.A(G50gat), .B1(new_n681_), .B2(new_n473_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n473_), .A2(G50gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n712_), .B2(new_n748_), .ZN(G1331gat));
  NAND4_X1  g548(.A1(new_n655_), .A2(new_n525_), .A3(new_n592_), .A4(new_n630_), .ZN(new_n750_));
  OAI21_X1  g549(.A(G57gat), .B1(new_n750_), .B2(new_n277_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n477_), .A2(new_n524_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n752_), .A2(new_n592_), .A3(new_n630_), .A4(new_n615_), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n635_), .A2(G57gat), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n751_), .B1(new_n753_), .B2(new_n754_), .ZN(G1332gat));
  OAI21_X1  g554(.A(G64gat), .B1(new_n750_), .B2(new_n472_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT48), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n472_), .A2(G64gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n753_), .B2(new_n758_), .ZN(G1333gat));
  OAI21_X1  g558(.A(G71gat), .B1(new_n750_), .B2(new_n476_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT49), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n476_), .A2(G71gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n761_), .B1(new_n753_), .B2(new_n762_), .ZN(G1334gat));
  OAI21_X1  g562(.A(G78gat), .B1(new_n750_), .B2(new_n414_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT50), .ZN(new_n765_));
  OR2_X1    g564(.A1(new_n414_), .A2(G78gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n753_), .B2(new_n766_), .ZN(G1335gat));
  NOR4_X1   g566(.A1(new_n477_), .A2(new_n591_), .A3(new_n524_), .A4(new_n679_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n768_), .A2(new_n539_), .A3(new_n634_), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n591_), .A2(new_n524_), .A3(new_n630_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n709_), .A2(new_n770_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n771_), .A2(new_n682_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n769_), .B1(new_n772_), .B2(new_n539_), .ZN(G1336gat));
  NAND3_X1  g572(.A1(new_n768_), .A2(new_n540_), .A3(new_n649_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n771_), .A2(new_n649_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(new_n540_), .ZN(G1337gat));
  NAND2_X1  g575(.A1(new_n771_), .A2(new_n443_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n476_), .A2(new_n544_), .ZN(new_n778_));
  AOI22_X1  g577(.A1(new_n777_), .A2(G99gat), .B1(new_n768_), .B2(new_n778_), .ZN(new_n779_));
  XOR2_X1   g578(.A(new_n779_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g579(.A1(new_n709_), .A2(new_n473_), .A3(new_n770_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(G106gat), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT117), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n781_), .A2(KEYINPUT117), .A3(G106gat), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n784_), .A2(KEYINPUT52), .A3(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT117), .B1(new_n781_), .B2(G106gat), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n414_), .A2(G106gat), .ZN(new_n789_));
  AOI22_X1  g588(.A1(new_n787_), .A2(new_n788_), .B1(new_n768_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n786_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT53), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n786_), .A2(new_n790_), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(G1339gat));
  AND3_X1   g594(.A1(new_n420_), .A2(new_n443_), .A3(new_n445_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n478_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n503_), .A2(new_n479_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n516_), .B1(new_n509_), .B2(new_n798_), .ZN(new_n799_));
  AOI22_X1  g598(.A1(new_n520_), .A2(new_n522_), .B1(new_n797_), .B2(new_n799_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n583_), .A2(new_n800_), .A3(new_n584_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n574_), .A2(new_n576_), .A3(new_n535_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT55), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n581_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n580_), .A2(KEYINPUT55), .A3(new_n534_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n531_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(KEYINPUT118), .B1(new_n806_), .B2(KEYINPUT56), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(KEYINPUT56), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n577_), .B1(KEYINPUT55), .B2(new_n802_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n805_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n532_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT56), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n811_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n807_), .A2(new_n808_), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n582_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n816_), .B1(new_n518_), .B2(new_n523_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n801_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(KEYINPUT119), .B1(new_n818_), .B2(new_n642_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n811_), .A2(KEYINPUT120), .A3(new_n813_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n800_), .A2(new_n582_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT120), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n808_), .A2(new_n822_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n806_), .A2(KEYINPUT56), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n820_), .B(new_n821_), .C1(new_n823_), .C2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT58), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n615_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n821_), .A2(new_n820_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n828_), .B(KEYINPUT58), .C1(new_n824_), .C2(new_n823_), .ZN(new_n829_));
  AOI22_X1  g628(.A1(new_n819_), .A2(KEYINPUT57), .B1(new_n827_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n831_));
  OAI211_X1 g630(.A(KEYINPUT119), .B(new_n831_), .C1(new_n818_), .C2(new_n642_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n630_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n591_), .A2(new_n525_), .A3(new_n630_), .A4(new_n615_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n834_), .B(new_n835_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n796_), .B(new_n634_), .C1(new_n833_), .C2(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(KEYINPUT121), .B2(KEYINPUT59), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n819_), .A2(KEYINPUT57), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n827_), .A2(new_n829_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n832_), .A3(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n629_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n834_), .B(KEYINPUT54), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n635_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  XOR2_X1   g643(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n844_), .A2(new_n796_), .A3(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n838_), .A2(new_n847_), .A3(new_n524_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(G113gat), .ZN(new_n849_));
  OR3_X1    g648(.A1(new_n837_), .A2(G113gat), .A3(new_n525_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1340gat));
  XOR2_X1   g650(.A(KEYINPUT122), .B(G120gat), .Z(new_n852_));
  OR2_X1    g651(.A1(new_n852_), .A2(KEYINPUT60), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n591_), .B2(KEYINPUT60), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n844_), .A2(new_n796_), .A3(new_n853_), .A4(new_n854_), .ZN(new_n855_));
  AND3_X1   g654(.A1(new_n838_), .A2(new_n592_), .A3(new_n847_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(new_n852_), .ZN(G1341gat));
  OAI21_X1  g656(.A(G127gat), .B1(new_n629_), .B2(KEYINPUT123), .ZN(new_n858_));
  OR2_X1    g657(.A1(KEYINPUT123), .A2(G127gat), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n838_), .A2(new_n847_), .A3(new_n858_), .A4(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n209_), .B1(new_n837_), .B2(new_n629_), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1342gat));
  XNOR2_X1  g661(.A(KEYINPUT124), .B(G134gat), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n838_), .A2(new_n847_), .A3(new_n697_), .A4(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n207_), .B1(new_n837_), .B2(new_n641_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n864_), .A2(new_n865_), .ZN(G1343gat));
  NOR3_X1   g665(.A1(new_n443_), .A2(new_n649_), .A3(new_n414_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n844_), .A2(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n525_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(new_n223_), .ZN(G1344gat));
  NOR2_X1   g669(.A1(new_n868_), .A2(new_n591_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(new_n224_), .ZN(G1345gat));
  XNOR2_X1  g671(.A(KEYINPUT61), .B(G155gat), .ZN(new_n873_));
  OR3_X1    g672(.A1(new_n868_), .A2(new_n629_), .A3(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n868_), .B2(new_n629_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(G1346gat));
  OR3_X1    g675(.A1(new_n868_), .A2(G162gat), .A3(new_n641_), .ZN(new_n877_));
  OAI21_X1  g676(.A(G162gat), .B1(new_n868_), .B2(new_n615_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(G1347gat));
  AOI21_X1  g678(.A(new_n472_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n634_), .A2(new_n473_), .A3(new_n476_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(G169gat), .B1(new_n882_), .B2(new_n525_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT125), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(KEYINPUT62), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n887_));
  OAI211_X1 g686(.A(G169gat), .B(new_n887_), .C1(new_n882_), .C2(new_n525_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT22), .B(G169gat), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n880_), .A2(new_n524_), .A3(new_n881_), .A4(new_n889_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n886_), .A2(new_n888_), .A3(new_n890_), .ZN(G1348gat));
  NAND3_X1  g690(.A1(new_n880_), .A2(new_n592_), .A3(new_n881_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g692(.A1(new_n880_), .A2(new_n630_), .A3(new_n881_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n894_), .A2(new_n299_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n895_), .B1(new_n321_), .B2(new_n894_), .ZN(G1350gat));
  OAI21_X1  g695(.A(G190gat), .B1(new_n882_), .B2(new_n615_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n642_), .A2(new_n300_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n882_), .B2(new_n898_), .ZN(G1351gat));
  NOR3_X1   g698(.A1(new_n682_), .A2(new_n443_), .A3(new_n414_), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n649_), .B(new_n900_), .C1(new_n833_), .C2(new_n836_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n901_), .A2(new_n525_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(new_n279_), .ZN(G1352gat));
  NOR2_X1   g702(.A1(new_n901_), .A2(new_n591_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n282_), .A2(KEYINPUT126), .ZN(new_n905_));
  XOR2_X1   g704(.A(new_n904_), .B(new_n905_), .Z(G1353gat));
  AOI21_X1  g705(.A(new_n629_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  OAI21_X1  g707(.A(KEYINPUT127), .B1(new_n901_), .B2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT127), .ZN(new_n910_));
  NAND4_X1  g709(.A1(new_n880_), .A2(new_n910_), .A3(new_n900_), .A4(new_n907_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  AND3_X1   g711(.A1(new_n909_), .A2(new_n911_), .A3(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n912_), .B1(new_n909_), .B2(new_n911_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1354gat));
  OAI21_X1  g714(.A(G218gat), .B1(new_n901_), .B2(new_n615_), .ZN(new_n916_));
  OR2_X1    g715(.A1(new_n641_), .A2(G218gat), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n901_), .B2(new_n917_), .ZN(G1355gat));
endmodule


