//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 0 0 1 1 1 1 1 1 0 1 1 0 0 1 1 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n845_, new_n846_, new_n848_, new_n849_, new_n850_, new_n852_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_;
  NAND2_X1  g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT2), .ZN(new_n203_));
  OR4_X1    g002(.A1(KEYINPUT87), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n204_));
  INV_X1    g003(.A(G141gat), .ZN(new_n205_));
  INV_X1    g004(.A(G148gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT3), .B1(new_n207_), .B2(KEYINPUT87), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n203_), .A2(new_n204_), .A3(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT86), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n209_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(KEYINPUT1), .ZN(new_n215_));
  OAI211_X1 g014(.A(new_n207_), .B(new_n202_), .C1(new_n211_), .C2(new_n215_), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT94), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G113gat), .B(G120gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT83), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  OR2_X1    g020(.A1(G113gat), .A2(G120gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G113gat), .A2(G120gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(KEYINPUT83), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n221_), .A2(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(G127gat), .B(G134gat), .Z(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n221_), .A2(new_n224_), .A3(new_n226_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n217_), .A2(new_n218_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n214_), .A2(new_n216_), .ZN(new_n232_));
  AND3_X1   g031(.A1(new_n221_), .A2(new_n224_), .A3(new_n226_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n226_), .B1(new_n221_), .B2(new_n224_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT94), .B1(new_n232_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n231_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT93), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT84), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n229_), .A2(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n240_), .B1(new_n235_), .B2(new_n239_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n238_), .B1(new_n241_), .B2(new_n217_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n240_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n243_), .B1(new_n230_), .B2(KEYINPUT84), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n244_), .A2(KEYINPUT93), .A3(new_n232_), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n237_), .A2(new_n242_), .A3(KEYINPUT4), .A4(new_n245_), .ZN(new_n246_));
  XOR2_X1   g045(.A(KEYINPUT96), .B(KEYINPUT4), .Z(new_n247_));
  NAND3_X1  g046(.A1(new_n244_), .A2(new_n232_), .A3(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G225gat), .A2(G233gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT95), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n246_), .A2(new_n248_), .A3(new_n250_), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n237_), .A2(new_n242_), .A3(new_n249_), .A4(new_n245_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT0), .B(G57gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(G85gat), .ZN(new_n255_));
  XOR2_X1   g054(.A(G1gat), .B(G29gat), .Z(new_n256_));
  XOR2_X1   g055(.A(new_n255_), .B(new_n256_), .Z(new_n257_));
  NAND2_X1  g056(.A1(new_n253_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n257_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n251_), .A2(new_n252_), .A3(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n258_), .A2(KEYINPUT101), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT101), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n251_), .A2(new_n262_), .A3(new_n252_), .A4(new_n259_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT103), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G230gat), .A2(G233gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G99gat), .A2(G106gat), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT6), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT64), .ZN(new_n274_));
  INV_X1    g073(.A(G99gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT10), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT10), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(G99gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(G106gat), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n274_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  AOI211_X1 g080(.A(KEYINPUT64), .B(G106gat), .C1(new_n276_), .C2(new_n278_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n273_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT65), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT9), .ZN(new_n285_));
  INV_X1    g084(.A(G85gat), .ZN(new_n286_));
  INV_X1    g085(.A(G92gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G85gat), .A2(G92gat), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n285_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n285_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n284_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n293_));
  AND2_X1   g092(.A1(G85gat), .A2(G92gat), .ZN(new_n294_));
  NOR2_X1   g093(.A1(G85gat), .A2(G92gat), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  OAI211_X1 g095(.A(KEYINPUT65), .B(new_n291_), .C1(new_n296_), .C2(new_n285_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n293_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT7), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n299_), .A2(new_n275_), .A3(new_n280_), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n300_), .A2(new_n271_), .A3(new_n272_), .A4(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT8), .ZN(new_n303_));
  AND3_X1   g102(.A1(new_n302_), .A2(new_n303_), .A3(new_n296_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n303_), .B1(new_n302_), .B2(new_n296_), .ZN(new_n305_));
  OAI22_X1  g104(.A1(new_n283_), .A2(new_n298_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT66), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n305_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n302_), .A2(new_n303_), .A3(new_n296_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT10), .B(G99gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT64), .B1(new_n312_), .B2(G106gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n279_), .A2(new_n274_), .A3(new_n280_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND4_X1  g114(.A1(new_n315_), .A2(new_n273_), .A3(new_n293_), .A4(new_n297_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n311_), .A2(new_n316_), .A3(KEYINPUT66), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G57gat), .B(G64gat), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n318_), .A2(KEYINPUT11), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(KEYINPUT11), .ZN(new_n320_));
  XOR2_X1   g119(.A(G71gat), .B(G78gat), .Z(new_n321_));
  NAND3_X1  g120(.A1(new_n319_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n320_), .A2(new_n321_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n308_), .A2(new_n317_), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT68), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n308_), .A2(KEYINPUT68), .A3(new_n317_), .A4(new_n325_), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT67), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n308_), .A2(new_n317_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n331_), .B1(new_n332_), .B2(new_n324_), .ZN(new_n333_));
  AOI211_X1 g132(.A(KEYINPUT67), .B(new_n325_), .C1(new_n308_), .C2(new_n317_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n268_), .B1(new_n330_), .B2(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n325_), .B1(new_n308_), .B2(new_n317_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT12), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n337_), .B1(new_n338_), .B2(new_n326_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n306_), .A2(new_n325_), .A3(KEYINPUT12), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n339_), .A2(new_n268_), .A3(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n267_), .B1(new_n336_), .B2(new_n341_), .ZN(new_n342_));
  XOR2_X1   g141(.A(G120gat), .B(G148gat), .Z(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(G204gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT5), .ZN(new_n345_));
  INV_X1    g144(.A(G176gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n317_), .ZN(new_n349_));
  AOI21_X1  g148(.A(KEYINPUT66), .B1(new_n311_), .B2(new_n316_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n324_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(KEYINPUT67), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n337_), .A2(new_n331_), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n352_), .A2(new_n353_), .A3(new_n328_), .A4(new_n329_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n268_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n339_), .A2(new_n268_), .A3(new_n340_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n356_), .A2(new_n357_), .A3(KEYINPUT69), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n342_), .A2(new_n348_), .A3(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT70), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n356_), .A2(new_n357_), .A3(new_n347_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT70), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n342_), .A2(new_n362_), .A3(new_n358_), .A4(new_n348_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n360_), .A2(new_n361_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT13), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT13), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n360_), .A2(new_n366_), .A3(new_n361_), .A4(new_n363_), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n365_), .A2(KEYINPUT71), .A3(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(KEYINPUT71), .B1(new_n365_), .B2(new_n367_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT78), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G15gat), .B(G22gat), .ZN(new_n371_));
  INV_X1    g170(.A(G1gat), .ZN(new_n372_));
  INV_X1    g171(.A(G8gat), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT14), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n371_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G1gat), .B(G8gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(G29gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT72), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT72), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(G29gat), .ZN(new_n381_));
  INV_X1    g180(.A(G36gat), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n379_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n382_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G43gat), .B(G50gat), .ZN(new_n386_));
  NOR3_X1   g185(.A1(new_n384_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n386_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n379_), .A2(new_n381_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(G36gat), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n388_), .B1(new_n390_), .B2(new_n383_), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT73), .B1(new_n387_), .B2(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n386_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n390_), .A2(new_n388_), .A3(new_n383_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT73), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n393_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  AND3_X1   g195(.A1(new_n392_), .A2(KEYINPUT15), .A3(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(KEYINPUT15), .B1(new_n392_), .B2(new_n396_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n377_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n387_), .A2(new_n391_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n399_), .B1(new_n401_), .B2(new_n377_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G229gat), .A2(G233gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  XOR2_X1   g204(.A(new_n400_), .B(new_n377_), .Z(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n404_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n370_), .B1(new_n405_), .B2(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G113gat), .B(G141gat), .ZN(new_n410_));
  INV_X1    g209(.A(G169gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(G197gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  OAI211_X1 g213(.A(KEYINPUT78), .B(new_n407_), .C1(new_n402_), .C2(new_n404_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n409_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT79), .ZN(new_n417_));
  OR3_X1    g216(.A1(new_n405_), .A2(new_n414_), .A3(new_n408_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT79), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n409_), .A2(new_n419_), .A3(new_n414_), .A4(new_n415_), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n417_), .A2(new_n418_), .A3(new_n420_), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n368_), .A2(new_n369_), .A3(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT16), .B(G183gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(G211gat), .ZN(new_n424_));
  XOR2_X1   g223(.A(G127gat), .B(G155gat), .Z(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G231gat), .A2(G233gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n377_), .B(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(new_n325_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n426_), .B1(new_n429_), .B2(KEYINPUT17), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n430_), .B1(KEYINPUT17), .B2(new_n426_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n429_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT77), .ZN(new_n433_));
  XOR2_X1   g232(.A(new_n431_), .B(new_n433_), .Z(new_n434_));
  INV_X1    g233(.A(new_n264_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(KEYINPUT82), .A2(KEYINPUT22), .ZN(new_n436_));
  OAI21_X1  g235(.A(G169gat), .B1(new_n436_), .B2(G176gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT22), .B(G169gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n346_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT82), .ZN(new_n440_));
  XOR2_X1   g239(.A(KEYINPUT80), .B(G183gat), .Z(new_n441_));
  NOR2_X1   g240(.A1(new_n441_), .A2(G190gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G183gat), .A2(G190gat), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT23), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  OAI221_X1 g244(.A(new_n437_), .B1(new_n439_), .B2(new_n440_), .C1(new_n442_), .C2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n411_), .A2(new_n346_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n447_), .A2(KEYINPUT24), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n445_), .A2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n450_), .B1(new_n441_), .B2(KEYINPUT25), .ZN(new_n451_));
  XOR2_X1   g250(.A(KEYINPUT26), .B(G190gat), .Z(new_n452_));
  OAI21_X1  g251(.A(new_n449_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G169gat), .A2(G176gat), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n447_), .A2(KEYINPUT24), .A3(new_n454_), .ZN(new_n455_));
  XOR2_X1   g254(.A(new_n455_), .B(KEYINPUT81), .Z(new_n456_));
  OAI21_X1  g255(.A(new_n446_), .B1(new_n453_), .B2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  AND2_X1   g257(.A1(G211gat), .A2(G218gat), .ZN(new_n459_));
  NOR2_X1   g258(.A1(G211gat), .A2(G218gat), .ZN(new_n460_));
  OAI21_X1  g259(.A(KEYINPUT89), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT21), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G197gat), .B(G204gat), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n461_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n464_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n463_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(new_n461_), .A3(KEYINPUT21), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n465_), .A2(KEYINPUT90), .A3(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(KEYINPUT90), .B1(new_n465_), .B2(new_n467_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n458_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(KEYINPUT25), .B(G183gat), .Z(new_n471_));
  OAI211_X1 g270(.A(new_n449_), .B(new_n455_), .C1(new_n452_), .C2(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(G183gat), .A2(G190gat), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n439_), .B(new_n454_), .C1(new_n445_), .C2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n465_), .A2(new_n467_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n470_), .A2(KEYINPUT20), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G226gat), .A2(G233gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT19), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n478_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT20), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n468_), .A2(new_n469_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n483_), .B1(new_n484_), .B2(new_n457_), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n475_), .A2(new_n476_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n482_), .B1(new_n481_), .B2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G8gat), .B(G36gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G64gat), .B(G92gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT32), .ZN(new_n495_));
  OR2_X1    g294(.A1(new_n488_), .A2(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n480_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n470_), .A2(KEYINPUT20), .A3(new_n480_), .A4(new_n477_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT100), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(new_n501_), .A3(new_n495_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n499_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n495_), .B1(new_n503_), .B2(new_n497_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT100), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n435_), .A2(KEYINPUT102), .A3(new_n496_), .A4(new_n506_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n506_), .A2(new_n261_), .A3(new_n263_), .A4(new_n496_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT102), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  XOR2_X1   g309(.A(KEYINPUT97), .B(KEYINPUT33), .Z(new_n511_));
  NAND2_X1  g310(.A1(new_n260_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT98), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  NOR3_X1   g313(.A1(new_n503_), .A2(new_n497_), .A3(new_n494_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n493_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n260_), .ZN(new_n517_));
  AOI211_X1 g316(.A(new_n515_), .B(new_n516_), .C1(KEYINPUT33), .C2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n246_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n519_), .B(KEYINPUT99), .Z(new_n520_));
  AND3_X1   g319(.A1(new_n237_), .A2(new_n242_), .A3(new_n245_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n259_), .B1(new_n521_), .B2(new_n250_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n514_), .A2(new_n518_), .A3(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n507_), .A2(new_n510_), .A3(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G227gat), .A2(G233gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(G15gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G71gat), .B(G99gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n527_), .B(new_n528_), .Z(new_n529_));
  NAND2_X1  g328(.A1(new_n457_), .A2(KEYINPUT30), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n457_), .A2(KEYINPUT30), .ZN(new_n532_));
  OAI21_X1  g331(.A(G43gat), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n532_), .ZN(new_n534_));
  INV_X1    g333(.A(G43gat), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n535_), .A3(new_n530_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n529_), .B1(new_n533_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n533_), .A2(new_n536_), .A3(new_n529_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n538_), .A2(KEYINPUT85), .A3(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT85), .ZN(new_n541_));
  INV_X1    g340(.A(new_n539_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n541_), .B1(new_n542_), .B2(new_n537_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n241_), .B(KEYINPUT31), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n540_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n544_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n538_), .A2(KEYINPUT85), .A3(new_n539_), .A4(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n232_), .A2(KEYINPUT29), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G22gat), .B(G50gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT28), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n549_), .B(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G228gat), .A2(G233gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n232_), .A2(KEYINPUT29), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n484_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n476_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n557_), .A2(G228gat), .A3(G233gat), .ZN(new_n558_));
  INV_X1    g357(.A(G78gat), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n556_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n559_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n280_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n556_), .A2(new_n558_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(G78gat), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n565_), .A2(G106gat), .A3(new_n560_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT88), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n563_), .A2(new_n566_), .A3(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT91), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT91), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n563_), .A2(new_n566_), .A3(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n553_), .B1(new_n569_), .B2(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n552_), .B1(new_n568_), .B2(KEYINPUT91), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n525_), .A2(new_n548_), .A3(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n516_), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n576_), .B(KEYINPUT27), .C1(new_n494_), .C2(new_n488_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT27), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n578_), .B1(new_n516_), .B2(new_n515_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n545_), .A2(new_n547_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n569_), .A2(new_n571_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(new_n552_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n573_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n581_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n572_), .A2(new_n548_), .A3(new_n573_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n266_), .B(new_n580_), .C1(new_n585_), .C2(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n434_), .B1(new_n575_), .B2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n422_), .A2(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n400_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n306_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT34), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n593_), .A2(KEYINPUT35), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n590_), .A2(new_n591_), .A3(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n590_), .A2(KEYINPUT74), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n596_), .A2(new_n597_), .A3(KEYINPUT35), .A4(new_n593_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n401_), .B1(new_n308_), .B2(new_n317_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT74), .ZN(new_n600_));
  OAI211_X1 g399(.A(KEYINPUT35), .B(new_n593_), .C1(new_n599_), .C2(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n599_), .A2(new_n594_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n601_), .A2(new_n591_), .A3(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n598_), .A2(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G190gat), .B(G218gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(G134gat), .ZN(new_n606_));
  INV_X1    g405(.A(G162gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n609_), .A2(KEYINPUT36), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(KEYINPUT36), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n604_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT75), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n610_), .B1(new_n598_), .B2(new_n603_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n616_), .A2(KEYINPUT75), .A3(new_n612_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT37), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n598_), .A2(new_n603_), .A3(new_n610_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n618_), .A2(KEYINPUT76), .A3(new_n619_), .A4(new_n620_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n615_), .A2(new_n619_), .A3(new_n620_), .A4(new_n617_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT76), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n619_), .B1(new_n613_), .B2(new_n620_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n622_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n621_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n589_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(KEYINPUT104), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT104), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n630_), .B1(new_n589_), .B2(new_n627_), .ZN(new_n631_));
  AOI211_X1 g430(.A(G1gat), .B(new_n266_), .C1(new_n629_), .C2(new_n631_), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n632_), .A2(KEYINPUT38), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n618_), .A2(new_n620_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n589_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(G1gat), .B1(new_n637_), .B2(new_n266_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n632_), .A2(KEYINPUT38), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n633_), .A2(new_n638_), .A3(new_n639_), .ZN(G1324gat));
  INV_X1    g439(.A(new_n580_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n373_), .B1(new_n636_), .B2(new_n641_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT39), .Z(new_n643_));
  AOI21_X1  g442(.A(G8gat), .B1(new_n629_), .B2(new_n631_), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n644_), .A2(KEYINPUT105), .A3(new_n641_), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT105), .B1(new_n644_), .B2(new_n641_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n643_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT40), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n643_), .B(KEYINPUT40), .C1(new_n645_), .C2(new_n646_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1325gat));
  INV_X1    g450(.A(G15gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n628_), .A2(new_n652_), .A3(new_n581_), .ZN(new_n653_));
  OAI21_X1  g452(.A(G15gat), .B1(new_n637_), .B2(new_n548_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT41), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n654_), .A2(new_n655_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n653_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT106), .Z(G1326gat));
  INV_X1    g458(.A(G22gat), .ZN(new_n660_));
  INV_X1    g459(.A(new_n574_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n636_), .B2(new_n661_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT42), .Z(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n660_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT107), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n628_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n663_), .A2(new_n666_), .ZN(G1327gat));
  INV_X1    g466(.A(new_n434_), .ZN(new_n668_));
  AOI211_X1 g467(.A(new_n634_), .B(new_n668_), .C1(new_n575_), .C2(new_n587_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n669_), .A2(new_n422_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n266_), .ZN(new_n671_));
  AOI21_X1  g470(.A(G29gat), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n575_), .A2(new_n587_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(new_n627_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n673_), .A2(KEYINPUT43), .A3(new_n627_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n676_), .A2(new_n422_), .A3(new_n434_), .A4(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(KEYINPUT43), .B1(new_n673_), .B2(new_n627_), .ZN(new_n681_));
  AOI211_X1 g480(.A(new_n675_), .B(new_n626_), .C1(new_n575_), .C2(new_n587_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n683_), .A2(KEYINPUT44), .A3(new_n422_), .A4(new_n434_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n680_), .A2(new_n684_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n685_), .A2(G29gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n672_), .B1(new_n686_), .B2(new_n671_), .ZN(G1328gat));
  NAND3_X1  g486(.A1(new_n670_), .A2(new_n382_), .A3(new_n641_), .ZN(new_n688_));
  XOR2_X1   g487(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n689_));
  XNOR2_X1  g488(.A(new_n688_), .B(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n680_), .A2(new_n684_), .A3(new_n641_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(G36gat), .ZN(new_n692_));
  AOI22_X1  g491(.A1(new_n690_), .A2(new_n692_), .B1(KEYINPUT109), .B2(KEYINPUT46), .ZN(new_n693_));
  NOR2_X1   g492(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(G1329gat));
  NAND3_X1  g494(.A1(new_n680_), .A2(new_n684_), .A3(new_n581_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(G43gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n670_), .A2(new_n535_), .A3(new_n581_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(KEYINPUT110), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT110), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n697_), .A2(new_n701_), .A3(new_n698_), .ZN(new_n702_));
  AOI21_X1  g501(.A(KEYINPUT47), .B1(new_n700_), .B2(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n701_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n698_), .ZN(new_n705_));
  AOI211_X1 g504(.A(KEYINPUT110), .B(new_n705_), .C1(new_n696_), .C2(G43gat), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT47), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n704_), .A2(new_n706_), .A3(new_n707_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n703_), .A2(new_n708_), .ZN(G1330gat));
  AOI21_X1  g508(.A(G50gat), .B1(new_n670_), .B2(new_n661_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n661_), .A2(G50gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n685_), .B2(new_n711_), .ZN(G1331gat));
  NOR2_X1   g511(.A1(new_n368_), .A2(new_n369_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n421_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(new_n588_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n716_), .A2(new_n627_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT111), .Z(new_n718_));
  AOI21_X1  g517(.A(G57gat), .B1(new_n718_), .B2(new_n671_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n716_), .A2(new_n635_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n671_), .A2(G57gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n719_), .B1(new_n720_), .B2(new_n721_), .ZN(G1332gat));
  INV_X1    g521(.A(G64gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n723_), .B1(new_n720_), .B2(new_n641_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT48), .Z(new_n725_));
  NAND3_X1  g524(.A1(new_n718_), .A2(new_n723_), .A3(new_n641_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1333gat));
  INV_X1    g526(.A(G71gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n720_), .B2(new_n581_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT49), .Z(new_n730_));
  NAND3_X1  g529(.A1(new_n718_), .A2(new_n728_), .A3(new_n581_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1334gat));
  NAND2_X1  g531(.A1(new_n661_), .A2(new_n559_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT113), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n718_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n720_), .ZN(new_n736_));
  OAI21_X1  g535(.A(G78gat), .B1(new_n736_), .B2(new_n574_), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n737_), .A2(KEYINPUT112), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(KEYINPUT112), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n738_), .A2(KEYINPUT50), .A3(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(KEYINPUT50), .B1(new_n738_), .B2(new_n739_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n735_), .B1(new_n740_), .B2(new_n741_), .ZN(G1335gat));
  AND2_X1   g541(.A1(new_n715_), .A2(new_n669_), .ZN(new_n743_));
  AOI21_X1  g542(.A(G85gat), .B1(new_n743_), .B2(new_n671_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT114), .Z(new_n745_));
  NAND4_X1  g544(.A1(new_n676_), .A2(new_n434_), .A3(new_n677_), .A4(new_n715_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n746_), .A2(new_n286_), .A3(new_n266_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n745_), .A2(new_n747_), .ZN(G1336gat));
  NOR3_X1   g547(.A1(new_n746_), .A2(new_n287_), .A3(new_n580_), .ZN(new_n749_));
  AOI21_X1  g548(.A(G92gat), .B1(new_n743_), .B2(new_n641_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1337gat));
  NAND3_X1  g550(.A1(new_n743_), .A2(new_n279_), .A3(new_n581_), .ZN(new_n752_));
  OAI21_X1  g551(.A(G99gat), .B1(new_n746_), .B2(new_n548_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT115), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n753_), .A2(new_n754_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n752_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g558(.A(KEYINPUT117), .ZN(new_n760_));
  OR3_X1    g559(.A1(new_n746_), .A2(new_n760_), .A3(new_n574_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n746_), .B2(new_n574_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n761_), .A2(G106gat), .A3(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n743_), .A2(new_n280_), .A3(new_n661_), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT116), .Z(new_n767_));
  NAND4_X1  g566(.A1(new_n761_), .A2(KEYINPUT52), .A3(G106gat), .A4(new_n762_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n765_), .A2(new_n767_), .A3(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(KEYINPUT53), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT53), .ZN(new_n771_));
  NAND4_X1  g570(.A1(new_n765_), .A2(new_n767_), .A3(new_n771_), .A4(new_n768_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(G1339gat));
  NOR2_X1   g572(.A1(new_n266_), .A2(new_n641_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n268_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n357_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n339_), .A2(KEYINPUT55), .A3(new_n268_), .A4(new_n340_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n347_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n780_), .A2(KEYINPUT56), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n406_), .A2(new_n403_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n414_), .B(new_n783_), .C1(new_n402_), .C2(new_n403_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n418_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT56), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n361_), .B1(new_n779_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n782_), .A2(new_n785_), .A3(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT58), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT58), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n782_), .A2(new_n791_), .A3(new_n785_), .A4(new_n788_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n626_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n364_), .A2(new_n785_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT119), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n714_), .A2(new_n782_), .A3(new_n788_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT119), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n364_), .A2(new_n797_), .A3(new_n785_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n795_), .A2(new_n796_), .A3(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n634_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n793_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n799_), .A2(KEYINPUT57), .A3(new_n634_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n668_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n365_), .A2(new_n367_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n434_), .B1(new_n621_), .B2(new_n625_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT118), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n805_), .A2(new_n806_), .A3(new_n807_), .A4(new_n421_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(KEYINPUT54), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n805_), .A2(new_n806_), .A3(new_n421_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(KEYINPUT118), .A3(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(KEYINPUT118), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n812_), .A2(KEYINPUT54), .A3(new_n808_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n813_), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n586_), .B(new_n774_), .C1(new_n804_), .C2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(G113gat), .B1(new_n816_), .B2(new_n714_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT59), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n815_), .A2(new_n818_), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n364_), .A2(new_n797_), .A3(new_n785_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n797_), .B1(new_n364_), .B2(new_n785_), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n421_), .A2(new_n781_), .A3(new_n787_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n820_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n801_), .B1(new_n823_), .B2(new_n635_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n793_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n824_), .A2(new_n825_), .A3(new_n803_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n434_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n809_), .B(new_n812_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n829_), .A2(KEYINPUT59), .A3(new_n586_), .A4(new_n774_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n421_), .B1(new_n819_), .B2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n817_), .B1(new_n831_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g631(.A(G120gat), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n833_), .B1(new_n713_), .B2(KEYINPUT60), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n816_), .B(new_n834_), .C1(KEYINPUT60), .C2(new_n833_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n713_), .B1(new_n819_), .B2(new_n830_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(new_n833_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT121), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n835_), .B(KEYINPUT121), .C1(new_n836_), .C2(new_n833_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(G1341gat));
  AOI21_X1  g640(.A(G127gat), .B1(new_n816_), .B2(new_n668_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n434_), .B1(new_n819_), .B2(new_n830_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g643(.A(G134gat), .B1(new_n816_), .B2(new_n635_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n626_), .B1(new_n819_), .B2(new_n830_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(G134gat), .ZN(G1343gat));
  AND2_X1   g646(.A1(new_n829_), .A2(new_n585_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n774_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n849_), .A2(new_n421_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(new_n205_), .ZN(G1344gat));
  NOR2_X1   g650(.A1(new_n849_), .A2(new_n713_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(new_n206_), .ZN(G1345gat));
  NOR2_X1   g652(.A1(new_n849_), .A2(new_n434_), .ZN(new_n854_));
  XOR2_X1   g653(.A(KEYINPUT61), .B(G155gat), .Z(new_n855_));
  XNOR2_X1  g654(.A(new_n854_), .B(new_n855_), .ZN(G1346gat));
  NOR3_X1   g655(.A1(new_n849_), .A2(new_n607_), .A3(new_n626_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n849_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n635_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n857_), .B1(new_n607_), .B2(new_n859_), .ZN(G1347gat));
  NOR2_X1   g659(.A1(new_n661_), .A2(new_n421_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n671_), .A2(new_n548_), .A3(new_n580_), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n861_), .B(new_n862_), .C1(new_n804_), .C2(new_n814_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT122), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n829_), .A2(new_n865_), .A3(new_n861_), .A4(new_n862_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n864_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT62), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n867_), .A2(KEYINPUT123), .A3(new_n868_), .A4(G169gat), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n864_), .A2(new_n866_), .A3(G169gat), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(KEYINPUT62), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT123), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n872_), .B1(new_n870_), .B2(KEYINPUT62), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n869_), .A2(new_n871_), .A3(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n671_), .A2(new_n580_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n829_), .A2(new_n586_), .A3(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT124), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n876_), .A2(new_n877_), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n714_), .B(new_n438_), .C1(new_n879_), .C2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n874_), .A2(new_n881_), .ZN(G1348gat));
  INV_X1    g681(.A(new_n713_), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n346_), .B(new_n883_), .C1(new_n879_), .C2(new_n880_), .ZN(new_n884_));
  OAI21_X1  g683(.A(G176gat), .B1(new_n876_), .B2(new_n713_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1349gat));
  INV_X1    g685(.A(new_n876_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n441_), .B1(new_n887_), .B2(new_n668_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n880_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n434_), .B1(new_n889_), .B2(new_n878_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n888_), .B1(new_n890_), .B2(new_n471_), .ZN(G1350gat));
  NOR2_X1   g690(.A1(new_n634_), .A2(new_n452_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n892_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n626_), .B1(new_n889_), .B2(new_n878_), .ZN(new_n894_));
  INV_X1    g693(.A(G190gat), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n893_), .B1(new_n894_), .B2(new_n895_), .ZN(G1351gat));
  NAND3_X1  g695(.A1(new_n829_), .A2(new_n585_), .A3(new_n875_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n421_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(new_n413_), .ZN(G1352gat));
  INV_X1    g698(.A(new_n897_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n883_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n901_), .B1(KEYINPUT125), .B2(G204gat), .ZN(new_n902_));
  NAND2_X1  g701(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n903_));
  MUX2_X1   g702(.A(new_n901_), .B(new_n902_), .S(new_n903_), .Z(G1353gat));
  INV_X1    g703(.A(KEYINPUT63), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n434_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  OR3_X1    g706(.A1(new_n897_), .A2(KEYINPUT126), .A3(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(G211gat), .ZN(new_n909_));
  OAI21_X1  g708(.A(KEYINPUT126), .B1(new_n897_), .B2(new_n907_), .ZN(new_n910_));
  AND4_X1   g709(.A1(new_n905_), .A2(new_n908_), .A3(new_n909_), .A4(new_n910_), .ZN(new_n911_));
  AOI22_X1  g710(.A1(new_n908_), .A2(new_n910_), .B1(new_n905_), .B2(new_n909_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1354gat));
  XNOR2_X1  g712(.A(KEYINPUT127), .B(G218gat), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n914_), .B1(new_n900_), .B2(new_n635_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n897_), .A2(new_n626_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n915_), .B1(new_n914_), .B2(new_n916_), .ZN(G1355gat));
endmodule


