//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 0 0 0 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0 0 1 0 1 0 0 1 0 1 0 1 0 0 0 0 0 0 0 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n905_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n938_, new_n939_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n949_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n956_, new_n957_, new_n958_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT4), .ZN(new_n203_));
  INV_X1    g002(.A(G134gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G127gat), .ZN(new_n205_));
  INV_X1    g004(.A(G127gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G134gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n205_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G120gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G113gat), .ZN(new_n210_));
  INV_X1    g009(.A(G113gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G120gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n208_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT83), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n205_), .A2(new_n207_), .A3(new_n210_), .A4(new_n212_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n208_), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n218_), .A2(KEYINPUT83), .A3(new_n210_), .A4(new_n212_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n221_));
  INV_X1    g020(.A(G141gat), .ZN(new_n222_));
  INV_X1    g021(.A(G148gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G141gat), .A2(G148gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT2), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n224_), .A2(new_n227_), .A3(new_n228_), .A4(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G155gat), .A2(G162gat), .ZN(new_n231_));
  OR2_X1    g030(.A1(G155gat), .A2(G162gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n222_), .A2(new_n223_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n231_), .A2(KEYINPUT1), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(new_n232_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n231_), .A2(KEYINPUT1), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n234_), .B(new_n225_), .C1(new_n236_), .C2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n233_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n220_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n214_), .A2(new_n216_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n233_), .A2(new_n241_), .A3(new_n238_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n203_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(KEYINPUT4), .B1(new_n220_), .B2(new_n239_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n202_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G1gat), .B(G29gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G57gat), .B(G85gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT95), .ZN(new_n252_));
  AOI22_X1  g051(.A1(new_n219_), .A2(new_n217_), .B1(new_n233_), .B2(new_n238_), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n233_), .A2(new_n241_), .A3(new_n238_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n252_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n240_), .A2(KEYINPUT95), .A3(new_n242_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n202_), .B(KEYINPUT93), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n245_), .A2(new_n251_), .A3(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n240_), .A2(new_n242_), .A3(new_n202_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n240_), .A2(new_n242_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n244_), .B1(new_n261_), .B2(KEYINPUT4), .ZN(new_n262_));
  INV_X1    g061(.A(new_n257_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n260_), .B(new_n250_), .C1(new_n262_), .C2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT33), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n257_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT33), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n266_), .A2(new_n267_), .A3(new_n260_), .A4(new_n250_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n259_), .B1(new_n265_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G226gat), .A2(G233gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT19), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G169gat), .A2(G176gat), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT80), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(G169gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n275_), .A2(KEYINPUT81), .A3(KEYINPUT22), .ZN(new_n276_));
  INV_X1    g075(.A(G176gat), .ZN(new_n277_));
  AND2_X1   g076(.A1(KEYINPUT81), .A2(KEYINPUT22), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n276_), .B(new_n277_), .C1(new_n275_), .C2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G183gat), .A2(G190gat), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT23), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n283_));
  INV_X1    g082(.A(G183gat), .ZN(new_n284_));
  INV_X1    g083(.A(G190gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n282_), .A2(new_n283_), .A3(new_n286_), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n274_), .A2(new_n279_), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT24), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT79), .B1(G169gat), .B2(G176gat), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NOR3_X1   g090(.A1(KEYINPUT79), .A2(G169gat), .A3(G176gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n289_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n280_), .A2(KEYINPUT23), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n281_), .A2(G183gat), .A3(G190gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n284_), .A2(KEYINPUT25), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT25), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(G183gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n285_), .A2(KEYINPUT26), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT26), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(G190gat), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n297_), .A2(new_n299_), .A3(new_n300_), .A4(new_n302_), .ZN(new_n303_));
  AND3_X1   g102(.A1(new_n293_), .A2(new_n296_), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n292_), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n274_), .A2(KEYINPUT24), .A3(new_n305_), .A4(new_n290_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n288_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(G204gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT85), .B1(new_n308_), .B2(G197gat), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT85), .ZN(new_n310_));
  INV_X1    g109(.A(G197gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n310_), .A2(new_n311_), .A3(G204gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n308_), .A2(G197gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n309_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT89), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G211gat), .B(G218gat), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT21), .B1(new_n317_), .B2(KEYINPUT88), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n318_), .B1(KEYINPUT88), .B2(new_n317_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n316_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n317_), .ZN(new_n321_));
  AND3_X1   g120(.A1(new_n309_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n322_));
  AND2_X1   g121(.A1(KEYINPUT86), .A2(KEYINPUT21), .ZN(new_n323_));
  NOR2_X1   g122(.A1(KEYINPUT86), .A2(KEYINPUT21), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n321_), .B1(new_n322_), .B2(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT84), .B1(new_n308_), .B2(G197gat), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT84), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n328_), .A2(new_n311_), .A3(G204gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n329_), .A3(new_n313_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT21), .ZN(new_n331_));
  AOI21_X1  g130(.A(KEYINPUT87), .B1(new_n326_), .B2(new_n331_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n325_), .A2(new_n313_), .A3(new_n309_), .A4(new_n312_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n331_), .A2(new_n333_), .A3(KEYINPUT87), .A4(new_n317_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n307_), .B(new_n320_), .C1(new_n332_), .C2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT20), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT87), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n333_), .A2(new_n317_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n330_), .A2(KEYINPUT21), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n338_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  AOI22_X1  g140(.A1(new_n341_), .A2(new_n334_), .B1(new_n316_), .B2(new_n319_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n305_), .A2(KEYINPUT24), .A3(new_n272_), .A4(new_n290_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n343_), .A2(new_n293_), .A3(new_n296_), .A4(new_n303_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT22), .B(G169gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(new_n277_), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n294_), .A2(new_n295_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT90), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n274_), .B(new_n346_), .C1(new_n347_), .C2(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n287_), .A2(KEYINPUT90), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n344_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n342_), .A2(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n271_), .B1(new_n337_), .B2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G8gat), .B(G36gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G64gat), .B(G92gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT20), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n320_), .B1(new_n332_), .B2(new_n335_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n307_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n360_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n271_), .B1(new_n342_), .B2(new_n352_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n354_), .A2(new_n359_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT92), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n354_), .A2(KEYINPUT92), .A3(new_n365_), .A4(new_n359_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n354_), .A2(new_n365_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n359_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n269_), .A2(new_n368_), .A3(new_n369_), .A4(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT96), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n359_), .B1(new_n354_), .B2(new_n365_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n375_), .B1(new_n367_), .B2(new_n366_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT96), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n376_), .A2(new_n377_), .A3(new_n369_), .A4(new_n269_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n359_), .A2(KEYINPUT32), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n354_), .A2(new_n365_), .A3(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT4), .B1(new_n253_), .B2(new_n254_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n244_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n263_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n260_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n251_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(new_n264_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n380_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT97), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n351_), .A2(new_n388_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n344_), .B(KEYINPUT97), .C1(new_n350_), .C2(new_n349_), .ZN(new_n390_));
  AND3_X1   g189(.A1(new_n342_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT20), .B1(new_n342_), .B2(new_n307_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n271_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n361_), .A2(new_n351_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n271_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n394_), .A2(KEYINPUT20), .A3(new_n395_), .A4(new_n336_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n379_), .B1(new_n393_), .B2(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n387_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n374_), .A2(new_n378_), .A3(new_n399_), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n239_), .A2(KEYINPUT29), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n401_), .A2(KEYINPUT28), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(KEYINPUT28), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n239_), .A2(KEYINPUT29), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n404_), .A2(new_n361_), .A3(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n361_), .A2(new_n405_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n407_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G228gat), .A2(G233gat), .ZN(new_n409_));
  INV_X1    g208(.A(G78gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(G106gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G22gat), .B(G50gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n406_), .A2(new_n408_), .A3(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n415_), .B1(new_n406_), .B2(new_n408_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n396_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n342_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n395_), .B1(new_n363_), .B2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n371_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT98), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT98), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n424_), .B(new_n371_), .C1(new_n419_), .C2(new_n421_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n366_), .A2(KEYINPUT27), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n368_), .A2(new_n369_), .A3(new_n372_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT27), .ZN(new_n429_));
  AOI22_X1  g228(.A1(new_n426_), .A2(new_n427_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n418_), .A2(new_n386_), .ZN(new_n431_));
  AOI22_X1  g230(.A1(new_n400_), .A2(new_n418_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n220_), .B(KEYINPUT31), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n433_), .A2(KEYINPUT82), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G227gat), .A2(G233gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(G15gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT30), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n307_), .B(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n434_), .B(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G71gat), .B(G99gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(G43gat), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n439_), .A2(new_n441_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT99), .B1(new_n432_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n430_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n418_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n444_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n449_), .A2(new_n386_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT99), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n398_), .B1(new_n373_), .B2(KEYINPUT96), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n447_), .B1(new_n453_), .B2(new_n378_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n426_), .A2(new_n427_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n428_), .A2(new_n429_), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n455_), .A2(new_n456_), .A3(new_n431_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n452_), .B(new_n449_), .C1(new_n454_), .C2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n445_), .A2(new_n451_), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT37), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT74), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n460_), .A2(KEYINPUT74), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G29gat), .B(G36gat), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G43gat), .B(G50gat), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n463_), .A2(new_n465_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT64), .B(G92gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(G85gat), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT9), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n475_), .A2(KEYINPUT65), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT65), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n477_), .B1(G85gat), .B2(G92gat), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n476_), .B1(new_n475_), .B2(new_n478_), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n474_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G99gat), .A2(G106gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT6), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT10), .B(G99gat), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n482_), .B1(G106gat), .B2(new_n483_), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n480_), .A2(new_n484_), .ZN(new_n485_));
  XOR2_X1   g284(.A(G85gat), .B(G92gat), .Z(new_n486_));
  OR2_X1    g285(.A1(G99gat), .A2(G106gat), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n482_), .B1(KEYINPUT7), .B2(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT66), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n486_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT8), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n492_), .A2(KEYINPUT67), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n491_), .A2(new_n493_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n470_), .B(new_n485_), .C1(new_n494_), .C2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT15), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n469_), .A2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n467_), .A2(KEYINPUT15), .A3(new_n468_), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n480_), .A2(new_n484_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n491_), .A2(new_n493_), .ZN(new_n502_));
  OAI221_X1 g301(.A(new_n486_), .B1(KEYINPUT67), .B2(new_n492_), .C1(new_n488_), .C2(new_n490_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n501_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n496_), .B1(new_n500_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT72), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G232gat), .A2(G233gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT34), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT35), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n506_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n505_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT69), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n509_), .A2(new_n510_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n512_), .A2(new_n513_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n505_), .A2(KEYINPUT69), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(new_n514_), .ZN(new_n518_));
  AOI21_X1  g317(.A(KEYINPUT69), .B1(new_n505_), .B2(new_n511_), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n516_), .B(KEYINPUT73), .C1(new_n518_), .C2(new_n519_), .ZN(new_n520_));
  XOR2_X1   g319(.A(G190gat), .B(G218gat), .Z(new_n521_));
  XNOR2_X1  g320(.A(G134gat), .B(G162gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(KEYINPUT70), .B(KEYINPUT71), .Z(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT36), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n516_), .B(new_n527_), .C1(new_n518_), .C2(new_n519_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n525_), .A2(new_n526_), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n520_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n520_), .B1(new_n529_), .B2(new_n528_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n461_), .B(new_n462_), .C1(new_n530_), .C2(new_n531_), .ZN(new_n532_));
  AOI211_X1 g331(.A(KEYINPUT69), .B(new_n514_), .C1(new_n505_), .C2(new_n511_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n518_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n519_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n533_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n529_), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n536_), .B(KEYINPUT73), .C1(new_n537_), .C2(new_n527_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n520_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n538_), .A2(KEYINPUT74), .A3(new_n460_), .A4(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n532_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G57gat), .B(G64gat), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n542_), .A2(KEYINPUT11), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(KEYINPUT11), .ZN(new_n544_));
  XOR2_X1   g343(.A(G71gat), .B(G78gat), .Z(new_n545_));
  NAND3_X1  g344(.A1(new_n543_), .A2(new_n544_), .A3(new_n545_), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n544_), .A2(new_n545_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G231gat), .A2(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT75), .B(G1gat), .ZN(new_n551_));
  INV_X1    g350(.A(G8gat), .ZN(new_n552_));
  OAI21_X1  g351(.A(KEYINPUT14), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G15gat), .B(G22gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G1gat), .B(G8gat), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n553_), .A2(new_n554_), .A3(new_n556_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n550_), .B(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(G127gat), .B(G155gat), .Z(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT16), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G183gat), .B(G211gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT17), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n565_), .A2(new_n566_), .ZN(new_n568_));
  NOR3_X1   g367(.A1(new_n561_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n561_), .A2(new_n567_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n541_), .A2(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(G120gat), .B(G148gat), .Z(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G176gat), .B(G204gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n485_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n548_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n504_), .A2(new_n548_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(KEYINPUT12), .A3(new_n583_), .ZN(new_n584_));
  OR3_X1    g383(.A1(new_n504_), .A2(KEYINPUT12), .A3(new_n548_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G230gat), .A2(G233gat), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n587_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n579_), .B1(new_n588_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n587_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n592_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n593_), .A2(new_n589_), .A3(new_n578_), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n591_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT13), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n591_), .A2(new_n594_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT13), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n560_), .A2(new_n469_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n498_), .A2(new_n559_), .A3(new_n558_), .A4(new_n499_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G229gat), .A2(G233gat), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n602_), .A2(new_n603_), .A3(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT76), .ZN(new_n606_));
  INV_X1    g405(.A(new_n604_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n602_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n560_), .A2(new_n469_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n607_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT76), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n602_), .A2(new_n603_), .A3(new_n611_), .A4(new_n604_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n606_), .A2(new_n610_), .A3(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G113gat), .B(G141gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT77), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G169gat), .B(G197gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n613_), .A2(new_n618_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n606_), .A2(new_n610_), .A3(new_n612_), .A4(new_n617_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT78), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n620_), .A2(new_n621_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n619_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n601_), .A2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n459_), .A2(new_n573_), .A3(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT100), .Z(new_n629_));
  NAND3_X1  g428(.A1(new_n629_), .A2(new_n551_), .A3(new_n386_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT38), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n530_), .A2(new_n531_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n459_), .A2(new_n633_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n597_), .A2(new_n599_), .A3(new_n571_), .A4(new_n625_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT101), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n386_), .ZN(new_n639_));
  OAI21_X1  g438(.A(G1gat), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n630_), .A2(new_n631_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n632_), .A2(new_n640_), .A3(new_n641_), .ZN(G1324gat));
  NAND3_X1  g441(.A1(new_n629_), .A2(new_n552_), .A3(new_n446_), .ZN(new_n643_));
  AND4_X1   g442(.A1(new_n633_), .A2(new_n636_), .A3(new_n459_), .A4(new_n446_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT102), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT39), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n552_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n646_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n647_), .B1(new_n646_), .B2(new_n648_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n643_), .B1(new_n649_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT40), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  OAI211_X1 g452(.A(KEYINPUT40), .B(new_n643_), .C1(new_n649_), .C2(new_n650_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1325gat));
  OAI21_X1  g454(.A(G15gat), .B1(new_n638_), .B2(new_n449_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n657_), .ZN(new_n659_));
  INV_X1    g458(.A(G15gat), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n629_), .A2(new_n660_), .A3(new_n444_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n658_), .A2(new_n659_), .A3(new_n661_), .ZN(G1326gat));
  INV_X1    g461(.A(G22gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n663_), .B1(new_n637_), .B2(new_n447_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n629_), .A2(new_n663_), .A3(new_n447_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1327gat));
  NOR2_X1   g467(.A1(new_n633_), .A2(new_n571_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n459_), .A2(new_n627_), .A3(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n459_), .A2(KEYINPUT106), .A3(new_n627_), .A4(new_n669_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(G29gat), .B1(new_n674_), .B2(new_n386_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n627_), .A2(new_n572_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n400_), .A2(new_n418_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n430_), .A2(new_n431_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n452_), .B1(new_n679_), .B2(new_n449_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n458_), .A2(new_n451_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n541_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT43), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT43), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n459_), .A2(new_n684_), .A3(new_n541_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n676_), .B1(new_n683_), .B2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(KEYINPUT105), .B1(new_n686_), .B2(KEYINPUT44), .ZN(new_n687_));
  INV_X1    g486(.A(new_n676_), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n459_), .A2(new_n684_), .A3(new_n541_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n684_), .B1(new_n459_), .B2(new_n541_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n688_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n691_), .A2(new_n692_), .A3(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n687_), .A2(new_n694_), .ZN(new_n695_));
  OAI211_X1 g494(.A(KEYINPUT44), .B(new_n688_), .C1(new_n689_), .C2(new_n690_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n386_), .A2(G29gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n675_), .B1(new_n698_), .B2(new_n699_), .ZN(G1328gat));
  INV_X1    g499(.A(KEYINPUT108), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n701_), .A2(KEYINPUT46), .ZN(new_n702_));
  INV_X1    g501(.A(G36gat), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n696_), .A2(new_n446_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n703_), .B1(new_n695_), .B2(new_n705_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n672_), .A2(new_n703_), .A3(new_n446_), .A4(new_n673_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n707_), .B(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n702_), .B1(new_n706_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n708_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n707_), .B(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n704_), .B1(new_n687_), .B2(new_n694_), .ZN(new_n713_));
  OAI221_X1 g512(.A(new_n712_), .B1(new_n701_), .B2(KEYINPUT46), .C1(new_n713_), .C2(new_n703_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n710_), .A2(new_n714_), .ZN(G1329gat));
  NAND2_X1  g514(.A1(new_n444_), .A2(G43gat), .ZN(new_n716_));
  INV_X1    g515(.A(new_n696_), .ZN(new_n717_));
  AOI211_X1 g516(.A(new_n716_), .B(new_n717_), .C1(new_n687_), .C2(new_n694_), .ZN(new_n718_));
  AOI21_X1  g517(.A(G43gat), .B1(new_n674_), .B2(new_n444_), .ZN(new_n719_));
  OAI21_X1  g518(.A(KEYINPUT47), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT47), .ZN(new_n721_));
  INV_X1    g520(.A(new_n719_), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n721_), .B(new_n722_), .C1(new_n697_), .C2(new_n716_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n720_), .A2(new_n723_), .ZN(G1330gat));
  AOI21_X1  g523(.A(G50gat), .B1(new_n674_), .B2(new_n447_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n447_), .A2(G50gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n698_), .B2(new_n726_), .ZN(G1331gat));
  NOR2_X1   g526(.A1(new_n572_), .A2(new_n625_), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n634_), .A2(new_n601_), .A3(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(new_n386_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(G57gat), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n459_), .A2(new_n626_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n600_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n459_), .A2(KEYINPUT109), .A3(new_n626_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(new_n573_), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n639_), .A2(G57gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n731_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT110), .ZN(G1332gat));
  INV_X1    g539(.A(G64gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n729_), .B2(new_n446_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT48), .Z(new_n743_));
  INV_X1    g542(.A(new_n737_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n744_), .A2(new_n741_), .A3(new_n446_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1333gat));
  NAND2_X1  g545(.A1(new_n729_), .A2(new_n444_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(G71gat), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT49), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n449_), .A2(G71gat), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n749_), .B1(new_n737_), .B2(new_n750_), .ZN(G1334gat));
  AOI21_X1  g550(.A(new_n410_), .B1(new_n729_), .B2(new_n447_), .ZN(new_n752_));
  XOR2_X1   g551(.A(new_n752_), .B(KEYINPUT50), .Z(new_n753_));
  NAND3_X1  g552(.A1(new_n744_), .A2(new_n410_), .A3(new_n447_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1335gat));
  NAND3_X1  g554(.A1(new_n734_), .A2(new_n669_), .A3(new_n735_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT111), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT111), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n734_), .A2(new_n758_), .A3(new_n669_), .A4(new_n735_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(G85gat), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n760_), .A2(new_n761_), .A3(new_n386_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n683_), .A2(new_n685_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n600_), .A2(new_n571_), .A3(new_n625_), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n763_), .A2(new_n386_), .A3(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n762_), .B1(new_n761_), .B2(new_n765_), .ZN(G1336gat));
  NAND4_X1  g565(.A1(new_n763_), .A2(new_n471_), .A3(new_n446_), .A4(new_n764_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n430_), .B1(new_n757_), .B2(new_n759_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(G92gat), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT112), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n767_), .B(KEYINPUT112), .C1(new_n768_), .C2(G92gat), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(G1337gat));
  OAI211_X1 g572(.A(new_n444_), .B(new_n764_), .C1(new_n689_), .C2(new_n690_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(G99gat), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT113), .ZN(new_n776_));
  INV_X1    g575(.A(new_n483_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n444_), .A2(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n778_), .B1(new_n757_), .B2(new_n759_), .ZN(new_n779_));
  OAI21_X1  g578(.A(KEYINPUT51), .B1(new_n776_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n775_), .B(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n779_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT51), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n782_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n780_), .A2(new_n785_), .ZN(G1338gat));
  NAND3_X1  g585(.A1(new_n763_), .A2(new_n447_), .A3(new_n764_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(G106gat), .ZN(new_n788_));
  XOR2_X1   g587(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n787_), .A2(G106gat), .A3(new_n789_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n447_), .A2(new_n412_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n794_), .B1(new_n757_), .B2(new_n759_), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT53), .B1(new_n793_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n795_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n797_), .A2(new_n798_), .A3(new_n792_), .A4(new_n791_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n796_), .A2(new_n799_), .ZN(G1339gat));
  NAND3_X1  g599(.A1(new_n448_), .A2(new_n444_), .A3(new_n386_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT58), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT56), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n803_), .A2(KEYINPUT119), .ZN(new_n804_));
  AND3_X1   g603(.A1(new_n584_), .A2(new_n592_), .A3(new_n585_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n805_), .A2(new_n593_), .A3(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n586_), .A2(new_n806_), .A3(new_n587_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n578_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n804_), .B1(new_n807_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n594_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n584_), .A2(new_n592_), .A3(new_n585_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n588_), .A2(KEYINPUT55), .A3(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n579_), .B1(new_n593_), .B2(new_n806_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n813_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n810_), .A2(new_n811_), .A3(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n818_));
  INV_X1    g617(.A(new_n624_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n622_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n604_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n602_), .A2(new_n603_), .A3(new_n607_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n821_), .A2(new_n618_), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n818_), .B1(new_n820_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n823_), .ZN(new_n825_));
  AOI211_X1 g624(.A(KEYINPUT116), .B(new_n825_), .C1(new_n819_), .C2(new_n622_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n824_), .A2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n802_), .B1(new_n817_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n813_), .A2(new_n814_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n594_), .B1(new_n829_), .B2(new_n804_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n823_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT116), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n820_), .A2(new_n818_), .A3(new_n823_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n830_), .A2(new_n834_), .A3(KEYINPUT58), .A4(new_n816_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n541_), .A2(new_n828_), .A3(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT120), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n541_), .A2(new_n828_), .A3(new_n835_), .A4(KEYINPUT120), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT117), .B1(new_n841_), .B2(KEYINPUT57), .ZN(new_n842_));
  NOR2_X1   g641(.A1(KEYINPUT115), .A2(KEYINPUT56), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n813_), .A2(new_n814_), .A3(new_n844_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n844_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n625_), .B(new_n811_), .C1(new_n845_), .C2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n595_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n842_), .B1(new_n849_), .B2(new_n633_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT117), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n811_), .A2(new_n625_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n829_), .A2(new_n843_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n813_), .A2(new_n814_), .A3(new_n844_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n852_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n598_), .B1(new_n833_), .B2(new_n832_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n851_), .B(new_n633_), .C1(new_n855_), .C2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n841_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n850_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n572_), .B1(new_n840_), .B2(new_n860_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n600_), .A2(new_n540_), .A3(new_n532_), .A4(new_n728_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT54), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n801_), .B1(new_n861_), .B2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(G113gat), .B1(new_n864_), .B2(new_n625_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n801_), .A2(KEYINPUT59), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n849_), .A2(new_n633_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n842_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n538_), .A2(new_n539_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n870_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n871_));
  AOI21_X1  g670(.A(KEYINPUT118), .B1(new_n871_), .B2(new_n851_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n869_), .B1(new_n872_), .B2(KEYINPUT57), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n571_), .B1(new_n873_), .B2(new_n836_), .ZN(new_n874_));
  XOR2_X1   g673(.A(new_n862_), .B(KEYINPUT54), .Z(new_n875_));
  OAI21_X1  g674(.A(new_n866_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n864_), .B2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n211_), .B1(new_n625_), .B2(KEYINPUT121), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n880_), .B1(KEYINPUT121), .B2(new_n211_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n865_), .B1(new_n879_), .B2(new_n881_), .ZN(G1340gat));
  OAI211_X1 g681(.A(new_n601_), .B(new_n876_), .C1(new_n864_), .C2(new_n877_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(G120gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n209_), .B1(new_n600_), .B2(KEYINPUT60), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n864_), .B(new_n885_), .C1(KEYINPUT60), .C2(new_n209_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT122), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n884_), .A2(KEYINPUT122), .A3(new_n886_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1341gat));
  OAI21_X1  g690(.A(G127gat), .B1(new_n878_), .B2(new_n572_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n864_), .A2(new_n206_), .A3(new_n571_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(G1342gat));
  AOI21_X1  g693(.A(G134gat), .B1(new_n864_), .B2(new_n870_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n541_), .ZN(new_n896_));
  XOR2_X1   g695(.A(KEYINPUT123), .B(G134gat), .Z(new_n897_));
  NOR2_X1   g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n895_), .B1(new_n879_), .B2(new_n898_), .ZN(G1343gat));
  NAND2_X1  g698(.A1(new_n861_), .A2(new_n863_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n444_), .A2(new_n639_), .A3(new_n418_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n900_), .A2(new_n430_), .A3(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(new_n626_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(new_n222_), .ZN(G1344gat));
  NOR2_X1   g703(.A1(new_n902_), .A2(new_n600_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(new_n223_), .ZN(G1345gat));
  NOR2_X1   g705(.A1(new_n902_), .A2(new_n572_), .ZN(new_n907_));
  XOR2_X1   g706(.A(KEYINPUT61), .B(G155gat), .Z(new_n908_));
  XNOR2_X1  g707(.A(new_n907_), .B(new_n908_), .ZN(G1346gat));
  OAI21_X1  g708(.A(G162gat), .B1(new_n902_), .B2(new_n896_), .ZN(new_n910_));
  OR2_X1    g709(.A1(new_n633_), .A2(G162gat), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n902_), .B2(new_n911_), .ZN(G1347gat));
  INV_X1    g711(.A(KEYINPUT124), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n446_), .A2(new_n418_), .A3(new_n450_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n916_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n917_), .A2(new_n626_), .ZN(new_n918_));
  OAI211_X1 g717(.A(new_n913_), .B(new_n914_), .C1(new_n918_), .C2(new_n275_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n345_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n275_), .B1(KEYINPUT124), .B2(KEYINPUT62), .ZN(new_n921_));
  OAI221_X1 g720(.A(new_n921_), .B1(KEYINPUT124), .B2(KEYINPUT62), .C1(new_n917_), .C2(new_n626_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n919_), .A2(new_n920_), .A3(new_n922_), .ZN(G1348gat));
  INV_X1    g722(.A(new_n917_), .ZN(new_n924_));
  AOI21_X1  g723(.A(G176gat), .B1(new_n924_), .B2(new_n601_), .ZN(new_n925_));
  NAND4_X1  g724(.A1(new_n900_), .A2(G176gat), .A3(new_n601_), .A4(new_n916_), .ZN(new_n926_));
  OR2_X1    g725(.A1(new_n926_), .A2(KEYINPUT125), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(KEYINPUT125), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n925_), .B1(new_n927_), .B2(new_n928_), .ZN(G1349gat));
  AND2_X1   g728(.A1(new_n861_), .A2(new_n863_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n930_), .A2(new_n915_), .ZN(new_n931_));
  AOI21_X1  g730(.A(G183gat), .B1(new_n931_), .B2(new_n571_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n572_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n934_));
  AND3_X1   g733(.A1(new_n924_), .A2(new_n933_), .A3(new_n934_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n933_), .B1(new_n924_), .B2(new_n934_), .ZN(new_n936_));
  NOR3_X1   g735(.A1(new_n932_), .A2(new_n935_), .A3(new_n936_), .ZN(G1350gat));
  OAI21_X1  g736(.A(G190gat), .B1(new_n917_), .B2(new_n896_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n870_), .A2(new_n300_), .A3(new_n302_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n938_), .B1(new_n917_), .B2(new_n939_), .ZN(G1351gat));
  INV_X1    g739(.A(KEYINPUT127), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n446_), .A2(new_n449_), .A3(new_n431_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n930_), .A2(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(new_n625_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n941_), .B1(new_n944_), .B2(new_n311_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n311_), .ZN(new_n946_));
  NAND4_X1  g745(.A1(new_n943_), .A2(KEYINPUT127), .A3(G197gat), .A4(new_n625_), .ZN(new_n947_));
  AND3_X1   g746(.A1(new_n945_), .A2(new_n946_), .A3(new_n947_), .ZN(G1352gat));
  NAND2_X1  g747(.A1(new_n943_), .A2(new_n601_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n949_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g749(.A1(new_n943_), .A2(new_n571_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n952_));
  AND2_X1   g751(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n953_));
  NOR3_X1   g752(.A1(new_n951_), .A2(new_n952_), .A3(new_n953_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n954_), .B1(new_n951_), .B2(new_n952_), .ZN(G1354gat));
  INV_X1    g754(.A(new_n943_), .ZN(new_n956_));
  OR3_X1    g755(.A1(new_n956_), .A2(G218gat), .A3(new_n633_), .ZN(new_n957_));
  OAI21_X1  g756(.A(G218gat), .B1(new_n956_), .B2(new_n896_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n957_), .A2(new_n958_), .ZN(G1355gat));
endmodule


