//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n766_, new_n767_, new_n768_, new_n769_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n897_, new_n898_, new_n899_, new_n900_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n933_, new_n934_, new_n936_, new_n937_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n954_, new_n955_;
  AND2_X1   g000(.A1(KEYINPUT83), .A2(G169gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(KEYINPUT83), .A2(G169gat), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT22), .B1(new_n202_), .B2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT84), .ZN(new_n205_));
  INV_X1    g004(.A(G176gat), .ZN(new_n206_));
  INV_X1    g005(.A(G169gat), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n207_), .A2(KEYINPUT22), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT84), .ZN(new_n209_));
  OAI211_X1 g008(.A(new_n209_), .B(KEYINPUT22), .C1(new_n202_), .C2(new_n203_), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n205_), .A2(new_n206_), .A3(new_n208_), .A4(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G183gat), .ZN(new_n214_));
  INV_X1    g013(.A(G190gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n213_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n211_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT24), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(new_n207_), .A3(new_n206_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n213_), .A2(new_n217_), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT82), .ZN(new_n225_));
  INV_X1    g024(.A(new_n217_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n226_), .A2(new_n212_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT82), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n228_), .A3(new_n223_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n230_));
  AND2_X1   g029(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n231_));
  AND2_X1   g030(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n233_));
  OAI22_X1  g032(.A1(new_n230_), .A2(new_n231_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n207_), .A2(new_n206_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(KEYINPUT24), .A3(new_n219_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n225_), .A2(new_n229_), .A3(new_n234_), .A4(new_n236_), .ZN(new_n237_));
  AND3_X1   g036(.A1(new_n221_), .A2(KEYINPUT85), .A3(new_n237_), .ZN(new_n238_));
  AOI21_X1  g037(.A(KEYINPUT85), .B1(new_n221_), .B2(new_n237_), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT86), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n221_), .A2(new_n237_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT85), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT86), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n221_), .A2(KEYINPUT85), .A3(new_n237_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n240_), .A2(new_n246_), .A3(KEYINPUT30), .ZN(new_n247_));
  AOI21_X1  g046(.A(KEYINPUT30), .B1(new_n240_), .B2(new_n246_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT87), .ZN(new_n249_));
  NOR3_X1   g048(.A1(new_n247_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT30), .ZN(new_n252_));
  NOR3_X1   g051(.A1(new_n238_), .A2(new_n239_), .A3(KEYINPUT86), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n244_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n252_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n240_), .A2(new_n246_), .A3(KEYINPUT30), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT87), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G15gat), .B(G43gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G71gat), .B(G99gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  AND2_X1   g059(.A1(G227gat), .A2(G233gat), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n260_), .B(new_n261_), .Z(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT31), .B1(new_n257_), .B2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G127gat), .B(G134gat), .ZN(new_n265_));
  INV_X1    g064(.A(G113gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(G120gat), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n249_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT31), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n269_), .A2(new_n270_), .A3(new_n262_), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n264_), .A2(new_n268_), .A3(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n268_), .B1(new_n264_), .B2(new_n271_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n251_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n268_), .ZN(new_n275_));
  NOR3_X1   g074(.A1(new_n257_), .A2(KEYINPUT31), .A3(new_n263_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n270_), .B1(new_n269_), .B2(new_n262_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n275_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n264_), .A2(new_n268_), .A3(new_n271_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(new_n250_), .A3(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n274_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G155gat), .A2(G162gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT1), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT1), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n284_), .A2(G155gat), .A3(G162gat), .ZN(new_n285_));
  OR2_X1    g084(.A1(G155gat), .A2(G162gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n283_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  OR2_X1    g086(.A1(G141gat), .A2(G148gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n287_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(new_n290_), .B(KEYINPUT88), .Z(new_n291_));
  XNOR2_X1  g090(.A(new_n288_), .B(KEYINPUT3), .ZN(new_n292_));
  XOR2_X1   g091(.A(new_n289_), .B(KEYINPUT2), .Z(new_n293_));
  OAI211_X1 g092(.A(new_n286_), .B(new_n282_), .C1(new_n292_), .C2(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT89), .B1(new_n291_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n291_), .A2(KEYINPUT89), .A3(new_n294_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NOR3_X1   g097(.A1(new_n298_), .A2(KEYINPUT93), .A3(KEYINPUT29), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT93), .ZN(new_n300_));
  INV_X1    g099(.A(new_n297_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n301_), .A2(new_n295_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT29), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n300_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n299_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(G204gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(G197gat), .ZN(new_n307_));
  INV_X1    g106(.A(G197gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(G204gat), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT92), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n307_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G211gat), .B(G218gat), .ZN(new_n312_));
  AND3_X1   g111(.A1(new_n311_), .A2(KEYINPUT21), .A3(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(KEYINPUT21), .B1(new_n311_), .B2(new_n312_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n307_), .A2(new_n309_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n315_), .A2(new_n312_), .ZN(new_n316_));
  NOR3_X1   g115(.A1(new_n313_), .A2(new_n314_), .A3(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(G233gat), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT91), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n319_), .A2(G228gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(G228gat), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n318_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n317_), .B(new_n324_), .C1(new_n302_), .C2(new_n303_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n291_), .A2(new_n294_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n317_), .B1(new_n327_), .B2(new_n303_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(new_n323_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n325_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n305_), .A2(new_n330_), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n329_), .B(new_n325_), .C1(new_n299_), .C2(new_n304_), .ZN(new_n332_));
  XOR2_X1   g131(.A(G22gat), .B(G50gat), .Z(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  XOR2_X1   g134(.A(G78gat), .B(G106gat), .Z(new_n336_));
  XOR2_X1   g135(.A(new_n335_), .B(new_n336_), .Z(new_n337_));
  AND3_X1   g136(.A1(new_n331_), .A2(new_n332_), .A3(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n337_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n281_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G225gat), .A2(G233gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT97), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT4), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n268_), .B1(new_n301_), .B2(new_n295_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n327_), .A2(new_n275_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n345_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT4), .B1(new_n298_), .B2(new_n268_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n344_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n346_), .A2(new_n342_), .A3(new_n347_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G1gat), .B(G29gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(G85gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT0), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(G57gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n350_), .A2(new_n351_), .A3(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n356_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G64gat), .B(G92gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G8gat), .B(G36gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n362_), .B(new_n363_), .Z(new_n364_));
  NAND2_X1  g163(.A1(G226gat), .A2(G233gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT19), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n207_), .A2(KEYINPUT22), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n208_), .A2(new_n368_), .A3(new_n206_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n218_), .A2(new_n369_), .A3(new_n219_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n234_), .A2(new_n227_), .A3(new_n223_), .A4(new_n236_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n317_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n243_), .A2(new_n245_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n373_), .B1(new_n374_), .B2(new_n317_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n367_), .B1(new_n375_), .B2(KEYINPUT20), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n311_), .A2(new_n312_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT21), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n316_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n311_), .A2(KEYINPUT21), .A3(new_n312_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n379_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n243_), .A2(new_n382_), .A3(new_n245_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n317_), .A2(new_n372_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n383_), .A2(KEYINPUT20), .A3(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n385_), .A2(new_n366_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n364_), .B1(new_n376_), .B2(new_n386_), .ZN(new_n387_));
  OR2_X1    g186(.A1(new_n387_), .A2(KEYINPUT100), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT27), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n389_), .B1(new_n387_), .B2(KEYINPUT100), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n374_), .A2(new_n317_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT20), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT94), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n393_), .B1(new_n317_), .B2(new_n372_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n382_), .A2(KEYINPUT94), .A3(new_n370_), .A4(new_n371_), .ZN(new_n395_));
  AOI211_X1 g194(.A(new_n392_), .B(new_n366_), .C1(new_n394_), .C2(new_n395_), .ZN(new_n396_));
  AOI22_X1  g195(.A1(new_n385_), .A2(new_n366_), .B1(new_n391_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n364_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  OR2_X1    g198(.A1(new_n399_), .A2(KEYINPUT101), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(KEYINPUT101), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n388_), .A2(new_n390_), .A3(new_n400_), .A4(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n385_), .A2(new_n366_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n391_), .A2(new_n396_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n405_), .A2(KEYINPUT96), .A3(new_n364_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT96), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n407_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n406_), .A2(new_n408_), .A3(new_n399_), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n409_), .A2(KEYINPUT102), .A3(new_n389_), .ZN(new_n410_));
  AOI21_X1  g209(.A(KEYINPUT102), .B1(new_n409_), .B2(new_n389_), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n359_), .B(new_n402_), .C1(new_n410_), .C2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n341_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n340_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n398_), .A2(KEYINPUT32), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n397_), .A2(new_n416_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n376_), .A2(new_n386_), .ZN(new_n418_));
  OAI221_X1 g217(.A(new_n417_), .B1(new_n418_), .B2(new_n416_), .C1(new_n357_), .C2(new_n358_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n342_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT99), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT99), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n422_), .B(new_n342_), .C1(new_n348_), .C2(new_n349_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n346_), .A2(new_n347_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n355_), .B1(new_n424_), .B2(new_n343_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT98), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  OAI211_X1 g226(.A(KEYINPUT98), .B(new_n355_), .C1(new_n424_), .C2(new_n343_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n421_), .A2(new_n423_), .A3(new_n427_), .A4(new_n428_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n429_), .A2(new_n399_), .A3(new_n408_), .A4(new_n406_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n350_), .A2(new_n351_), .A3(new_n356_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT33), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n340_), .B(new_n419_), .C1(new_n430_), .C2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n281_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n415_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT103), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n281_), .B1(new_n414_), .B2(new_n412_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT103), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(new_n439_), .A3(new_n434_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n413_), .B1(new_n437_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G230gat), .A2(G233gat), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NOR3_X1   g243(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT67), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  AND3_X1   g245(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT7), .ZN(new_n450_));
  INV_X1    g249(.A(G99gat), .ZN(new_n451_));
  INV_X1    g250(.A(G106gat), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT67), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n453_), .A2(new_n454_), .A3(new_n443_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n446_), .A2(new_n449_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(G85gat), .ZN(new_n457_));
  INV_X1    g256(.A(G92gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G85gat), .A2(G92gat), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n456_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT68), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n456_), .A2(KEYINPUT68), .A3(new_n461_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(KEYINPUT8), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT64), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n467_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G99gat), .A2(G106gat), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT6), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(KEYINPUT64), .A3(new_n472_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n468_), .A2(new_n473_), .A3(new_n443_), .A4(new_n453_), .ZN(new_n474_));
  XOR2_X1   g273(.A(KEYINPUT65), .B(KEYINPUT8), .Z(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(new_n475_), .A3(new_n461_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT66), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT66), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n474_), .A2(new_n478_), .A3(new_n475_), .A4(new_n461_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n466_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT69), .ZN(new_n482_));
  AND2_X1   g281(.A1(new_n468_), .A2(new_n473_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n451_), .A2(KEYINPUT10), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n451_), .A2(KEYINPUT10), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n452_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n461_), .A2(KEYINPUT9), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n483_), .A2(new_n486_), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT9), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n489_), .A2(G85gat), .A3(G92gat), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n482_), .B1(new_n488_), .B2(new_n491_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n487_), .A2(new_n486_), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n493_), .A2(new_n483_), .A3(KEYINPUT69), .A4(new_n490_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n481_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G57gat), .B(G64gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT11), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G71gat), .B(G78gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n497_), .A2(KEYINPUT11), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n496_), .A2(KEYINPUT12), .A3(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n488_), .A2(new_n491_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n505_), .B1(new_n466_), .B2(new_n480_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(new_n502_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT12), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n508_), .B1(new_n506_), .B2(new_n502_), .ZN(new_n509_));
  AND4_X1   g308(.A1(new_n442_), .A2(new_n504_), .A3(new_n507_), .A4(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n442_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n507_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n506_), .A2(new_n502_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n512_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n511_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G120gat), .B(G148gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT71), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G176gat), .B(G204gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n520_), .B(new_n521_), .Z(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n516_), .A2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n511_), .A2(new_n515_), .A3(new_n522_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  AND2_X1   g325(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n526_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G229gat), .A2(G233gat), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(G50gat), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G29gat), .A2(G36gat), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(G29gat), .A2(G36gat), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT73), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(G43gat), .ZN(new_n539_));
  INV_X1    g338(.A(G29gat), .ZN(new_n540_));
  INV_X1    g339(.A(G36gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT73), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n542_), .A2(new_n543_), .A3(new_n535_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n538_), .A2(new_n539_), .A3(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n539_), .B1(new_n538_), .B2(new_n544_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n534_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n547_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n549_), .A2(G50gat), .A3(new_n545_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G15gat), .B(G22gat), .ZN(new_n553_));
  INV_X1    g352(.A(G1gat), .ZN(new_n554_));
  INV_X1    g353(.A(G8gat), .ZN(new_n555_));
  OAI21_X1  g354(.A(KEYINPUT14), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n553_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G1gat), .B(G8gat), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n557_), .B(new_n558_), .Z(new_n559_));
  NOR2_X1   g358(.A1(new_n552_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n559_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n551_), .A2(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n533_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n563_));
  AND3_X1   g362(.A1(new_n548_), .A2(new_n550_), .A3(KEYINPUT15), .ZN(new_n564_));
  AOI21_X1  g363(.A(KEYINPUT15), .B1(new_n548_), .B2(new_n550_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  OR3_X1    g365(.A1(new_n566_), .A2(KEYINPUT79), .A3(new_n559_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n562_), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT79), .B1(new_n566_), .B2(new_n559_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n567_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n563_), .B1(new_n570_), .B2(new_n533_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G113gat), .B(G141gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT81), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(G169gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(new_n308_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(KEYINPUT80), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n571_), .B(new_n576_), .Z(new_n577_));
  NAND2_X1  g376(.A1(new_n531_), .A2(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n441_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G232gat), .A2(G233gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT34), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT35), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n506_), .A2(KEYINPUT75), .A3(new_n552_), .ZN(new_n585_));
  AOI21_X1  g384(.A(KEYINPUT75), .B1(new_n506_), .B2(new_n552_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  AOI22_X1  g386(.A1(new_n466_), .A2(new_n480_), .B1(new_n492_), .B2(new_n494_), .ZN(new_n588_));
  OAI21_X1  g387(.A(KEYINPUT74), .B1(new_n588_), .B2(new_n566_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n565_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n548_), .A2(new_n550_), .A3(KEYINPUT15), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT74), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n496_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n589_), .A2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n584_), .B1(new_n587_), .B2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n581_), .B(KEYINPUT35), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n597_), .B1(new_n496_), .B2(new_n592_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n598_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT76), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT76), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n598_), .B(new_n601_), .C1(new_n585_), .C2(new_n586_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n596_), .A2(new_n600_), .A3(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT77), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G190gat), .B(G218gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(G134gat), .ZN(new_n606_));
  INV_X1    g405(.A(G162gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT36), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT77), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n596_), .A2(new_n600_), .A3(new_n610_), .A4(new_n602_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n604_), .A2(new_n609_), .A3(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT37), .ZN(new_n613_));
  INV_X1    g412(.A(new_n608_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n614_), .A2(KEYINPUT36), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n596_), .A2(new_n600_), .A3(new_n615_), .A4(new_n602_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n612_), .A2(new_n613_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT78), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n603_), .A2(new_n609_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n616_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n618_), .B1(new_n620_), .B2(KEYINPUT37), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n617_), .A2(new_n621_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n612_), .A2(new_n618_), .A3(new_n613_), .A4(new_n616_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G231gat), .A2(G233gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n559_), .B(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(new_n502_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G127gat), .B(G155gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT16), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(new_n214_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(G211gat), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT17), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n631_), .A2(new_n632_), .ZN(new_n634_));
  OR3_X1    g433(.A1(new_n627_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n627_), .A2(new_n634_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n624_), .A2(new_n637_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n579_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n359_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n639_), .A2(new_n554_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT38), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n612_), .A2(new_n616_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n645_), .A2(new_n637_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n579_), .A2(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G1gat), .B1(new_n647_), .B2(new_n359_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n641_), .A2(new_n642_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n643_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(KEYINPUT104), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT104), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n643_), .A2(new_n652_), .A3(new_n648_), .A4(new_n649_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(G1324gat));
  OR2_X1    g453(.A1(new_n410_), .A2(new_n411_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(new_n402_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n639_), .A2(new_n555_), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n656_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G8gat), .B1(new_n647_), .B2(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n659_), .A2(KEYINPUT39), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(KEYINPUT39), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n657_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT40), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(G1325gat));
  INV_X1    g463(.A(G15gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n639_), .A2(new_n665_), .A3(new_n281_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n413_), .ZN(new_n667_));
  AND4_X1   g466(.A1(new_n439_), .A2(new_n415_), .A3(new_n434_), .A4(new_n435_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n439_), .B1(new_n438_), .B2(new_n434_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n667_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n577_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n671_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n670_), .A2(new_n672_), .A3(new_n281_), .A4(new_n646_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(G15gat), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT105), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT105), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n673_), .A2(new_n676_), .A3(G15gat), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n675_), .A2(KEYINPUT41), .A3(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(KEYINPUT41), .B1(new_n675_), .B2(new_n677_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n666_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT106), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  OAI211_X1 g481(.A(KEYINPUT106), .B(new_n666_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1326gat));
  OAI21_X1  g483(.A(G22gat), .B1(new_n647_), .B2(new_n340_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT42), .ZN(new_n686_));
  INV_X1    g485(.A(G22gat), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n639_), .A2(new_n687_), .A3(new_n414_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(G1327gat));
  INV_X1    g488(.A(new_n637_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n644_), .A2(new_n690_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n579_), .A2(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(G29gat), .B1(new_n692_), .B2(new_n640_), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT107), .B1(new_n578_), .B2(new_n690_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT107), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n672_), .A2(new_n695_), .A3(new_n637_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT109), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n624_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n441_), .A2(KEYINPUT43), .A3(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n704_), .B1(new_n670_), .B2(new_n624_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n701_), .B1(new_n703_), .B2(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT109), .B1(new_n698_), .B2(KEYINPUT108), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(KEYINPUT43), .B1(new_n441_), .B2(new_n702_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n670_), .A2(new_n704_), .A3(new_n624_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n707_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n711_), .A2(new_n712_), .A3(new_n701_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n359_), .B1(new_n708_), .B2(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n693_), .B1(new_n714_), .B2(G29gat), .ZN(G1328gat));
  XNOR2_X1  g514(.A(new_n656_), .B(KEYINPUT110), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n692_), .A2(KEYINPUT45), .A3(new_n541_), .A4(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n579_), .A2(new_n541_), .A3(new_n691_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n719_), .B1(new_n720_), .B2(new_n716_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n718_), .A2(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n658_), .B1(new_n708_), .B2(new_n713_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(new_n723_), .B2(new_n541_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT46), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n722_), .B(KEYINPUT46), .C1(new_n723_), .C2(new_n541_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(G1329gat));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n712_), .B1(new_n711_), .B2(new_n701_), .ZN(new_n730_));
  AOI211_X1 g529(.A(new_n707_), .B(new_n700_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n281_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(G43gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n692_), .A2(new_n539_), .A3(new_n281_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n729_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n734_), .ZN(new_n736_));
  AOI211_X1 g535(.A(KEYINPUT47), .B(new_n736_), .C1(new_n732_), .C2(G43gat), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1330gat));
  NAND2_X1  g537(.A1(new_n414_), .A2(new_n534_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT111), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n692_), .A2(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n340_), .B1(new_n708_), .B2(new_n713_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n741_), .B1(new_n742_), .B2(new_n534_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  OAI211_X1 g544(.A(KEYINPUT112), .B(new_n741_), .C1(new_n742_), .C2(new_n534_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1331gat));
  NOR3_X1   g546(.A1(new_n441_), .A2(new_n577_), .A3(new_n531_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n748_), .A2(new_n638_), .ZN(new_n749_));
  INV_X1    g548(.A(G57gat), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n749_), .A2(new_n750_), .A3(new_n640_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n748_), .A2(new_n646_), .ZN(new_n752_));
  OAI21_X1  g551(.A(G57gat), .B1(new_n752_), .B2(new_n359_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(new_n754_));
  XOR2_X1   g553(.A(new_n754_), .B(KEYINPUT113), .Z(G1332gat));
  OAI21_X1  g554(.A(G64gat), .B1(new_n752_), .B2(new_n716_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT48), .ZN(new_n757_));
  INV_X1    g556(.A(G64gat), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n749_), .A2(new_n758_), .A3(new_n717_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(G1333gat));
  OAI21_X1  g559(.A(G71gat), .B1(new_n752_), .B2(new_n435_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT49), .ZN(new_n762_));
  INV_X1    g561(.A(G71gat), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n749_), .A2(new_n763_), .A3(new_n281_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(G1334gat));
  OAI21_X1  g564(.A(G78gat), .B1(new_n752_), .B2(new_n340_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT50), .ZN(new_n767_));
  INV_X1    g566(.A(G78gat), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n749_), .A2(new_n768_), .A3(new_n414_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1335gat));
  INV_X1    g569(.A(new_n531_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n771_), .A2(new_n671_), .A3(new_n637_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n772_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n774_), .A2(new_n457_), .A3(new_n359_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n748_), .A2(new_n691_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n776_), .B(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n640_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n775_), .B1(new_n779_), .B2(new_n457_), .ZN(G1336gat));
  NOR3_X1   g579(.A1(new_n774_), .A2(new_n458_), .A3(new_n716_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n778_), .A2(new_n656_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n782_), .B2(new_n458_), .ZN(G1337gat));
  AOI21_X1  g582(.A(new_n451_), .B1(new_n773_), .B2(new_n281_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n484_), .A2(new_n485_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n435_), .A2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n784_), .B1(new_n778_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n787_), .B(new_n788_), .ZN(G1338gat));
  INV_X1    g588(.A(KEYINPUT52), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n773_), .A2(new_n414_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(G106gat), .ZN(new_n792_));
  AOI211_X1 g591(.A(KEYINPUT52), .B(new_n452_), .C1(new_n773_), .C2(new_n414_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n776_), .B(KEYINPUT114), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n414_), .A2(new_n452_), .ZN(new_n795_));
  OAI22_X1  g594(.A1(new_n792_), .A2(new_n793_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT53), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n798_));
  OAI221_X1 g597(.A(new_n798_), .B1(new_n794_), .B2(new_n795_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n799_), .ZN(G1339gat));
  NAND3_X1  g599(.A1(new_n504_), .A2(new_n507_), .A3(new_n509_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n512_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n510_), .B1(KEYINPUT55), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n801_), .A2(new_n804_), .A3(new_n512_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n523_), .B1(new_n803_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT56), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT56), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n808_), .B(new_n523_), .C1(new_n803_), .C2(new_n805_), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n807_), .A2(new_n525_), .A3(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n571_), .A2(new_n575_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n567_), .A2(new_n533_), .A3(new_n568_), .A4(new_n569_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n532_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n812_), .A2(new_n575_), .A3(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT116), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT116), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n812_), .A2(new_n816_), .A3(new_n575_), .A4(new_n813_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n811_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n810_), .A2(KEYINPUT117), .A3(KEYINPUT58), .A4(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n807_), .A2(new_n818_), .A3(new_n525_), .A4(new_n809_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT58), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n820_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n822_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n819_), .A2(new_n624_), .A3(new_n823_), .A4(new_n824_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n807_), .A2(new_n577_), .A3(new_n525_), .A4(new_n809_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n818_), .A2(new_n526_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n644_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n828_), .A2(KEYINPUT57), .A3(new_n644_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n825_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n637_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n622_), .A2(new_n671_), .A3(new_n690_), .A4(new_n623_), .ZN(new_n836_));
  OAI211_X1 g635(.A(KEYINPUT115), .B(new_n835_), .C1(new_n836_), .C2(new_n771_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n836_), .ZN(new_n838_));
  OR2_X1    g637(.A1(new_n835_), .A2(KEYINPUT115), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n835_), .A2(KEYINPUT115), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n838_), .A2(new_n531_), .A3(new_n839_), .A4(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n834_), .A2(new_n837_), .A3(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n341_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n844_), .A2(new_n845_), .A3(new_n640_), .A4(new_n658_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n842_), .A2(new_n640_), .A3(new_n843_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT59), .B1(new_n847_), .B2(new_n656_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n577_), .A2(G113gat), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(KEYINPUT119), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT118), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n844_), .A2(new_n640_), .A3(new_n658_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n852_), .B(new_n266_), .C1(new_n853_), .C2(new_n671_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n847_), .A2(new_n671_), .A3(new_n656_), .ZN(new_n855_));
  OAI21_X1  g654(.A(KEYINPUT118), .B1(new_n855_), .B2(G113gat), .ZN(new_n856_));
  AOI22_X1  g655(.A1(new_n849_), .A2(new_n851_), .B1(new_n854_), .B2(new_n856_), .ZN(G1340gat));
  NAND3_X1  g656(.A1(new_n846_), .A2(new_n771_), .A3(new_n848_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(G120gat), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n847_), .A2(new_n656_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT60), .ZN(new_n861_));
  AOI21_X1  g660(.A(G120gat), .B1(new_n771_), .B2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(G120gat), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n860_), .A2(new_n863_), .A3(new_n864_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n865_), .A2(KEYINPUT120), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n865_), .A2(KEYINPUT120), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n859_), .B1(new_n866_), .B2(new_n867_), .ZN(G1341gat));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n869_));
  OAI21_X1  g668(.A(G127gat), .B1(new_n637_), .B2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(G127gat), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(KEYINPUT121), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n846_), .A2(new_n848_), .A3(new_n870_), .A4(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n871_), .B1(new_n853_), .B2(new_n637_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1342gat));
  AOI21_X1  g674(.A(G134gat), .B1(new_n860_), .B2(new_n645_), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n624_), .A2(G134gat), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n876_), .B1(new_n849_), .B2(new_n877_), .ZN(G1343gat));
  XNOR2_X1  g677(.A(KEYINPUT123), .B(G141gat), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n842_), .A2(new_n640_), .A3(new_n414_), .A4(new_n435_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n882_), .B2(new_n717_), .ZN(new_n883_));
  AND3_X1   g682(.A1(new_n828_), .A2(KEYINPUT57), .A3(new_n644_), .ZN(new_n884_));
  AOI21_X1  g683(.A(KEYINPUT57), .B1(new_n828_), .B2(new_n644_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n690_), .B1(new_n886_), .B2(new_n825_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n841_), .A2(new_n837_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n414_), .B(new_n435_), .C1(new_n887_), .C2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n890_), .A2(KEYINPUT122), .A3(new_n640_), .A4(new_n716_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n883_), .A2(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n880_), .B1(new_n892_), .B2(new_n577_), .ZN(new_n893_));
  AOI211_X1 g692(.A(new_n671_), .B(new_n879_), .C1(new_n883_), .C2(new_n891_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1344gat));
  NOR2_X1   g694(.A1(new_n889_), .A2(new_n359_), .ZN(new_n896_));
  AOI21_X1  g695(.A(KEYINPUT122), .B1(new_n896_), .B2(new_n716_), .ZN(new_n897_));
  NOR4_X1   g696(.A1(new_n889_), .A2(new_n881_), .A3(new_n359_), .A4(new_n717_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n771_), .B1(new_n897_), .B2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(G148gat), .ZN(new_n900_));
  INV_X1    g699(.A(G148gat), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n892_), .A2(new_n901_), .A3(new_n771_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n900_), .A2(new_n902_), .ZN(G1345gat));
  XNOR2_X1  g702(.A(KEYINPUT61), .B(G155gat), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n904_), .B1(new_n892_), .B2(new_n690_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n904_), .ZN(new_n906_));
  AOI211_X1 g705(.A(new_n637_), .B(new_n906_), .C1(new_n883_), .C2(new_n891_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n905_), .A2(new_n907_), .ZN(G1346gat));
  AOI21_X1  g707(.A(G162gat), .B1(new_n892_), .B2(new_n645_), .ZN(new_n909_));
  AOI211_X1 g708(.A(new_n607_), .B(new_n702_), .C1(new_n883_), .C2(new_n891_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1347gat));
  NOR2_X1   g710(.A1(new_n716_), .A2(new_n640_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n844_), .A2(new_n577_), .A3(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT62), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n913_), .A2(new_n914_), .A3(G169gat), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n914_), .B1(new_n913_), .B2(G169gat), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n844_), .A2(new_n912_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n577_), .A2(new_n208_), .A3(new_n368_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(KEYINPUT124), .ZN(new_n920_));
  OAI22_X1  g719(.A1(new_n916_), .A2(new_n917_), .B1(new_n918_), .B2(new_n920_), .ZN(G1348gat));
  NOR2_X1   g720(.A1(new_n918_), .A2(new_n531_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(new_n206_), .ZN(G1349gat));
  INV_X1    g722(.A(new_n918_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n231_), .A2(new_n230_), .ZN(new_n926_));
  NAND4_X1  g725(.A1(new_n924_), .A2(new_n925_), .A3(new_n926_), .A4(new_n690_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n844_), .A2(new_n690_), .A3(new_n912_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(new_n214_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n926_), .ZN(new_n930_));
  OAI21_X1  g729(.A(KEYINPUT125), .B1(new_n928_), .B2(new_n930_), .ZN(new_n931_));
  AND3_X1   g730(.A1(new_n927_), .A2(new_n929_), .A3(new_n931_), .ZN(G1350gat));
  OAI21_X1  g731(.A(G190gat), .B1(new_n918_), .B2(new_n702_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n645_), .B1(new_n233_), .B2(new_n232_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n933_), .B1(new_n918_), .B2(new_n934_), .ZN(G1351gat));
  NAND4_X1  g734(.A1(new_n842_), .A2(new_n414_), .A3(new_n435_), .A4(new_n912_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n936_), .A2(new_n671_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(new_n308_), .ZN(G1352gat));
  NOR3_X1   g737(.A1(new_n889_), .A2(new_n640_), .A3(new_n716_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n939_), .A2(new_n306_), .A3(new_n771_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT127), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(new_n942_));
  OAI21_X1  g741(.A(KEYINPUT126), .B1(new_n936_), .B2(new_n531_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT126), .ZN(new_n944_));
  NAND4_X1  g743(.A1(new_n890_), .A2(new_n944_), .A3(new_n771_), .A4(new_n912_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n943_), .A2(new_n945_), .A3(G204gat), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n942_), .A2(new_n946_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n947_), .B1(KEYINPUT127), .B2(new_n946_), .ZN(G1353gat));
  NAND2_X1  g747(.A1(new_n939_), .A2(new_n690_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n950_));
  AND2_X1   g749(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n951_));
  NOR3_X1   g750(.A1(new_n949_), .A2(new_n950_), .A3(new_n951_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n952_), .B1(new_n949_), .B2(new_n950_), .ZN(G1354gat));
  AND3_X1   g752(.A1(new_n939_), .A2(G218gat), .A3(new_n624_), .ZN(new_n954_));
  AOI21_X1  g753(.A(G218gat), .B1(new_n939_), .B2(new_n645_), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n954_), .A2(new_n955_), .ZN(G1355gat));
endmodule


