//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 0 1 1 0 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 0 0 0 0 0 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n933_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_, new_n945_;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n205_), .B(KEYINPUT97), .Z(new_n206_));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n208_), .A2(KEYINPUT23), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n209_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n212_), .A2(KEYINPUT24), .A3(new_n213_), .ZN(new_n214_));
  OR3_X1    g013(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT25), .B(G183gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT26), .B(G190gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n211_), .A2(new_n214_), .A3(new_n215_), .A4(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n207_), .A2(KEYINPUT23), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n210_), .A2(new_n207_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n220_), .B1(new_n221_), .B2(KEYINPUT84), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT84), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n210_), .A2(new_n223_), .A3(new_n207_), .ZN(new_n224_));
  INV_X1    g023(.A(G183gat), .ZN(new_n225_));
  INV_X1    g024(.A(G190gat), .ZN(new_n226_));
  AOI22_X1  g025(.A1(new_n222_), .A2(new_n224_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(G169gat), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n219_), .B1(new_n227_), .B2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT96), .ZN(new_n232_));
  OR2_X1    g031(.A1(G197gat), .A2(G204gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G197gat), .A2(G204gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(KEYINPUT21), .A3(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G211gat), .B(G218gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT90), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n237_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n233_), .A2(new_n234_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT21), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n235_), .A2(new_n236_), .ZN(new_n244_));
  AOI22_X1  g043(.A1(new_n239_), .A2(new_n240_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT96), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n246_), .B(new_n219_), .C1(new_n227_), .C2(new_n230_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n232_), .A2(new_n245_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT20), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n222_), .A2(new_n224_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n214_), .A2(new_n215_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n216_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT26), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n253_), .B1(KEYINPUT82), .B2(G190gat), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n253_), .A2(KEYINPUT82), .A3(G190gat), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n251_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n250_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n225_), .A2(new_n226_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n211_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(new_n229_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n244_), .A2(new_n243_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n240_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n263_), .B1(new_n264_), .B2(new_n238_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n249_), .B1(new_n262_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n248_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G226gat), .A2(G233gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT19), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  AOI22_X1  g069(.A1(new_n250_), .A2(new_n257_), .B1(new_n260_), .B2(new_n229_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n249_), .B1(new_n271_), .B2(new_n245_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n231_), .A2(new_n265_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n269_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n272_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n206_), .B1(new_n270_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n272_), .A2(new_n273_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n269_), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n245_), .B(new_n219_), .C1(new_n227_), .C2(new_n230_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n266_), .A2(new_n274_), .A3(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n278_), .A2(new_n205_), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT27), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n276_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT27), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n262_), .A2(new_n265_), .ZN(new_n285_));
  AND4_X1   g084(.A1(KEYINPUT20), .A2(new_n285_), .A3(new_n274_), .A4(new_n279_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n274_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n205_), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n286_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n205_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n284_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT98), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n288_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n281_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT98), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(new_n295_), .A3(new_n284_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n283_), .B1(new_n292_), .B2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G1gat), .B(G29gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT94), .B(G85gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT0), .B(G57gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G225gat), .A2(G233gat), .ZN(new_n303_));
  XOR2_X1   g102(.A(G127gat), .B(G134gat), .Z(new_n304_));
  XOR2_X1   g103(.A(G113gat), .B(G120gat), .Z(new_n305_));
  XOR2_X1   g104(.A(new_n304_), .B(new_n305_), .Z(new_n306_));
  NOR2_X1   g105(.A1(G155gat), .A2(G162gat), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NOR3_X1   g109(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT89), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G141gat), .A2(G148gat), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT2), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n316_), .A2(new_n317_), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n310_), .B1(new_n313_), .B2(new_n320_), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n309_), .A2(KEYINPUT1), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n309_), .A2(KEYINPUT1), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n322_), .A2(new_n308_), .A3(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(G141gat), .A2(G148gat), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n324_), .A2(new_n326_), .A3(new_n314_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n306_), .B1(new_n321_), .B2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n311_), .B(KEYINPUT89), .ZN(new_n330_));
  OAI211_X1 g129(.A(new_n309_), .B(new_n308_), .C1(new_n330_), .C2(new_n319_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n304_), .B(new_n305_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n331_), .A2(new_n332_), .A3(new_n327_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n329_), .A2(new_n333_), .A3(KEYINPUT4), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n331_), .A2(new_n327_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT4), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(new_n336_), .A3(new_n306_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n303_), .B1(new_n334_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n303_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n339_), .B1(new_n329_), .B2(new_n333_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n302_), .B1(new_n338_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NOR3_X1   g141(.A1(new_n338_), .A2(new_n302_), .A3(new_n340_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n332_), .B(KEYINPUT31), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G227gat), .A2(G233gat), .ZN(new_n346_));
  INV_X1    g145(.A(G71gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(G99gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n262_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G15gat), .B(G43gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT85), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT30), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n350_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n271_), .B(new_n349_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n353_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(KEYINPUT86), .B1(new_n354_), .B2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n345_), .B1(new_n358_), .B2(KEYINPUT87), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n345_), .A2(KEYINPUT87), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n354_), .B(new_n357_), .C1(KEYINPUT86), .C2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT29), .B1(new_n321_), .B2(new_n328_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n245_), .B1(new_n364_), .B2(KEYINPUT92), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT29), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n366_), .B1(new_n331_), .B2(new_n327_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT92), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n365_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(G228gat), .ZN(new_n371_));
  INV_X1    g170(.A(G233gat), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n370_), .A2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G78gat), .B(G106gat), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT91), .ZN(new_n377_));
  INV_X1    g176(.A(new_n373_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n265_), .A2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n377_), .B1(new_n379_), .B2(new_n367_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n364_), .A2(KEYINPUT91), .A3(new_n265_), .A4(new_n378_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n374_), .A2(new_n376_), .A3(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT93), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n335_), .A2(KEYINPUT29), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G22gat), .B(G50gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT28), .ZN(new_n387_));
  XOR2_X1   g186(.A(new_n385_), .B(new_n387_), .Z(new_n388_));
  AND2_X1   g187(.A1(new_n380_), .A2(new_n381_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n378_), .B1(new_n365_), .B2(new_n369_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n375_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n384_), .A2(new_n388_), .B1(new_n391_), .B2(new_n383_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT93), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n391_), .A2(new_n383_), .A3(new_n393_), .A4(new_n388_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n392_), .A2(new_n395_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n297_), .A2(new_n344_), .A3(new_n363_), .A4(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n344_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n384_), .A2(new_n388_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n391_), .A2(new_n383_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n398_), .B1(new_n401_), .B2(new_n394_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n329_), .A2(new_n333_), .A3(new_n339_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n302_), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n334_), .A2(new_n303_), .A3(new_n337_), .ZN(new_n406_));
  AOI21_X1  g205(.A(KEYINPUT95), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n405_), .A2(new_n406_), .A3(KEYINPUT95), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n293_), .B(new_n281_), .C1(new_n407_), .C2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT33), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n341_), .A2(new_n410_), .ZN(new_n411_));
  OAI211_X1 g210(.A(KEYINPUT33), .B(new_n302_), .C1(new_n338_), .C2(new_n340_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n205_), .A2(KEYINPUT32), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n278_), .A2(new_n280_), .A3(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n415_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n414_), .B1(new_n270_), .B2(new_n275_), .ZN(new_n417_));
  OAI22_X1  g216(.A1(new_n409_), .A2(new_n413_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n297_), .A2(new_n402_), .B1(new_n396_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT88), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n362_), .B(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n397_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G1gat), .B(G8gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT75), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G15gat), .B(G22gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G1gat), .A2(G8gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT14), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n426_), .A2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n425_), .A2(new_n429_), .ZN(new_n430_));
  OR2_X1    g229(.A1(new_n424_), .A2(KEYINPUT75), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n424_), .A2(KEYINPUT75), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n431_), .A2(new_n428_), .A3(new_n426_), .A4(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n430_), .A2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G29gat), .B(G36gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G43gat), .B(G50gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n434_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT80), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT81), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n438_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n440_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n443_));
  OAI22_X1  g242(.A1(new_n442_), .A2(new_n443_), .B1(new_n434_), .B2(new_n437_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n443_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n434_), .A2(new_n437_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n445_), .A2(new_n446_), .A3(new_n441_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G229gat), .A2(G233gat), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n444_), .A2(new_n447_), .A3(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(new_n437_), .B(KEYINPUT15), .Z(new_n451_));
  OR2_X1    g250(.A1(new_n451_), .A2(new_n434_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n452_), .A2(new_n448_), .A3(new_n438_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G113gat), .B(G141gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G169gat), .B(G197gat), .ZN(new_n455_));
  XOR2_X1   g254(.A(new_n454_), .B(new_n455_), .Z(new_n456_));
  AND3_X1   g255(.A1(new_n450_), .A2(new_n453_), .A3(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n456_), .B1(new_n450_), .B2(new_n453_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n423_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT69), .ZN(new_n461_));
  INV_X1    g260(.A(G106gat), .ZN(new_n462_));
  AND2_X1   g261(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n463_));
  NOR2_X1   g262(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT64), .ZN(new_n465_));
  NOR3_X1   g264(.A1(new_n463_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  OR2_X1    g265(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n468_));
  AOI21_X1  g267(.A(KEYINPUT64), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n462_), .B1(new_n466_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G85gat), .A2(G92gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(G85gat), .A2(G92gat), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT9), .ZN(new_n474_));
  NOR3_X1   g273(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G99gat), .A2(G106gat), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT6), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n474_), .A2(G85gat), .A3(G92gat), .ZN(new_n479_));
  NAND3_X1  g278(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n475_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n470_), .A2(KEYINPUT65), .A3(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT65), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n467_), .A2(KEYINPUT64), .A3(new_n468_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n465_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n486_));
  AOI21_X1  g285(.A(G106gat), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  AND3_X1   g286(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n488_));
  AOI21_X1  g287(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(G85gat), .ZN(new_n491_));
  INV_X1    g290(.A(G92gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n493_), .A2(KEYINPUT9), .A3(new_n471_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n490_), .A2(new_n494_), .A3(new_n479_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n484_), .B1(new_n487_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n483_), .A2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G57gat), .B(G64gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT11), .ZN(new_n499_));
  XOR2_X1   g298(.A(G71gat), .B(G78gat), .Z(new_n500_));
  OR2_X1    g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n498_), .A2(KEYINPUT11), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n499_), .A2(new_n500_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n501_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT8), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n477_), .A2(KEYINPUT67), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT67), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT6), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n509_), .A2(G99gat), .A3(G106gat), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT7), .ZN(new_n511_));
  INV_X1    g310(.A(G99gat), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n512_), .A3(new_n462_), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n506_), .A2(new_n508_), .A3(new_n476_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n510_), .A2(new_n513_), .A3(new_n514_), .A4(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n472_), .A2(new_n473_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n505_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n513_), .A2(new_n478_), .A3(new_n480_), .A4(new_n514_), .ZN(new_n519_));
  NOR3_X1   g318(.A1(new_n472_), .A2(new_n473_), .A3(KEYINPUT8), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT66), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n519_), .A2(KEYINPUT66), .A3(new_n520_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n497_), .B(new_n504_), .C1(new_n518_), .C2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G230gat), .A2(G233gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n515_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n476_), .B1(new_n506_), .B2(new_n508_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n517_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT8), .ZN(new_n532_));
  AND3_X1   g331(.A1(new_n519_), .A2(KEYINPUT66), .A3(new_n520_), .ZN(new_n533_));
  AOI21_X1  g332(.A(KEYINPUT66), .B1(new_n519_), .B2(new_n520_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  AOI22_X1  g334(.A1(new_n532_), .A2(new_n535_), .B1(new_n496_), .B2(new_n483_), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT12), .B1(new_n536_), .B2(new_n504_), .ZN(new_n537_));
  AOI21_X1  g336(.A(KEYINPUT65), .B1(new_n470_), .B2(new_n482_), .ZN(new_n538_));
  NOR3_X1   g337(.A1(new_n487_), .A2(new_n495_), .A3(new_n484_), .ZN(new_n539_));
  OAI22_X1  g338(.A1(new_n518_), .A2(new_n525_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT12), .ZN(new_n541_));
  INV_X1    g340(.A(new_n504_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n540_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n528_), .B1(new_n537_), .B2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n540_), .A2(new_n542_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(new_n526_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n527_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(KEYINPUT68), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT68), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n546_), .A2(new_n550_), .A3(new_n547_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n544_), .B1(new_n549_), .B2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G120gat), .B(G148gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT5), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G176gat), .B(G204gat), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n554_), .B(new_n555_), .Z(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n461_), .B1(new_n552_), .B2(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n547_), .B1(new_n536_), .B2(new_n504_), .ZN(new_n559_));
  NOR3_X1   g358(.A1(new_n536_), .A2(KEYINPUT12), .A3(new_n504_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n541_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n559_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n550_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n563_));
  AOI211_X1 g362(.A(KEYINPUT68), .B(new_n527_), .C1(new_n545_), .C2(new_n526_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n562_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n565_), .A2(KEYINPUT69), .A3(new_n556_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n558_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n552_), .A2(KEYINPUT70), .A3(new_n557_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT70), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n569_), .B1(new_n565_), .B2(new_n556_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n567_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT13), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n567_), .A2(new_n571_), .A3(KEYINPUT13), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n536_), .A2(new_n437_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n577_), .B1(new_n451_), .B2(new_n536_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G232gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT34), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n580_), .A2(KEYINPUT35), .ZN(new_n581_));
  AOI21_X1  g380(.A(KEYINPUT71), .B1(new_n536_), .B2(new_n437_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(KEYINPUT35), .ZN(new_n583_));
  OAI22_X1  g382(.A1(new_n578_), .A2(new_n581_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n451_), .A2(new_n536_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n583_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n585_), .A2(KEYINPUT71), .A3(new_n577_), .A4(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(G190gat), .B(G218gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT72), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G134gat), .B(G162gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT36), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n584_), .A2(new_n587_), .A3(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT73), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n584_), .A2(new_n587_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n591_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n596_), .A2(KEYINPUT36), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT37), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT73), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n584_), .A2(new_n600_), .A3(new_n587_), .A4(new_n592_), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n594_), .A2(new_n598_), .A3(new_n599_), .A4(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT74), .ZN(new_n603_));
  INV_X1    g402(.A(new_n593_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n597_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n605_), .B1(new_n584_), .B2(new_n587_), .ZN(new_n606_));
  OAI21_X1  g405(.A(KEYINPUT37), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  AND3_X1   g406(.A1(new_n602_), .A2(new_n603_), .A3(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n603_), .B1(new_n602_), .B2(new_n607_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n504_), .B(KEYINPUT76), .Z(new_n611_));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n434_), .B(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n611_), .B(new_n613_), .ZN(new_n614_));
  XOR2_X1   g413(.A(G127gat), .B(G155gat), .Z(new_n615_));
  XNOR2_X1  g414(.A(G183gat), .B(G211gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n619_), .B(KEYINPUT17), .Z(new_n620_));
  NAND2_X1  g419(.A1(new_n614_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT78), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n619_), .A2(KEYINPUT17), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n614_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT78), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n614_), .A2(new_n625_), .A3(new_n620_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n622_), .A2(new_n624_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT79), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n576_), .A2(new_n610_), .A3(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n460_), .A2(new_n630_), .ZN(new_n631_));
  NOR3_X1   g430(.A1(new_n631_), .A2(G1gat), .A3(new_n344_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n574_), .A2(new_n575_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n629_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n459_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n635_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n638_), .A2(KEYINPUT100), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(KEYINPUT100), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n594_), .A2(new_n601_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(new_n598_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT101), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n423_), .A2(new_n644_), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n639_), .A2(new_n640_), .A3(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(new_n398_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(G1gat), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n634_), .A2(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT102), .ZN(G1324gat));
  INV_X1    g449(.A(KEYINPUT39), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n295_), .B1(new_n294_), .B2(new_n284_), .ZN(new_n652_));
  AOI211_X1 g451(.A(KEYINPUT98), .B(KEYINPUT27), .C1(new_n293_), .C2(new_n281_), .ZN(new_n653_));
  OAI22_X1  g452(.A1(new_n652_), .A2(new_n653_), .B1(new_n276_), .B2(new_n282_), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n639_), .A2(new_n640_), .A3(new_n654_), .A4(new_n645_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n651_), .B1(new_n655_), .B2(G8gat), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n655_), .A2(new_n651_), .A3(G8gat), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  OR3_X1    g458(.A1(new_n631_), .A2(G8gat), .A3(new_n297_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n659_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n661_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1325gat));
  INV_X1    g464(.A(G15gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(new_n646_), .B2(new_n421_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT41), .ZN(new_n668_));
  INV_X1    g467(.A(new_n631_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n666_), .A3(new_n421_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(G1326gat));
  OR3_X1    g470(.A1(new_n631_), .A2(G22gat), .A3(new_n396_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n396_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n646_), .A2(new_n673_), .ZN(new_n674_));
  XOR2_X1   g473(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n675_));
  AND3_X1   g474(.A1(new_n674_), .A2(G22gat), .A3(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n674_), .B2(G22gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n672_), .B1(new_n676_), .B2(new_n677_), .ZN(G1327gat));
  NOR3_X1   g477(.A1(new_n576_), .A2(new_n636_), .A3(new_n642_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n460_), .A2(new_n679_), .ZN(new_n680_));
  OR3_X1    g479(.A1(new_n680_), .A2(G29gat), .A3(new_n344_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n602_), .A2(new_n607_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT74), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT43), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n602_), .A2(new_n603_), .A3(new_n607_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n684_), .A2(new_n685_), .A3(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n396_), .A2(new_n418_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n344_), .B1(new_n392_), .B2(new_n395_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(new_n654_), .B2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n362_), .B(KEYINPUT88), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n687_), .B1(new_n692_), .B2(new_n397_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT106), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n694_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n684_), .A2(KEYINPUT106), .A3(new_n686_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(new_n422_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n693_), .B1(new_n698_), .B2(KEYINPUT43), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n574_), .A2(new_n629_), .A3(new_n637_), .A4(new_n575_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT105), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n700_), .B(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n682_), .B1(new_n699_), .B2(new_n702_), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n635_), .A2(new_n701_), .A3(new_n629_), .A4(new_n637_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n700_), .A2(KEYINPUT105), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n685_), .B1(new_n697_), .B2(new_n422_), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n706_), .B(KEYINPUT44), .C1(new_n707_), .C2(new_n693_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n703_), .A2(new_n398_), .A3(new_n708_), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n709_), .A2(KEYINPUT107), .A3(G29gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(KEYINPUT107), .B1(new_n709_), .B2(G29gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n681_), .B1(new_n710_), .B2(new_n711_), .ZN(G1328gat));
  NOR3_X1   g511(.A1(new_n680_), .A2(G36gat), .A3(new_n297_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT45), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n713_), .B(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n703_), .A2(new_n654_), .A3(new_n708_), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n716_), .A2(KEYINPUT108), .A3(G36gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(KEYINPUT108), .B1(new_n716_), .B2(G36gat), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n715_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT46), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n715_), .B(KEYINPUT46), .C1(new_n717_), .C2(new_n718_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1329gat));
  NAND4_X1  g522(.A1(new_n703_), .A2(new_n708_), .A3(G43gat), .A4(new_n363_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n680_), .A2(new_n691_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(G43gat), .B2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g526(.A1(new_n703_), .A2(new_n673_), .A3(new_n708_), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n728_), .A2(KEYINPUT109), .A3(G50gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(KEYINPUT109), .B1(new_n728_), .B2(G50gat), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n396_), .A2(G50gat), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT110), .ZN(new_n732_));
  OAI22_X1  g531(.A1(new_n729_), .A2(new_n730_), .B1(new_n680_), .B2(new_n732_), .ZN(G1331gat));
  NOR3_X1   g532(.A1(new_n423_), .A2(new_n637_), .A3(new_n635_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n610_), .A2(new_n629_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(G57gat), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n736_), .A2(new_n737_), .A3(new_n398_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n635_), .A2(new_n637_), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n645_), .A2(new_n636_), .A3(new_n739_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n740_), .A2(new_n398_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n738_), .B1(new_n741_), .B2(new_n737_), .ZN(G1332gat));
  INV_X1    g541(.A(G64gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n740_), .B2(new_n654_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT48), .Z(new_n745_));
  NOR2_X1   g544(.A1(new_n297_), .A2(G64gat), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT111), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n736_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n745_), .A2(new_n748_), .ZN(G1333gat));
  AOI21_X1  g548(.A(new_n347_), .B1(new_n740_), .B2(new_n421_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT49), .Z(new_n751_));
  NAND3_X1  g550(.A1(new_n736_), .A2(new_n347_), .A3(new_n421_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1334gat));
  INV_X1    g552(.A(G78gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n754_), .B1(new_n740_), .B2(new_n673_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT50), .Z(new_n756_));
  NAND3_X1  g555(.A1(new_n736_), .A2(new_n754_), .A3(new_n673_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(G1335gat));
  NAND2_X1  g557(.A1(new_n739_), .A2(new_n629_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n699_), .A2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(G85gat), .B1(new_n761_), .B2(new_n344_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n642_), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n734_), .A2(new_n629_), .A3(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n764_), .A2(new_n491_), .A3(new_n398_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n762_), .A2(new_n765_), .ZN(G1336gat));
  NAND3_X1  g565(.A1(new_n764_), .A2(new_n492_), .A3(new_n654_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n760_), .A2(new_n654_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n767_), .B1(new_n769_), .B2(new_n492_), .ZN(G1337gat));
  NAND2_X1  g569(.A1(new_n760_), .A2(new_n421_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n362_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n772_));
  AOI22_X1  g571(.A1(new_n771_), .A2(G99gat), .B1(new_n764_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n774_), .A2(KEYINPUT113), .A3(KEYINPUT51), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT113), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n773_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT112), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n779_), .B1(new_n774_), .B2(KEYINPUT51), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n773_), .A2(KEYINPUT112), .A3(new_n777_), .ZN(new_n781_));
  OAI22_X1  g580(.A1(new_n775_), .A2(new_n778_), .B1(new_n780_), .B2(new_n781_), .ZN(G1338gat));
  INV_X1    g581(.A(new_n759_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n783_), .B(new_n673_), .C1(new_n707_), .C2(new_n693_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(G106gat), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT114), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n784_), .A2(new_n787_), .A3(G106gat), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n786_), .A2(KEYINPUT52), .A3(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n787_), .B1(new_n784_), .B2(G106gat), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n396_), .A2(G106gat), .ZN(new_n792_));
  AOI22_X1  g591(.A1(new_n790_), .A2(new_n791_), .B1(new_n764_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n789_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT53), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n789_), .A2(new_n793_), .A3(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(G1339gat));
  INV_X1    g597(.A(KEYINPUT119), .ZN(new_n799_));
  XOR2_X1   g598(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n800_));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n526_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n802_));
  AOI22_X1  g601(.A1(new_n801_), .A2(new_n562_), .B1(new_n802_), .B2(new_n547_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n544_), .A2(KEYINPUT55), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n557_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(KEYINPUT115), .B1(new_n805_), .B2(KEYINPUT56), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n802_), .A2(new_n547_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n562_), .A2(new_n801_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n808_), .A3(new_n804_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n556_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT56), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n810_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n809_), .A2(KEYINPUT56), .A3(new_n556_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n809_), .A2(KEYINPUT116), .A3(KEYINPUT56), .A4(new_n556_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n806_), .A2(new_n813_), .A3(new_n816_), .A4(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT117), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n459_), .B1(new_n570_), .B2(new_n568_), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n818_), .A2(new_n819_), .A3(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n819_), .B1(new_n818_), .B2(new_n820_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n444_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n448_), .B1(new_n434_), .B2(new_n437_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n456_), .B1(new_n452_), .B2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n457_), .B1(new_n823_), .B2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n572_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n821_), .A2(new_n822_), .A3(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n800_), .B1(new_n829_), .B2(new_n763_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n810_), .A2(new_n812_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n814_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(new_n571_), .A3(new_n826_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT58), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n832_), .A2(KEYINPUT58), .A3(new_n571_), .A4(new_n826_), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n835_), .A2(new_n836_), .A3(new_n610_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n818_), .A2(new_n820_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT117), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n818_), .A2(new_n819_), .A3(new_n820_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n840_), .A3(new_n827_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n642_), .A2(KEYINPUT57), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n837_), .B1(new_n841_), .B2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n636_), .B1(new_n830_), .B2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n735_), .A2(new_n459_), .A3(new_n635_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n846_), .B(new_n847_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n845_), .A2(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n654_), .A2(new_n673_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n850_), .A2(new_n398_), .A3(new_n363_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n799_), .B1(new_n849_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(G113gat), .ZN(new_n853_));
  INV_X1    g652(.A(new_n837_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n829_), .B2(new_n842_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n800_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(new_n841_), .B2(new_n642_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n629_), .B1(new_n855_), .B2(new_n857_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n846_), .B(KEYINPUT54), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n851_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(KEYINPUT119), .A3(new_n861_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n852_), .A2(new_n853_), .A3(new_n637_), .A4(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT59), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n864_), .B1(new_n849_), .B2(new_n851_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n860_), .A2(KEYINPUT59), .A3(new_n861_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n459_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n863_), .B1(new_n867_), .B2(new_n853_), .ZN(G1340gat));
  INV_X1    g667(.A(G120gat), .ZN(new_n869_));
  OR2_X1    g668(.A1(new_n869_), .A2(KEYINPUT60), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n635_), .B2(KEYINPUT60), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n852_), .A2(new_n862_), .A3(new_n870_), .A4(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n635_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(new_n869_), .ZN(G1341gat));
  NAND3_X1  g673(.A1(new_n852_), .A2(new_n636_), .A3(new_n862_), .ZN(new_n875_));
  INV_X1    g674(.A(G127gat), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n865_), .A2(new_n866_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n629_), .A2(new_n876_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(KEYINPUT120), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n875_), .A2(new_n876_), .B1(new_n877_), .B2(new_n879_), .ZN(G1342gat));
  NAND3_X1  g679(.A1(new_n852_), .A2(new_n644_), .A3(new_n862_), .ZN(new_n881_));
  INV_X1    g680(.A(G134gat), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n610_), .A2(G134gat), .ZN(new_n883_));
  XOR2_X1   g682(.A(new_n883_), .B(KEYINPUT121), .Z(new_n884_));
  AOI22_X1  g683(.A1(new_n881_), .A2(new_n882_), .B1(new_n877_), .B2(new_n884_), .ZN(G1343gat));
  NAND2_X1  g684(.A1(new_n691_), .A2(new_n673_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n297_), .A2(new_n398_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n887_), .B(new_n889_), .C1(new_n845_), .C2(new_n848_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n637_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n576_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n896_), .B1(new_n890_), .B2(new_n629_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n886_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n898_));
  NAND4_X1  g697(.A1(new_n898_), .A2(KEYINPUT122), .A3(new_n636_), .A4(new_n889_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(KEYINPUT61), .B(G155gat), .ZN(new_n900_));
  AND3_X1   g699(.A1(new_n897_), .A2(new_n899_), .A3(new_n900_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n900_), .B1(new_n897_), .B2(new_n899_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1346gat));
  AOI21_X1  g702(.A(G162gat), .B1(new_n891_), .B2(new_n644_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n697_), .A2(G162gat), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n904_), .B1(new_n891_), .B2(new_n905_), .ZN(G1347gat));
  AND2_X1   g705(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n297_), .A2(new_n398_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n421_), .A2(new_n908_), .A3(new_n396_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n860_), .A2(new_n910_), .ZN(new_n911_));
  OAI211_X1 g710(.A(G169gat), .B(new_n907_), .C1(new_n911_), .C2(new_n459_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(KEYINPUT22), .B(G169gat), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n637_), .A2(new_n913_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(KEYINPUT124), .ZN(new_n915_));
  INV_X1    g714(.A(G169gat), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n849_), .A2(new_n909_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(new_n637_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n919_));
  OAI221_X1 g718(.A(new_n912_), .B1(new_n911_), .B2(new_n915_), .C1(new_n918_), .C2(new_n919_), .ZN(G1348gat));
  NAND2_X1  g719(.A1(new_n917_), .A2(new_n576_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g721(.A1(new_n860_), .A2(new_n636_), .A3(new_n910_), .ZN(new_n923_));
  OR3_X1    g722(.A1(new_n923_), .A2(KEYINPUT125), .A3(new_n216_), .ZN(new_n924_));
  OAI21_X1  g723(.A(KEYINPUT125), .B1(new_n923_), .B2(new_n216_), .ZN(new_n925_));
  AND2_X1   g724(.A1(new_n923_), .A2(new_n225_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n924_), .B1(new_n925_), .B2(new_n926_), .ZN(G1350gat));
  NAND3_X1  g726(.A1(new_n917_), .A2(new_n644_), .A3(new_n217_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n860_), .A2(new_n610_), .A3(new_n910_), .ZN(new_n929_));
  AND3_X1   g728(.A1(new_n929_), .A2(KEYINPUT126), .A3(G190gat), .ZN(new_n930_));
  AOI21_X1  g729(.A(KEYINPUT126), .B1(new_n929_), .B2(G190gat), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n928_), .B1(new_n930_), .B2(new_n931_), .ZN(G1351gat));
  NAND3_X1  g731(.A1(new_n898_), .A2(new_n637_), .A3(new_n908_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g733(.A1(new_n898_), .A2(new_n576_), .A3(new_n908_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g735(.A(new_n629_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n898_), .A2(new_n908_), .A3(new_n937_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(KEYINPUT127), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n938_), .B(new_n940_), .ZN(G1354gat));
  NAND2_X1  g740(.A1(new_n898_), .A2(new_n908_), .ZN(new_n942_));
  INV_X1    g741(.A(new_n610_), .ZN(new_n943_));
  OAI21_X1  g742(.A(G218gat), .B1(new_n942_), .B2(new_n943_), .ZN(new_n944_));
  OR2_X1    g743(.A1(new_n643_), .A2(G218gat), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n944_), .B1(new_n942_), .B2(new_n945_), .ZN(G1355gat));
endmodule


