//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 0 0 1 0 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n765_, new_n766_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n782_, new_n783_, new_n784_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n803_, new_n804_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n919_, new_n921_, new_n922_, new_n924_, new_n925_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n942_, new_n944_, new_n945_, new_n946_, new_n947_, new_n949_,
    new_n950_, new_n952_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n959_, new_n960_;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G141gat), .A2(G148gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT90), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT1), .ZN(new_n210_));
  OAI211_X1 g009(.A(new_n205_), .B(new_n206_), .C1(new_n208_), .C2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT90), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n207_), .B(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n204_), .B(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n206_), .B(new_n216_), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n213_), .B(new_n209_), .C1(new_n215_), .C2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n211_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT29), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G197gat), .B(G204gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G211gat), .B(G218gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT21), .ZN(new_n223_));
  OR3_X1    g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n221_), .A2(new_n223_), .ZN(new_n225_));
  INV_X1    g024(.A(G197gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n226_), .A2(G204gat), .ZN(new_n227_));
  INV_X1    g026(.A(G204gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n228_), .A2(G197gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT21), .B1(new_n227_), .B2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n225_), .A2(new_n230_), .A3(new_n222_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n224_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n220_), .A2(KEYINPUT92), .A3(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT29), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n235_), .B1(new_n211_), .B2(new_n218_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT91), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n236_), .A2(new_n237_), .A3(new_n232_), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n203_), .B(new_n234_), .C1(new_n238_), .C2(KEYINPUT92), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n220_), .A2(KEYINPUT91), .A3(new_n233_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT92), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n240_), .A2(new_n241_), .A3(new_n202_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n239_), .A2(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G78gat), .B(G106gat), .Z(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n244_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n239_), .A2(new_n242_), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n219_), .A2(KEYINPUT29), .ZN(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT28), .B(G22gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(G50gat), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n249_), .B(new_n251_), .Z(new_n252_));
  AOI21_X1  g051(.A(new_n246_), .B1(new_n239_), .B2(new_n242_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n252_), .B1(new_n253_), .B2(KEYINPUT93), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n248_), .A2(new_n254_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n245_), .A2(KEYINPUT93), .A3(new_n247_), .A4(new_n252_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT88), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G169gat), .A2(G176gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT87), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT87), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(G169gat), .A3(G176gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT24), .ZN(new_n267_));
  INV_X1    g066(.A(G169gat), .ZN(new_n268_));
  INV_X1    g067(.A(G176gat), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n267_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G183gat), .A2(G190gat), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT23), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n274_));
  AND3_X1   g073(.A1(new_n270_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT86), .ZN(new_n276_));
  INV_X1    g075(.A(G190gat), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT26), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(KEYINPUT85), .A2(G183gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(KEYINPUT25), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT25), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n281_), .A2(KEYINPUT85), .A3(G183gat), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT26), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n283_), .A2(KEYINPUT86), .A3(G190gat), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n278_), .A2(new_n280_), .A3(new_n282_), .A4(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n266_), .A2(new_n275_), .A3(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT30), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT22), .B(G169gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n269_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n273_), .B(new_n274_), .C1(G183gat), .C2(G190gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n289_), .A2(new_n290_), .A3(new_n263_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n286_), .A2(new_n287_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n287_), .B1(new_n286_), .B2(new_n291_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n258_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT31), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT31), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n258_), .B(new_n297_), .C1(new_n293_), .C2(new_n294_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n294_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n299_), .A2(KEYINPUT88), .A3(new_n292_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT89), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G71gat), .B(G99gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G15gat), .B(G43gat), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n302_), .B(new_n303_), .Z(new_n304_));
  NAND2_X1  g103(.A1(G227gat), .A2(G233gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  AND3_X1   g105(.A1(new_n300_), .A2(new_n301_), .A3(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n301_), .B1(new_n300_), .B2(new_n306_), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n296_), .B(new_n298_), .C1(new_n307_), .C2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n308_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n300_), .A2(new_n301_), .A3(new_n306_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n296_), .A2(new_n298_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n310_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(G120gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G127gat), .B(G134gat), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n315_), .A2(G113gat), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n315_), .A2(G113gat), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n314_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n315_), .A2(G113gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n315_), .A2(G113gat), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(G120gat), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n318_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  AND3_X1   g122(.A1(new_n309_), .A2(new_n313_), .A3(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n323_), .B1(new_n309_), .B2(new_n313_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n257_), .A2(new_n326_), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n255_), .B(new_n256_), .C1(new_n324_), .C2(new_n325_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n322_), .A2(new_n219_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n211_), .A2(new_n318_), .A3(new_n321_), .A4(new_n218_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n330_), .A2(KEYINPUT4), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G225gat), .A2(G233gat), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT4), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n322_), .A2(new_n219_), .A3(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n332_), .A2(new_n334_), .A3(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n330_), .A2(new_n333_), .A3(new_n331_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT99), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n337_), .A2(new_n340_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n332_), .A2(new_n339_), .A3(new_n334_), .A4(new_n336_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G1gat), .B(G29gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(G85gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT0), .ZN(new_n346_));
  INV_X1    g145(.A(G57gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n343_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n341_), .A2(new_n348_), .A3(new_n342_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT27), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n232_), .A2(new_n286_), .A3(new_n291_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n275_), .B(KEYINPUT95), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n265_), .A2(new_n259_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT25), .B(G183gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT26), .B(G190gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n356_), .A2(KEYINPUT96), .A3(new_n357_), .A4(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n275_), .A2(KEYINPUT95), .ZN(new_n362_));
  AND4_X1   g161(.A1(KEYINPUT95), .A2(new_n270_), .A3(new_n273_), .A4(new_n274_), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n357_), .B(new_n360_), .C1(new_n362_), .C2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT96), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n263_), .A2(KEYINPUT97), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT97), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n260_), .A2(new_n262_), .A3(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n367_), .A2(new_n289_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(KEYINPUT98), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT98), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n367_), .A2(new_n372_), .A3(new_n289_), .A4(new_n369_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  AOI22_X1  g173(.A1(new_n361_), .A2(new_n366_), .B1(new_n290_), .B2(new_n374_), .ZN(new_n375_));
  OAI211_X1 g174(.A(KEYINPUT20), .B(new_n355_), .C1(new_n375_), .C2(new_n232_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G226gat), .A2(G233gat), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n377_), .B(KEYINPUT94), .Z(new_n378_));
  XOR2_X1   g177(.A(new_n378_), .B(KEYINPUT19), .Z(new_n379_));
  AOI21_X1  g178(.A(new_n379_), .B1(new_n375_), .B2(new_n232_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT20), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n286_), .A2(new_n291_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n381_), .B1(new_n233_), .B2(new_n382_), .ZN(new_n383_));
  AOI22_X1  g182(.A1(new_n376_), .A2(new_n379_), .B1(new_n380_), .B2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G8gat), .B(G36gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT18), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(G64gat), .ZN(new_n387_));
  INV_X1    g186(.A(G92gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(KEYINPUT103), .B1(new_n384_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n376_), .A2(new_n379_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n380_), .A2(new_n383_), .ZN(new_n392_));
  AND4_X1   g191(.A1(KEYINPUT103), .A2(new_n391_), .A3(new_n389_), .A4(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n390_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n361_), .A2(new_n366_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n374_), .A2(new_n290_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n381_), .B1(new_n397_), .B2(new_n233_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n379_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n398_), .A2(KEYINPUT102), .A3(new_n399_), .A4(new_n355_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT102), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n401_), .B1(new_n376_), .B2(new_n379_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n396_), .A2(new_n232_), .A3(new_n364_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n383_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n379_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n400_), .A2(new_n402_), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n389_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n354_), .B1(new_n394_), .B2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n391_), .A2(new_n392_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(new_n407_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n384_), .A2(new_n389_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(new_n354_), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n329_), .B(new_n353_), .C1(new_n409_), .C2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n326_), .ZN(new_n416_));
  OR2_X1    g215(.A1(KEYINPUT100), .A2(KEYINPUT33), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n351_), .B(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n332_), .A2(new_n333_), .A3(new_n336_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT101), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n420_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n330_), .A2(new_n334_), .A3(new_n331_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n421_), .A2(new_n349_), .A3(new_n422_), .A4(new_n423_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n418_), .A2(new_n412_), .A3(new_n411_), .A4(new_n424_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n389_), .A2(KEYINPUT32), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n406_), .A2(new_n426_), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n410_), .A2(new_n426_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n427_), .A2(new_n428_), .A3(new_n352_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n416_), .B1(new_n425_), .B2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n257_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n415_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT13), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G230gat), .A2(G233gat), .ZN(new_n435_));
  INV_X1    g234(.A(G99gat), .ZN(new_n436_));
  INV_X1    g235(.A(G106gat), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(new_n437_), .A3(KEYINPUT7), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT7), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n439_), .B1(G99gat), .B2(G106gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n438_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G99gat), .A2(G106gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT6), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT6), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n444_), .A2(G99gat), .A3(G106gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n441_), .A2(new_n446_), .A3(KEYINPUT65), .ZN(new_n447_));
  INV_X1    g246(.A(G85gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n388_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G85gat), .A2(G92gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n451_), .A2(KEYINPUT66), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n447_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT8), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n436_), .A2(KEYINPUT10), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n436_), .A2(KEYINPUT10), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n437_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT9), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT64), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT64), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT9), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n449_), .A2(new_n460_), .A3(new_n462_), .A4(new_n450_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n459_), .A2(G85gat), .A3(G92gat), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n458_), .A2(new_n463_), .A3(new_n446_), .A4(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n441_), .A2(new_n446_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n451_), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT65), .B1(new_n454_), .B2(KEYINPUT66), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n455_), .A2(new_n465_), .A3(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G71gat), .B(G78gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G57gat), .B(G64gat), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(KEYINPUT11), .A3(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(KEYINPUT11), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(new_n471_), .ZN(new_n476_));
  OR2_X1    g275(.A1(new_n473_), .A2(KEYINPUT11), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n474_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT68), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT68), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n474_), .A2(new_n476_), .A3(new_n480_), .A4(new_n477_), .ZN(new_n481_));
  AND4_X1   g280(.A1(KEYINPUT12), .A2(new_n470_), .A3(new_n479_), .A4(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT67), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n455_), .A2(new_n483_), .A3(new_n465_), .A4(new_n469_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n469_), .A2(new_n465_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT8), .B1(new_n447_), .B2(new_n452_), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT67), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n478_), .B1(new_n484_), .B2(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n482_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n484_), .A2(new_n487_), .A3(new_n478_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT12), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n490_), .A2(KEYINPUT69), .A3(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT69), .B1(new_n490_), .B2(new_n491_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n435_), .B(new_n489_), .C1(new_n492_), .C2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT70), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n490_), .A2(new_n491_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT69), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n490_), .A2(KEYINPUT69), .A3(new_n491_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT70), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n500_), .A2(new_n501_), .A3(new_n435_), .A4(new_n489_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n495_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n478_), .ZN(new_n504_));
  AND2_X1   g303(.A1(new_n469_), .A2(new_n465_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n483_), .B1(new_n505_), .B2(new_n455_), .ZN(new_n506_));
  NOR3_X1   g305(.A1(new_n485_), .A2(new_n486_), .A3(KEYINPUT67), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n504_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(new_n490_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n435_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G120gat), .B(G148gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT5), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G176gat), .B(G204gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n515_), .B(new_n516_), .Z(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n503_), .A2(new_n511_), .A3(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n518_), .B1(new_n503_), .B2(new_n511_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n434_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n503_), .A2(new_n511_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(new_n517_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n503_), .A2(new_n511_), .A3(new_n518_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(new_n524_), .A3(KEYINPUT13), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n521_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT81), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G229gat), .A2(G233gat), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT14), .ZN(new_n530_));
  XNOR2_X1  g329(.A(KEYINPUT79), .B(G8gat), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n530_), .B1(new_n531_), .B2(G1gat), .ZN(new_n532_));
  XOR2_X1   g331(.A(G15gat), .B(G22gat), .Z(new_n533_));
  NOR3_X1   g332(.A1(new_n532_), .A2(G1gat), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(G1gat), .ZN(new_n535_));
  INV_X1    g334(.A(G8gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT79), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT79), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(G8gat), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n537_), .A2(new_n539_), .A3(G1gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT14), .ZN(new_n541_));
  INV_X1    g340(.A(new_n533_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n535_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  NOR3_X1   g342(.A1(new_n534_), .A2(new_n543_), .A3(new_n536_), .ZN(new_n544_));
  OAI21_X1  g343(.A(G1gat), .B1(new_n532_), .B2(new_n533_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n541_), .A2(new_n542_), .A3(new_n535_), .ZN(new_n546_));
  AOI21_X1  g345(.A(G8gat), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n544_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT15), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G29gat), .A2(G36gat), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(G29gat), .A2(G36gat), .ZN(new_n552_));
  OAI21_X1  g351(.A(G43gat), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(G29gat), .ZN(new_n554_));
  INV_X1    g353(.A(G36gat), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(G43gat), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n556_), .A2(new_n557_), .A3(new_n550_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n553_), .A2(G50gat), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(G50gat), .B1(new_n553_), .B2(new_n558_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n549_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n561_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n563_), .A2(KEYINPUT15), .A3(new_n559_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n548_), .A2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n536_), .B1(new_n534_), .B2(new_n543_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n545_), .A2(G8gat), .A3(new_n546_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n563_), .A2(new_n559_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(KEYINPUT80), .B1(new_n569_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT80), .ZN(new_n573_));
  AOI211_X1 g372(.A(new_n573_), .B(new_n570_), .C1(new_n567_), .C2(new_n568_), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n529_), .B(new_n566_), .C1(new_n572_), .C2(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n569_), .A2(new_n571_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n573_), .B1(new_n548_), .B2(new_n570_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n569_), .A2(KEYINPUT80), .A3(new_n571_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n576_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n528_), .B(new_n575_), .C1(new_n579_), .C2(new_n529_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT83), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G113gat), .B(G141gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT82), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(new_n268_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(new_n226_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n582_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n586_), .ZN(new_n588_));
  AOI21_X1  g387(.A(KEYINPUT81), .B1(new_n588_), .B2(new_n581_), .ZN(new_n589_));
  OAI22_X1  g388(.A1(new_n572_), .A2(new_n574_), .B1(new_n569_), .B2(new_n571_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n529_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n589_), .B1(new_n592_), .B2(new_n575_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(KEYINPUT84), .B1(new_n587_), .B2(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n588_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT84), .ZN(new_n597_));
  NOR3_X1   g396(.A1(new_n596_), .A2(new_n597_), .A3(new_n593_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n595_), .A2(new_n598_), .ZN(new_n599_));
  NOR3_X1   g398(.A1(new_n433_), .A2(new_n527_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT104), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n569_), .B(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(new_n504_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G127gat), .B(G155gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT16), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(G183gat), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n607_), .B(G211gat), .Z(new_n608_));
  INV_X1    g407(.A(KEYINPUT17), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n608_), .A2(new_n609_), .ZN(new_n611_));
  OR3_X1    g410(.A1(new_n604_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n479_), .A2(new_n481_), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n603_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n603_), .A2(new_n613_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n614_), .A2(new_n610_), .A3(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n612_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G232gat), .A2(G233gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT73), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT34), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT74), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n565_), .A2(new_n621_), .A3(new_n470_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n621_), .B1(new_n565_), .B2(new_n470_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n570_), .B1(new_n484_), .B2(new_n487_), .ZN(new_n625_));
  OAI211_X1 g424(.A(KEYINPUT35), .B(new_n620_), .C1(new_n624_), .C2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n565_), .A2(new_n470_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT74), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n565_), .A2(new_n470_), .A3(new_n621_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n620_), .A2(KEYINPUT35), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n620_), .A2(KEYINPUT35), .ZN(new_n632_));
  INV_X1    g431(.A(new_n625_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n630_), .A2(new_n631_), .A3(new_n632_), .A4(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n626_), .A2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(G190gat), .B(G218gat), .ZN(new_n636_));
  INV_X1    g435(.A(G134gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(G162gat), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT36), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT76), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  OR2_X1    g442(.A1(new_n641_), .A2(new_n642_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n635_), .A2(new_n643_), .A3(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT77), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n635_), .A2(KEYINPUT77), .A3(new_n643_), .A4(new_n644_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n639_), .A2(new_n640_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n626_), .A2(new_n649_), .A3(new_n634_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(KEYINPUT75), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT75), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n626_), .A2(new_n652_), .A3(new_n634_), .A4(new_n649_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n647_), .A2(new_n648_), .A3(new_n651_), .A4(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT37), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT37), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n645_), .A2(new_n656_), .A3(new_n650_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT78), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT78), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n645_), .A2(new_n659_), .A3(new_n656_), .A4(new_n650_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n617_), .B1(new_n655_), .B2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n600_), .A2(new_n601_), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n599_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n526_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n415_), .A2(new_n432_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n655_), .A2(new_n661_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n617_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(KEYINPUT104), .B1(new_n667_), .B2(new_n670_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n663_), .A2(new_n671_), .A3(new_n535_), .A4(new_n352_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT38), .ZN(new_n673_));
  OR3_X1    g472(.A1(new_n672_), .A2(KEYINPUT105), .A3(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n645_), .A2(new_n650_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n667_), .A2(new_n676_), .A3(new_n617_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n535_), .B1(new_n677_), .B2(new_n352_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n672_), .B1(new_n678_), .B2(new_n673_), .ZN(new_n679_));
  OAI21_X1  g478(.A(KEYINPUT105), .B1(new_n672_), .B2(new_n673_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n674_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n681_), .B(new_n682_), .ZN(G1324gat));
  NAND2_X1  g482(.A1(new_n663_), .A2(new_n671_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n390_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n393_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n685_), .A2(new_n686_), .A3(new_n408_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT27), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(new_n413_), .ZN(new_n689_));
  OR3_X1    g488(.A1(new_n684_), .A2(new_n531_), .A3(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n689_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n617_), .A2(new_n676_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n600_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(G8gat), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT107), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT39), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n693_), .A2(new_n697_), .A3(G8gat), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n695_), .A2(new_n696_), .A3(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n696_), .B1(new_n695_), .B2(new_n698_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n690_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT40), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  OAI211_X1 g502(.A(new_n690_), .B(KEYINPUT40), .C1(new_n699_), .C2(new_n700_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1325gat));
  NAND2_X1  g504(.A1(new_n677_), .A2(new_n416_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(G15gat), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT41), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT41), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n706_), .A2(new_n709_), .A3(G15gat), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n326_), .A2(G15gat), .ZN(new_n711_));
  OAI211_X1 g510(.A(new_n708_), .B(new_n710_), .C1(new_n684_), .C2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n712_), .B(new_n713_), .ZN(G1326gat));
  NAND2_X1  g513(.A1(new_n677_), .A2(new_n257_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(G22gat), .ZN(new_n716_));
  XNOR2_X1  g515(.A(KEYINPUT109), .B(KEYINPUT42), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n716_), .B(new_n717_), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n684_), .A2(G22gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n431_), .B2(new_n719_), .ZN(G1327gat));
  NOR3_X1   g519(.A1(new_n667_), .A2(new_n675_), .A3(new_n669_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n721_), .A2(new_n554_), .A3(new_n352_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT43), .ZN(new_n723_));
  INV_X1    g522(.A(new_n668_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n666_), .A2(new_n723_), .A3(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n723_), .B1(new_n666_), .B2(new_n724_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n665_), .B(new_n617_), .C1(new_n725_), .C2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n666_), .A2(new_n724_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT43), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n666_), .A2(new_n723_), .A3(new_n724_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n733_), .A2(KEYINPUT44), .A3(new_n665_), .A4(new_n617_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n729_), .A2(new_n734_), .A3(new_n352_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT110), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n735_), .A2(new_n736_), .A3(G29gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n735_), .B2(G29gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n722_), .B1(new_n737_), .B2(new_n738_), .ZN(G1328gat));
  NAND3_X1  g538(.A1(new_n729_), .A2(new_n734_), .A3(new_n691_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(G36gat), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT113), .ZN(new_n742_));
  XNOR2_X1  g541(.A(KEYINPUT111), .B(KEYINPUT112), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT45), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n721_), .A2(new_n555_), .A3(new_n691_), .A4(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n744_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n669_), .A2(new_n675_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n600_), .A2(new_n555_), .A3(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n746_), .B1(new_n748_), .B2(new_n689_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n745_), .A2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n741_), .A2(new_n742_), .A3(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n689_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n555_), .B1(new_n752_), .B2(new_n734_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n745_), .A2(new_n749_), .ZN(new_n754_));
  OAI21_X1  g553(.A(KEYINPUT113), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n751_), .A2(new_n755_), .A3(KEYINPUT46), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT46), .B1(new_n751_), .B2(new_n755_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n756_), .A2(new_n757_), .ZN(G1329gat));
  INV_X1    g557(.A(new_n721_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n557_), .B1(new_n759_), .B2(new_n326_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n734_), .A2(G43gat), .A3(new_n416_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n729_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n760_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g563(.A(G50gat), .B1(new_n721_), .B2(new_n257_), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n729_), .A2(G50gat), .A3(new_n257_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(new_n734_), .ZN(G1331gat));
  NOR3_X1   g566(.A1(new_n433_), .A2(new_n664_), .A3(new_n526_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n692_), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n769_), .A2(new_n347_), .A3(new_n353_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n662_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(new_n352_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n770_), .B1(new_n347_), .B2(new_n773_), .ZN(G1332gat));
  OR3_X1    g573(.A1(new_n771_), .A2(G64gat), .A3(new_n689_), .ZN(new_n775_));
  OAI21_X1  g574(.A(G64gat), .B1(new_n769_), .B2(new_n689_), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n776_), .A2(KEYINPUT114), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(KEYINPUT114), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n777_), .A2(KEYINPUT48), .A3(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(KEYINPUT48), .B1(new_n777_), .B2(new_n778_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n775_), .B1(new_n779_), .B2(new_n780_), .ZN(G1333gat));
  OAI21_X1  g580(.A(G71gat), .B1(new_n769_), .B2(new_n326_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT49), .ZN(new_n783_));
  OR2_X1    g582(.A1(new_n326_), .A2(G71gat), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n783_), .B1(new_n771_), .B2(new_n784_), .ZN(G1334gat));
  OR3_X1    g584(.A1(new_n771_), .A2(G78gat), .A3(new_n431_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n768_), .A2(new_n257_), .A3(new_n692_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n787_), .A2(G78gat), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(new_n789_), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n790_), .A2(KEYINPUT50), .A3(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT50), .B1(new_n790_), .B2(new_n791_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n786_), .B1(new_n792_), .B2(new_n793_), .ZN(G1335gat));
  AND2_X1   g593(.A1(new_n768_), .A2(new_n747_), .ZN(new_n795_));
  AOI21_X1  g594(.A(G85gat), .B1(new_n795_), .B2(new_n352_), .ZN(new_n796_));
  OR3_X1    g595(.A1(new_n725_), .A2(new_n726_), .A3(KEYINPUT116), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n733_), .A2(KEYINPUT116), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n526_), .A2(new_n664_), .A3(new_n669_), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n797_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n353_), .A2(new_n448_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n796_), .B1(new_n800_), .B2(new_n801_), .ZN(G1336gat));
  AOI21_X1  g601(.A(G92gat), .B1(new_n795_), .B2(new_n691_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n689_), .A2(new_n388_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n803_), .B1(new_n800_), .B2(new_n804_), .ZN(G1337gat));
  NAND4_X1  g604(.A1(new_n797_), .A2(new_n798_), .A3(new_n416_), .A4(new_n799_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(G99gat), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n456_), .A2(new_n457_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n326_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n795_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n807_), .A2(new_n810_), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n811_), .A2(KEYINPUT117), .A3(KEYINPUT51), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT117), .B1(new_n811_), .B2(KEYINPUT51), .ZN(new_n813_));
  XNOR2_X1  g612(.A(KEYINPUT118), .B(KEYINPUT51), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n811_), .A2(KEYINPUT119), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT119), .ZN(new_n816_));
  AOI22_X1  g615(.A1(new_n806_), .A2(G99gat), .B1(new_n795_), .B2(new_n809_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n814_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n816_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  OAI22_X1  g618(.A1(new_n812_), .A2(new_n813_), .B1(new_n815_), .B2(new_n819_), .ZN(G1338gat));
  NAND3_X1  g619(.A1(new_n795_), .A2(new_n437_), .A3(new_n257_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n733_), .A2(new_n257_), .A3(new_n799_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n822_), .A2(new_n823_), .A3(G106gat), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n823_), .B1(new_n822_), .B2(G106gat), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n821_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g626(.A1(new_n599_), .A2(new_n521_), .A3(new_n525_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n670_), .A2(KEYINPUT54), .A3(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830_));
  INV_X1    g629(.A(new_n828_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n830_), .B1(new_n831_), .B2(new_n662_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n829_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n592_), .A2(new_n575_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n588_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n591_), .B(new_n566_), .C1(new_n572_), .C2(new_n574_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n836_), .B1(new_n579_), .B2(new_n591_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n586_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n835_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n613_), .A2(KEYINPUT12), .A3(new_n470_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n508_), .A2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n842_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n501_), .B1(new_n843_), .B2(new_n435_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n494_), .A2(KEYINPUT70), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n840_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n843_), .A2(KEYINPUT55), .A3(new_n435_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n489_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n510_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n847_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n846_), .A2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT56), .B1(new_n851_), .B2(new_n517_), .ZN(new_n852_));
  AOI21_X1  g651(.A(KEYINPUT55), .B1(new_n495_), .B2(new_n502_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n847_), .A2(new_n849_), .ZN(new_n854_));
  OAI211_X1 g653(.A(KEYINPUT56), .B(new_n517_), .C1(new_n853_), .C2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n524_), .B(new_n839_), .C1(new_n852_), .C2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT58), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n517_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT56), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n855_), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n863_), .A2(KEYINPUT58), .A3(new_n524_), .A4(new_n839_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n859_), .A2(new_n724_), .A3(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n866_));
  AOI22_X1  g665(.A1(new_n523_), .A2(new_n524_), .B1(new_n838_), .B2(new_n835_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n598_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n597_), .B1(new_n596_), .B2(new_n593_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n519_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n867_), .B1(new_n870_), .B2(new_n863_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n866_), .B1(new_n871_), .B2(new_n676_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n524_), .B1(new_n595_), .B2(new_n598_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n873_), .B1(new_n862_), .B2(new_n855_), .ZN(new_n874_));
  OAI211_X1 g673(.A(KEYINPUT57), .B(new_n675_), .C1(new_n874_), .C2(new_n867_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n865_), .A2(new_n872_), .A3(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n833_), .B1(new_n876_), .B2(new_n617_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n691_), .A2(new_n353_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n877_), .A2(new_n328_), .A3(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(G113gat), .B1(new_n880_), .B2(new_n664_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT59), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n876_), .A2(new_n617_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n833_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n328_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n882_), .B1(new_n885_), .B2(new_n878_), .ZN(new_n886_));
  NOR4_X1   g685(.A1(new_n877_), .A2(KEYINPUT59), .A3(new_n328_), .A4(new_n879_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n664_), .A2(G113gat), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n881_), .B1(new_n888_), .B2(new_n889_), .ZN(G1340gat));
  XOR2_X1   g689(.A(KEYINPUT120), .B(G120gat), .Z(new_n891_));
  OAI21_X1  g690(.A(new_n891_), .B1(new_n526_), .B2(KEYINPUT60), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n880_), .B(new_n892_), .C1(KEYINPUT60), .C2(new_n891_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n886_), .A2(new_n887_), .A3(new_n526_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n894_), .B2(new_n891_), .ZN(G1341gat));
  INV_X1    g694(.A(KEYINPUT122), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n669_), .A2(G127gat), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(KEYINPUT121), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n886_), .A2(new_n887_), .A3(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(G127gat), .B1(new_n880_), .B2(new_n669_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n896_), .B1(new_n900_), .B2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n885_), .A2(new_n878_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(KEYINPUT59), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n880_), .A2(new_n882_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n904_), .A2(new_n905_), .A3(new_n898_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n901_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n906_), .A2(KEYINPUT122), .A3(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n902_), .A2(new_n908_), .ZN(G1342gat));
  OAI21_X1  g708(.A(new_n637_), .B1(new_n903_), .B2(new_n675_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(KEYINPUT123), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n904_), .A2(G134gat), .A3(new_n905_), .A4(new_n724_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT123), .ZN(new_n913_));
  OAI211_X1 g712(.A(new_n913_), .B(new_n637_), .C1(new_n903_), .C2(new_n675_), .ZN(new_n914_));
  AND3_X1   g713(.A1(new_n911_), .A2(new_n912_), .A3(new_n914_), .ZN(G1343gat));
  NOR3_X1   g714(.A1(new_n877_), .A2(new_n327_), .A3(new_n879_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n664_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g717(.A1(new_n916_), .A2(new_n527_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g719(.A1(new_n916_), .A2(new_n669_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(KEYINPUT61), .B(G155gat), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n921_), .B(new_n922_), .ZN(G1346gat));
  AOI21_X1  g722(.A(G162gat), .B1(new_n916_), .B2(new_n676_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n724_), .A2(G162gat), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(KEYINPUT124), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n924_), .B1(new_n916_), .B2(new_n926_), .ZN(G1347gat));
  NOR2_X1   g726(.A1(new_n877_), .A2(new_n257_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n689_), .A2(new_n352_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n930_), .A2(new_n599_), .A3(new_n326_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n928_), .A2(new_n288_), .A3(new_n931_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n931_), .B(KEYINPUT125), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n268_), .B1(new_n928_), .B2(new_n933_), .ZN(new_n934_));
  XOR2_X1   g733(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n935_));
  AND2_X1   g734(.A1(new_n934_), .A2(new_n935_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n934_), .A2(new_n935_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n932_), .B1(new_n936_), .B2(new_n937_), .ZN(G1348gat));
  NOR3_X1   g737(.A1(new_n877_), .A2(new_n328_), .A3(new_n930_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(new_n527_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g740(.A1(new_n939_), .A2(new_n669_), .ZN(new_n942_));
  MUX2_X1   g741(.A(new_n358_), .B(G183gat), .S(new_n942_), .Z(G1350gat));
  NAND2_X1  g742(.A1(new_n676_), .A2(new_n359_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(KEYINPUT127), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n939_), .A2(new_n945_), .ZN(new_n946_));
  AND2_X1   g745(.A1(new_n939_), .A2(new_n724_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n946_), .B1(new_n947_), .B2(new_n277_), .ZN(G1351gat));
  NOR3_X1   g747(.A1(new_n877_), .A2(new_n327_), .A3(new_n930_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n949_), .A2(new_n664_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g750(.A1(new_n949_), .A2(new_n527_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n952_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g752(.A1(new_n949_), .A2(new_n669_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n955_));
  AND2_X1   g754(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n956_));
  NOR3_X1   g755(.A1(new_n954_), .A2(new_n955_), .A3(new_n956_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n957_), .B1(new_n954_), .B2(new_n955_), .ZN(G1354gat));
  AOI21_X1  g757(.A(G218gat), .B1(new_n949_), .B2(new_n676_), .ZN(new_n959_));
  AND2_X1   g758(.A1(new_n724_), .A2(G218gat), .ZN(new_n960_));
  AOI21_X1  g759(.A(new_n959_), .B1(new_n949_), .B2(new_n960_), .ZN(G1355gat));
endmodule


