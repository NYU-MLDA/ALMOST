//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 1 1 0 1 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n793_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n800_, new_n802_, new_n803_, new_n805_, new_n806_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n821_, new_n822_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n830_, new_n831_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  AND2_X1   g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT84), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G155gat), .ZN(new_n207_));
  INV_X1    g006(.A(G162gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT84), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n209_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n206_), .A2(new_n212_), .ZN(new_n213_));
  AOI21_X1  g012(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n214_), .A2(KEYINPUT83), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(KEYINPUT83), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n213_), .B1(new_n217_), .B2(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n205_), .B1(KEYINPUT1), .B2(new_n211_), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n211_), .A2(KEYINPUT1), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  XOR2_X1   g026(.A(G141gat), .B(G148gat), .Z(new_n228_));
  AND2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n224_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT29), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT90), .ZN(new_n233_));
  INV_X1    g032(.A(G211gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n234_), .A2(G218gat), .ZN(new_n235_));
  INV_X1    g034(.A(G218gat), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n236_), .A2(G211gat), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n233_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n236_), .A2(G211gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n234_), .A2(G218gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n240_), .A3(KEYINPUT90), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(G204gat), .ZN(new_n243_));
  OAI21_X1  g042(.A(KEYINPUT88), .B1(new_n243_), .B2(G197gat), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT88), .ZN(new_n245_));
  INV_X1    g044(.A(G197gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(new_n246_), .A3(G204gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n243_), .A2(G197gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n244_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT21), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n242_), .A2(new_n250_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n244_), .A2(new_n248_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT89), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT21), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n252_), .A2(new_n253_), .A3(new_n254_), .A4(new_n247_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n244_), .A2(new_n247_), .A3(new_n254_), .A4(new_n248_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT89), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT87), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G197gat), .B(G204gat), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n259_), .B1(new_n260_), .B2(new_n254_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n246_), .A2(G204gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(new_n248_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n263_), .A2(KEYINPUT87), .A3(KEYINPUT21), .ZN(new_n264_));
  AOI22_X1  g063(.A1(new_n261_), .A2(new_n264_), .B1(new_n238_), .B2(new_n241_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n251_), .B1(new_n258_), .B2(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n203_), .B1(new_n232_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT91), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT91), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n269_), .B(new_n203_), .C1(new_n232_), .C2(new_n266_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n251_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n256_), .B(new_n253_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n261_), .A2(new_n264_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(new_n242_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n272_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT85), .B1(new_n224_), .B2(new_n229_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n227_), .A2(new_n228_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT85), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n280_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n278_), .B(new_n279_), .C1(new_n281_), .C2(new_n213_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n277_), .A2(new_n282_), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n202_), .B(new_n276_), .C1(new_n283_), .C2(new_n231_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G78gat), .B(G106gat), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n271_), .A2(new_n284_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n286_), .B1(new_n271_), .B2(new_n284_), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT92), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n271_), .A2(new_n284_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(new_n285_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT92), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n292_), .A2(new_n293_), .A3(new_n287_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n283_), .A2(new_n231_), .ZN(new_n295_));
  XOR2_X1   g094(.A(G22gat), .B(G50gat), .Z(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n295_), .A2(new_n297_), .ZN(new_n300_));
  XOR2_X1   g099(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n301_));
  OR3_X1    g100(.A1(new_n299_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n301_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n290_), .A2(new_n294_), .A3(new_n305_), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n304_), .A2(new_n293_), .A3(new_n287_), .A4(new_n292_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G169gat), .A2(G176gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT77), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT77), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n312_), .A2(G169gat), .A3(G176gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(G183gat), .ZN(new_n315_));
  INV_X1    g114(.A(G190gat), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT23), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT23), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(G183gat), .A3(G190gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n315_), .A2(new_n316_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n314_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT80), .ZN(new_n323_));
  INV_X1    g122(.A(G169gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT22), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT22), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(G169gat), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n323_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n323_), .B1(new_n326_), .B2(G169gat), .ZN(new_n329_));
  INV_X1    g128(.A(G176gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NOR3_X1   g130(.A1(new_n328_), .A2(new_n331_), .A3(KEYINPUT81), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT81), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n326_), .A2(G169gat), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n324_), .A2(KEYINPUT22), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT80), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(G176gat), .B1(new_n325_), .B2(new_n323_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n333_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n322_), .B1(new_n332_), .B2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT79), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n319_), .A2(KEYINPUT78), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT78), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n342_), .A2(new_n318_), .A3(G183gat), .A4(G190gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(new_n317_), .A3(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n324_), .A2(new_n330_), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n345_), .A2(KEYINPUT24), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n340_), .B1(new_n344_), .B2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n344_), .A2(new_n340_), .A3(new_n346_), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n311_), .A2(new_n313_), .A3(new_n345_), .A4(KEYINPUT24), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n315_), .A2(KEYINPUT25), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT25), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(G183gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n316_), .A2(KEYINPUT26), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT26), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(G190gat), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n350_), .A2(new_n352_), .A3(new_n353_), .A4(new_n355_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n349_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n348_), .A2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n339_), .B1(new_n347_), .B2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT30), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G71gat), .B(G99gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(G43gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G227gat), .A2(G233gat), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n363_), .B(G15gat), .Z(new_n364_));
  XNOR2_X1  g163(.A(new_n362_), .B(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n360_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G127gat), .B(G134gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G113gat), .B(G120gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n369_), .B(KEYINPUT31), .Z(new_n370_));
  NOR2_X1   g169(.A1(new_n370_), .A2(KEYINPUT82), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n366_), .B(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n369_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n277_), .A2(new_n374_), .A3(new_n282_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G225gat), .A2(G233gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n230_), .A2(new_n369_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G1gat), .B(G29gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT0), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(G57gat), .ZN(new_n381_));
  OR2_X1    g180(.A1(new_n379_), .A2(KEYINPUT0), .ZN(new_n382_));
  INV_X1    g181(.A(G57gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n379_), .A2(KEYINPUT0), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n381_), .A2(new_n385_), .A3(G85gat), .ZN(new_n386_));
  AOI21_X1  g185(.A(G85gat), .B1(new_n381_), .B2(new_n385_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n375_), .A2(KEYINPUT4), .A3(new_n377_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n369_), .A2(KEYINPUT4), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n277_), .A2(new_n282_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n376_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n378_), .B(new_n389_), .C1(new_n390_), .C2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n375_), .A2(KEYINPUT4), .A3(new_n377_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n397_), .A2(new_n393_), .A3(new_n392_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n389_), .B1(new_n398_), .B2(new_n378_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n396_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G226gat), .A2(G233gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT19), .ZN(new_n402_));
  XOR2_X1   g201(.A(new_n402_), .B(KEYINPUT93), .Z(new_n403_));
  NOR2_X1   g202(.A1(new_n359_), .A2(new_n276_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n346_), .A2(new_n356_), .A3(new_n320_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n310_), .A2(KEYINPUT24), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n406_), .A2(KEYINPUT94), .B1(new_n324_), .B2(new_n330_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n407_), .B1(KEYINPUT94), .B2(new_n406_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n344_), .A2(new_n321_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n334_), .A2(new_n335_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n314_), .B1(new_n410_), .B2(new_n330_), .ZN(new_n411_));
  AOI22_X1  g210(.A1(new_n405_), .A2(new_n408_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT20), .B1(new_n266_), .B2(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n403_), .B1(new_n404_), .B2(new_n413_), .ZN(new_n414_));
  XOR2_X1   g213(.A(G8gat), .B(G36gat), .Z(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT18), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G64gat), .B(G92gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n359_), .A2(new_n276_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT20), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n420_), .B1(new_n266_), .B2(new_n412_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n402_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n419_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n414_), .A2(new_n418_), .A3(new_n423_), .ZN(new_n424_));
  NOR3_X1   g223(.A1(new_n404_), .A2(new_n413_), .A3(new_n403_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n422_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  OAI211_X1 g226(.A(KEYINPUT27), .B(new_n424_), .C1(new_n427_), .C2(new_n418_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT95), .ZN(new_n429_));
  AOI211_X1 g228(.A(new_n429_), .B(new_n418_), .C1(new_n414_), .C2(new_n423_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n418_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n414_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n423_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n431_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n424_), .A2(KEYINPUT95), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n430_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  OAI211_X1 g235(.A(new_n400_), .B(new_n428_), .C1(new_n436_), .C2(KEYINPUT27), .ZN(new_n437_));
  NOR3_X1   g236(.A1(new_n309_), .A2(new_n373_), .A3(new_n437_), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n397_), .A2(new_n376_), .A3(new_n392_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n375_), .A2(new_n393_), .A3(new_n377_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(new_n388_), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT96), .B1(new_n439_), .B2(new_n441_), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n440_), .A2(new_n388_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT96), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n397_), .A2(new_n376_), .A3(new_n392_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n443_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT33), .ZN(new_n447_));
  AOI22_X1  g246(.A1(new_n442_), .A2(new_n446_), .B1(new_n447_), .B2(new_n395_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n398_), .A2(KEYINPUT33), .A3(new_n378_), .A4(new_n389_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n436_), .A2(new_n448_), .A3(KEYINPUT97), .A4(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n418_), .A2(KEYINPUT32), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n414_), .A2(new_n423_), .A3(new_n451_), .ZN(new_n452_));
  OAI221_X1 g251(.A(new_n452_), .B1(new_n427_), .B2(new_n451_), .C1(new_n396_), .C2(new_n399_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n450_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n395_), .A2(new_n447_), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n443_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n444_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n449_), .B(new_n455_), .C1(new_n456_), .C2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(KEYINPUT97), .B1(new_n459_), .B2(new_n436_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n308_), .B1(new_n454_), .B2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT98), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT98), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n308_), .B(new_n463_), .C1(new_n454_), .C2(new_n460_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n308_), .A2(new_n437_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n462_), .A2(new_n464_), .A3(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n438_), .B1(new_n467_), .B2(new_n373_), .ZN(new_n468_));
  XOR2_X1   g267(.A(G71gat), .B(G78gat), .Z(new_n469_));
  XNOR2_X1  g268(.A(G57gat), .B(G64gat), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n469_), .B1(KEYINPUT11), .B2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT67), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(KEYINPUT11), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT8), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G99gat), .A2(G106gat), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT6), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT66), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n476_), .B(KEYINPUT6), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT66), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(G99gat), .A2(G106gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT7), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n479_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G85gat), .B(G92gat), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n475_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(KEYINPUT65), .B(KEYINPUT8), .Z(new_n489_));
  AOI211_X1 g288(.A(new_n486_), .B(new_n489_), .C1(new_n484_), .C2(new_n480_), .ZN(new_n490_));
  INV_X1    g289(.A(G106gat), .ZN(new_n491_));
  XOR2_X1   g290(.A(KEYINPUT10), .B(G99gat), .Z(new_n492_));
  AOI21_X1  g291(.A(new_n478_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n494_), .B1(new_n486_), .B2(KEYINPUT9), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT64), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n495_), .A2(KEYINPUT64), .ZN(new_n498_));
  OAI22_X1  g297(.A1(new_n488_), .A2(new_n490_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n474_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT12), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n474_), .A2(new_n499_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n474_), .A2(KEYINPUT12), .A3(new_n499_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  AND2_X1   g304(.A1(G230gat), .A2(G233gat), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n503_), .A2(new_n500_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(new_n506_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G120gat), .B(G148gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT5), .ZN(new_n512_));
  XOR2_X1   g311(.A(G176gat), .B(G204gat), .Z(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n510_), .A2(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n510_), .A2(new_n514_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT13), .ZN(new_n518_));
  OR2_X1    g317(.A1(new_n518_), .A2(KEYINPUT68), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(KEYINPUT68), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n517_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  OAI211_X1 g320(.A(KEYINPUT68), .B(new_n518_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G113gat), .B(G141gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G169gat), .B(G197gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G15gat), .B(G22gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT71), .B(G8gat), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n530_), .A2(G1gat), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT14), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n529_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G1gat), .B(G8gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(G29gat), .B(G36gat), .Z(new_n536_));
  XNOR2_X1  g335(.A(G43gat), .B(G50gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n535_), .A2(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n538_), .B(KEYINPUT15), .Z(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n535_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G229gat), .A2(G233gat), .ZN(new_n543_));
  XOR2_X1   g342(.A(new_n543_), .B(KEYINPUT75), .Z(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n535_), .B(new_n538_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT73), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n543_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n545_), .B1(new_n550_), .B2(KEYINPUT74), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(KEYINPUT74), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n528_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n553_), .ZN(new_n555_));
  NOR3_X1   g354(.A1(new_n555_), .A2(new_n551_), .A3(new_n527_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT76), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n552_), .A2(new_n553_), .A3(new_n528_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n527_), .B1(new_n555_), .B2(new_n551_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT76), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n559_), .A2(new_n563_), .ZN(new_n564_));
  NOR3_X1   g363(.A1(new_n468_), .A2(new_n524_), .A3(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(G190gat), .B(G218gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(G134gat), .B(G162gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G232gat), .A2(G233gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT34), .ZN(new_n570_));
  OAI22_X1  g369(.A1(new_n499_), .A2(new_n538_), .B1(KEYINPUT35), .B2(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n571_), .B1(new_n499_), .B2(new_n540_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(KEYINPUT35), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n568_), .B1(new_n574_), .B2(KEYINPUT69), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT36), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n575_), .B(new_n576_), .C1(new_n568_), .C2(new_n574_), .ZN(new_n577_));
  OAI211_X1 g376(.A(KEYINPUT36), .B(new_n568_), .C1(new_n574_), .C2(KEYINPUT69), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(KEYINPUT70), .B(KEYINPUT37), .Z(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n580_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n577_), .A2(new_n578_), .A3(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n474_), .B(new_n585_), .Z(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(new_n535_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G127gat), .B(G155gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT16), .ZN(new_n589_));
  XOR2_X1   g388(.A(G183gat), .B(G211gat), .Z(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n587_), .B1(KEYINPUT17), .B2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n592_), .A2(KEYINPUT72), .A3(KEYINPUT17), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n584_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n565_), .A2(new_n597_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n598_), .A2(G1gat), .A3(new_n400_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT38), .Z(new_n600_));
  AND3_X1   g399(.A1(new_n577_), .A2(KEYINPUT99), .A3(new_n578_), .ZN(new_n601_));
  AOI21_X1  g400(.A(KEYINPUT99), .B1(new_n577_), .B2(new_n578_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n468_), .A2(new_n604_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n605_), .A2(new_n562_), .A3(new_n523_), .A4(new_n595_), .ZN(new_n606_));
  OAI21_X1  g405(.A(G1gat), .B1(new_n606_), .B2(new_n400_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n600_), .A2(new_n607_), .ZN(G1324gat));
  OAI21_X1  g407(.A(new_n428_), .B1(new_n436_), .B2(KEYINPUT27), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(G8gat), .B1(new_n606_), .B2(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(new_n611_), .B(KEYINPUT39), .Z(new_n612_));
  NOR3_X1   g411(.A1(new_n598_), .A2(new_n610_), .A3(new_n530_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT40), .ZN(G1325gat));
  NOR3_X1   g414(.A1(new_n598_), .A2(G15gat), .A3(new_n373_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT100), .Z(new_n617_));
  OAI21_X1  g416(.A(G15gat), .B1(new_n606_), .B2(new_n373_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT41), .Z(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(G1326gat));
  NOR2_X1   g419(.A1(new_n308_), .A2(G22gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT103), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n598_), .A2(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(G22gat), .B1(new_n606_), .B2(new_n308_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT102), .ZN(new_n625_));
  XOR2_X1   g424(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n626_));
  AOI21_X1  g425(.A(new_n623_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n627_), .B1(new_n625_), .B2(new_n626_), .ZN(G1327gat));
  NOR3_X1   g427(.A1(new_n524_), .A2(new_n557_), .A3(new_n595_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n584_), .ZN(new_n630_));
  OAI211_X1 g429(.A(KEYINPUT104), .B(KEYINPUT43), .C1(new_n468_), .C2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT43), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n465_), .B1(new_n461_), .B2(KEYINPUT98), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n372_), .B1(new_n633_), .B2(new_n464_), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n584_), .B(new_n632_), .C1(new_n634_), .C2(new_n438_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n631_), .A2(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n584_), .B1(new_n634_), .B2(new_n438_), .ZN(new_n637_));
  AOI21_X1  g436(.A(KEYINPUT104), .B1(new_n637_), .B2(KEYINPUT43), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n629_), .B1(new_n636_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT44), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n400_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n641_), .A2(G29gat), .A3(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n639_), .A2(new_n640_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n603_), .A2(new_n595_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n565_), .A2(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n647_), .A2(new_n400_), .ZN(new_n648_));
  OAI22_X1  g447(.A1(new_n643_), .A2(new_n645_), .B1(G29gat), .B2(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT105), .ZN(G1328gat));
  NAND3_X1  g449(.A1(new_n641_), .A2(new_n609_), .A3(new_n644_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(G36gat), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n647_), .A2(G36gat), .A3(new_n610_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n652_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT46), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n656_), .B(new_n657_), .ZN(G1329gat));
  NAND4_X1  g457(.A1(new_n641_), .A2(G43gat), .A3(new_n372_), .A4(new_n644_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n647_), .A2(new_n373_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n659_), .B1(G43gat), .B2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g461(.A1(new_n647_), .A2(G50gat), .A3(new_n308_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n641_), .A2(KEYINPUT107), .A3(new_n309_), .A4(new_n644_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n664_), .A2(G50gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n641_), .A2(new_n309_), .A3(new_n644_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT107), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(KEYINPUT108), .B1(new_n665_), .B2(new_n668_), .ZN(new_n669_));
  AND4_X1   g468(.A1(KEYINPUT108), .A2(new_n668_), .A3(G50gat), .A4(new_n664_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n663_), .B1(new_n669_), .B2(new_n670_), .ZN(G1331gat));
  AOI21_X1  g470(.A(new_n596_), .B1(new_n559_), .B2(new_n563_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n605_), .A2(new_n524_), .A3(new_n672_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n673_), .A2(new_n383_), .A3(new_n400_), .ZN(new_n674_));
  NOR3_X1   g473(.A1(new_n468_), .A2(new_n562_), .A3(new_n523_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(new_n597_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n400_), .B1(new_n676_), .B2(KEYINPUT109), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n677_), .B1(KEYINPUT109), .B2(new_n676_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n674_), .B1(new_n678_), .B2(new_n383_), .ZN(G1332gat));
  OAI21_X1  g478(.A(G64gat), .B1(new_n673_), .B2(new_n610_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT48), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n610_), .A2(G64gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n681_), .B1(new_n676_), .B2(new_n682_), .ZN(G1333gat));
  OAI21_X1  g482(.A(G71gat), .B1(new_n673_), .B2(new_n373_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT49), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n373_), .A2(G71gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n685_), .B1(new_n676_), .B2(new_n686_), .ZN(G1334gat));
  OAI21_X1  g486(.A(G78gat), .B1(new_n673_), .B2(new_n308_), .ZN(new_n688_));
  XOR2_X1   g487(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n689_));
  XNOR2_X1  g488(.A(new_n688_), .B(new_n689_), .ZN(new_n690_));
  OR2_X1    g489(.A1(new_n308_), .A2(G78gat), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n690_), .B1(new_n676_), .B2(new_n691_), .ZN(G1335gat));
  NAND2_X1  g491(.A1(new_n675_), .A2(new_n646_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n693_), .A2(G85gat), .A3(new_n400_), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n523_), .A2(new_n562_), .A3(new_n595_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT111), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n695_), .B(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n697_), .B1(new_n636_), .B2(new_n638_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT112), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n697_), .B(KEYINPUT112), .C1(new_n636_), .C2(new_n638_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(new_n642_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n694_), .B1(new_n703_), .B2(G85gat), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT113), .ZN(G1336gat));
  INV_X1    g504(.A(new_n693_), .ZN(new_n706_));
  INV_X1    g505(.A(G92gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n706_), .A2(new_n707_), .A3(new_n609_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n610_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n708_), .B1(new_n709_), .B2(new_n707_), .ZN(G1337gat));
  INV_X1    g509(.A(KEYINPUT114), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n706_), .A2(new_n372_), .A3(new_n492_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n373_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n713_));
  INV_X1    g512(.A(G99gat), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n711_), .B(new_n712_), .C1(new_n713_), .C2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT51), .ZN(new_n716_));
  OAI211_X1 g515(.A(KEYINPUT115), .B(new_n712_), .C1(new_n713_), .C2(new_n714_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT114), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n716_), .B(new_n718_), .ZN(G1338gat));
  NAND3_X1  g518(.A1(new_n706_), .A2(new_n491_), .A3(new_n309_), .ZN(new_n720_));
  OR2_X1    g519(.A1(new_n698_), .A2(new_n308_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT52), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n721_), .A2(new_n722_), .A3(G106gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n721_), .B2(G106gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n720_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  XOR2_X1   g524(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n726_));
  XNOR2_X1  g525(.A(new_n725_), .B(new_n726_), .ZN(G1339gat));
  NAND2_X1  g526(.A1(new_n610_), .A2(new_n642_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n728_), .A2(new_n373_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n630_), .A2(new_n672_), .A3(new_n523_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n730_), .A2(KEYINPUT117), .A3(KEYINPUT54), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(KEYINPUT117), .B1(new_n730_), .B2(KEYINPUT54), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n730_), .A2(KEYINPUT54), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n732_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT55), .ZN(new_n736_));
  OR2_X1    g535(.A1(new_n507_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n507_), .A2(new_n736_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n505_), .A2(new_n506_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n737_), .A2(new_n738_), .A3(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(new_n514_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT56), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n740_), .A2(KEYINPUT56), .A3(new_n514_), .ZN(new_n744_));
  AOI211_X1 g543(.A(new_n516_), .B(new_n557_), .C1(new_n743_), .C2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n548_), .A2(new_n544_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n542_), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n746_), .B(new_n527_), .C1(new_n747_), .C2(new_n544_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n560_), .A2(new_n748_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n749_), .A2(new_n517_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n603_), .B1(new_n745_), .B2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT57), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n560_), .B(new_n748_), .C1(new_n510_), .C2(new_n514_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n754_), .A2(KEYINPUT58), .ZN(new_n755_));
  AOI22_X1  g554(.A1(new_n754_), .A2(KEYINPUT58), .B1(new_n581_), .B2(new_n583_), .ZN(new_n756_));
  AOI22_X1  g555(.A1(new_n751_), .A2(new_n752_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  OAI211_X1 g556(.A(KEYINPUT57), .B(new_n603_), .C1(new_n745_), .C2(new_n750_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n595_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n308_), .B(new_n729_), .C1(new_n735_), .C2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(G113gat), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n761_), .A2(new_n762_), .A3(new_n562_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT59), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n760_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n751_), .A2(new_n752_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n755_), .A2(new_n756_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n766_), .A2(new_n758_), .A3(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n768_), .A2(new_n596_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n733_), .A2(new_n734_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n731_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n769_), .A2(new_n771_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n772_), .A2(KEYINPUT59), .A3(new_n308_), .A4(new_n729_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n564_), .B1(new_n765_), .B2(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n763_), .B1(new_n774_), .B2(new_n762_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT118), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT118), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n777_), .B(new_n763_), .C1(new_n774_), .C2(new_n762_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(G1340gat));
  INV_X1    g578(.A(KEYINPUT60), .ZN(new_n780_));
  INV_X1    g579(.A(G120gat), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n524_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n782_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n761_), .A2(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n523_), .B1(new_n765_), .B2(new_n773_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n784_), .B1(new_n785_), .B2(new_n781_), .ZN(G1341gat));
  INV_X1    g585(.A(G127gat), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n761_), .A2(new_n787_), .A3(new_n595_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n596_), .B1(new_n765_), .B2(new_n773_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n788_), .B1(new_n789_), .B2(new_n787_), .ZN(G1342gat));
  INV_X1    g589(.A(G134gat), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n761_), .A2(new_n791_), .A3(new_n604_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n630_), .B1(new_n765_), .B2(new_n773_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n792_), .B1(new_n793_), .B2(new_n791_), .ZN(G1343gat));
  NOR2_X1   g593(.A1(new_n308_), .A2(new_n372_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  AOI211_X1 g595(.A(new_n728_), .B(new_n796_), .C1(new_n769_), .C2(new_n771_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n562_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g598(.A1(new_n797_), .A2(new_n524_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g600(.A1(new_n797_), .A2(new_n595_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(KEYINPUT61), .B(G155gat), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n802_), .B(new_n803_), .ZN(G1346gat));
  NAND3_X1  g603(.A1(new_n797_), .A2(new_n208_), .A3(new_n604_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n797_), .A2(new_n584_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(new_n208_), .ZN(G1347gat));
  INV_X1    g606(.A(KEYINPUT62), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n309_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n610_), .A2(new_n642_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n811_), .A2(new_n373_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n809_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n562_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n808_), .B1(new_n815_), .B2(G169gat), .ZN(new_n816_));
  AOI211_X1 g615(.A(KEYINPUT62), .B(new_n324_), .C1(new_n814_), .C2(new_n562_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n562_), .A2(new_n410_), .ZN(new_n818_));
  XOR2_X1   g617(.A(new_n818_), .B(KEYINPUT119), .Z(new_n819_));
  OAI22_X1  g618(.A1(new_n816_), .A2(new_n817_), .B1(new_n813_), .B2(new_n819_), .ZN(G1348gat));
  NOR2_X1   g619(.A1(new_n813_), .A2(new_n523_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(KEYINPUT120), .B(G176gat), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n821_), .B(new_n822_), .ZN(G1349gat));
  NAND2_X1  g622(.A1(new_n350_), .A2(new_n352_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n814_), .A2(new_n824_), .A3(new_n595_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n825_), .A2(KEYINPUT121), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(KEYINPUT121), .ZN(new_n827_));
  AOI21_X1  g626(.A(G183gat), .B1(new_n814_), .B2(new_n595_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n826_), .A2(new_n827_), .A3(new_n828_), .ZN(G1350gat));
  OAI21_X1  g628(.A(G190gat), .B1(new_n813_), .B2(new_n630_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n604_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n813_), .B2(new_n831_), .ZN(G1351gat));
  NOR2_X1   g631(.A1(new_n796_), .A2(new_n811_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n834_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n562_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(KEYINPUT122), .B(G197gat), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n836_), .B(new_n837_), .ZN(G1352gat));
  NAND2_X1  g637(.A1(new_n835_), .A2(new_n524_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g639(.A(KEYINPUT63), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n595_), .B1(new_n841_), .B2(new_n234_), .ZN(new_n842_));
  XOR2_X1   g641(.A(new_n842_), .B(KEYINPUT123), .Z(new_n843_));
  NAND2_X1  g642(.A1(new_n835_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(KEYINPUT124), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT124), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n835_), .A2(new_n847_), .A3(new_n843_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n848_), .A2(KEYINPUT125), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(KEYINPUT125), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n846_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n851_), .ZN(new_n853_));
  AOI22_X1  g652(.A1(new_n844_), .A2(KEYINPUT124), .B1(new_n841_), .B2(new_n234_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n853_), .A2(new_n854_), .A3(new_n849_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n852_), .A2(new_n855_), .ZN(G1354gat));
  INV_X1    g655(.A(new_n835_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n857_), .A2(new_n236_), .A3(new_n630_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n857_), .A2(KEYINPUT126), .A3(new_n603_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(G218gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(KEYINPUT126), .B1(new_n857_), .B2(new_n603_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n858_), .B1(new_n860_), .B2(new_n861_), .ZN(G1355gat));
endmodule


