//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 1 1 1 0 1 0 0 1 0 0 0 0 0 1 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n773_, new_n774_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_;
  OAI21_X1  g000(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT94), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  OR3_X1    g003(.A1(KEYINPUT93), .A2(G141gat), .A3(G148gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT93), .B1(G141gat), .B2(G148gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT2), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n204_), .A2(new_n208_), .A3(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n211_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT1), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n214_), .B1(new_n213_), .B2(new_n217_), .ZN(new_n218_));
  AND3_X1   g017(.A1(new_n212_), .A2(KEYINPUT92), .A3(KEYINPUT1), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT92), .B1(new_n212_), .B2(KEYINPUT1), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n218_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G141gat), .ZN(new_n222_));
  INV_X1    g021(.A(G148gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n221_), .A2(new_n224_), .A3(new_n209_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n216_), .A2(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(G113gat), .B(G120gat), .Z(new_n227_));
  XNOR2_X1  g026(.A(G127gat), .B(G134gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  XOR2_X1   g028(.A(G127gat), .B(G134gat), .Z(new_n230_));
  XNOR2_X1  g029(.A(G113gat), .B(G120gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n229_), .A2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT90), .B(KEYINPUT91), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n229_), .A2(new_n232_), .A3(new_n234_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n226_), .A2(new_n238_), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n216_), .A2(new_n236_), .A3(new_n225_), .A4(new_n237_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G225gat), .A2(G233gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT101), .ZN(new_n243_));
  AOI22_X1  g042(.A1(new_n216_), .A2(new_n225_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT4), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n243_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  AND4_X1   g045(.A1(new_n243_), .A2(new_n226_), .A3(new_n238_), .A4(new_n245_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n239_), .A2(KEYINPUT4), .A3(new_n240_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n241_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n242_), .B1(new_n248_), .B2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G1gat), .B(G29gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(G85gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT0), .B(G57gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n252_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n256_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n242_), .B(new_n258_), .C1(new_n248_), .C2(new_n251_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n257_), .A2(KEYINPUT106), .A3(new_n259_), .ZN(new_n260_));
  OR2_X1    g059(.A1(G197gat), .A2(G204gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G197gat), .A2(G204gat), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n261_), .A2(KEYINPUT21), .A3(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT21), .ZN(new_n264_));
  AND2_X1   g063(.A1(G197gat), .A2(G204gat), .ZN(new_n265_));
  NOR2_X1   g064(.A1(G197gat), .A2(G204gat), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n264_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G211gat), .B(G218gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n263_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  NOR3_X1   g068(.A1(new_n265_), .A2(new_n266_), .A3(new_n264_), .ZN(new_n270_));
  XOR2_X1   g069(.A(G211gat), .B(G218gat), .Z(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n269_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G169gat), .A2(G176gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G183gat), .A2(G190gat), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT23), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(G183gat), .ZN(new_n278_));
  INV_X1    g077(.A(G190gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n277_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT85), .ZN(new_n283_));
  INV_X1    g082(.A(G169gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n283_), .B1(new_n284_), .B2(KEYINPUT22), .ZN(new_n285_));
  INV_X1    g084(.A(G176gat), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT22), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n287_), .A2(KEYINPUT85), .A3(G169gat), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n285_), .A2(new_n286_), .A3(new_n288_), .ZN(new_n289_));
  OR2_X1    g088(.A1(KEYINPUT84), .A2(G169gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(KEYINPUT84), .A2(G169gat), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n287_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n274_), .B(new_n282_), .C1(new_n289_), .C2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT86), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n278_), .A2(KEYINPUT25), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT25), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(G183gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n279_), .A2(KEYINPUT26), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT26), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(G190gat), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n295_), .A2(new_n297_), .A3(new_n298_), .A4(new_n300_), .ZN(new_n301_));
  AND3_X1   g100(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n302_));
  AOI21_X1  g101(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n284_), .A2(new_n286_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n305_), .A2(KEYINPUT24), .A3(new_n274_), .ZN(new_n306_));
  OR3_X1    g105(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n301_), .A2(new_n304_), .A3(new_n306_), .A4(new_n307_), .ZN(new_n308_));
  AND3_X1   g107(.A1(new_n293_), .A2(new_n294_), .A3(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n294_), .B1(new_n293_), .B2(new_n308_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n273_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(KEYINPUT104), .B(KEYINPUT20), .Z(new_n312_));
  AND2_X1   g111(.A1(new_n269_), .A2(new_n272_), .ZN(new_n313_));
  AND3_X1   g112(.A1(new_n277_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n287_), .A2(G169gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n284_), .A2(KEYINPUT22), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n315_), .A2(new_n316_), .A3(new_n286_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n274_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n314_), .B1(new_n318_), .B2(KEYINPUT97), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT97), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n317_), .A2(new_n320_), .A3(new_n274_), .ZN(new_n321_));
  AND3_X1   g120(.A1(new_n304_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT96), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n299_), .A2(G190gat), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n279_), .A2(KEYINPUT26), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n323_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n295_), .A2(new_n297_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n298_), .A2(new_n300_), .A3(KEYINPUT96), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  AOI22_X1  g128(.A1(new_n319_), .A2(new_n321_), .B1(new_n322_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT105), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n313_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n318_), .A2(KEYINPUT97), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n333_), .A2(new_n282_), .A3(new_n321_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n322_), .A2(new_n329_), .ZN(new_n335_));
  AND3_X1   g134(.A1(new_n334_), .A2(new_n331_), .A3(new_n335_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n311_), .B(new_n312_), .C1(new_n332_), .C2(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(KEYINPUT19), .A2(G226gat), .A3(G233gat), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(KEYINPUT19), .B1(G226gat), .B2(G233gat), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NOR3_X1   g140(.A1(new_n309_), .A2(new_n310_), .A3(new_n273_), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT20), .B1(new_n330_), .B2(new_n313_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n341_), .B(KEYINPUT95), .Z(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n337_), .A2(new_n341_), .B1(new_n344_), .B2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n345_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n293_), .A2(new_n308_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT86), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n293_), .A2(new_n294_), .A3(new_n308_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n313_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n334_), .A2(new_n313_), .A3(new_n335_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT20), .B1(new_n339_), .B2(new_n340_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT98), .B1(new_n352_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT98), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n311_), .A2(new_n358_), .A3(new_n353_), .A4(new_n355_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n348_), .A2(new_n357_), .A3(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G64gat), .B(G92gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT100), .ZN(new_n362_));
  XOR2_X1   g161(.A(KEYINPUT99), .B(KEYINPUT18), .Z(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G8gat), .B(G36gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT32), .ZN(new_n367_));
  MUX2_X1   g166(.A(new_n347_), .B(new_n360_), .S(new_n367_), .Z(new_n368_));
  INV_X1    g167(.A(KEYINPUT106), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n252_), .A2(new_n369_), .A3(new_n256_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n260_), .A2(new_n368_), .A3(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n239_), .A2(new_n240_), .A3(new_n250_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(new_n256_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n249_), .A2(new_n241_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT101), .B1(new_n239_), .B2(KEYINPUT4), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n244_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n373_), .B1(new_n374_), .B2(new_n377_), .ZN(new_n378_));
  XOR2_X1   g177(.A(KEYINPUT103), .B(KEYINPUT33), .Z(new_n379_));
  AOI21_X1  g178(.A(new_n378_), .B1(new_n259_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT33), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT102), .B1(new_n259_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n366_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n360_), .A2(new_n383_), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n348_), .A2(new_n366_), .A3(new_n357_), .A4(new_n359_), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n242_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n249_), .A2(new_n250_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n387_), .B1(new_n388_), .B2(new_n377_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT102), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n389_), .A2(new_n390_), .A3(KEYINPUT33), .A4(new_n258_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n380_), .A2(new_n382_), .A3(new_n386_), .A4(new_n391_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n371_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G228gat), .A2(G233gat), .ZN(new_n394_));
  INV_X1    g193(.A(G78gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(G106gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G22gat), .B(G50gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  OR2_X1    g200(.A1(new_n226_), .A2(KEYINPUT29), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT28), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n313_), .B1(new_n226_), .B2(KEYINPUT29), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT28), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n402_), .B(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n404_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n401_), .B1(new_n405_), .B2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n403_), .A2(new_n404_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n407_), .A2(new_n408_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(new_n412_), .A3(new_n400_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n410_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n384_), .A2(new_n385_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT27), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  OAI211_X1 g216(.A(KEYINPUT27), .B(new_n385_), .C1(new_n347_), .C2(new_n366_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n260_), .A2(new_n370_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n414_), .ZN(new_n421_));
  OAI22_X1  g220(.A1(new_n393_), .A2(new_n414_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G227gat), .A2(G233gat), .ZN(new_n423_));
  INV_X1    g222(.A(G71gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(G99gat), .ZN(new_n426_));
  XOR2_X1   g225(.A(G15gat), .B(G43gat), .Z(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(KEYINPUT88), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n426_), .B(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(KEYINPUT87), .B(KEYINPUT30), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n431_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n350_), .A2(new_n351_), .A3(new_n430_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT89), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n429_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(KEYINPUT89), .B1(new_n432_), .B2(new_n433_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n238_), .B(KEYINPUT31), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  AOI211_X1 g240(.A(KEYINPUT89), .B(new_n429_), .C1(new_n433_), .C2(new_n432_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n439_), .A2(new_n441_), .A3(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n440_), .B1(new_n438_), .B2(new_n442_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n414_), .ZN(new_n448_));
  AOI22_X1  g247(.A1(new_n260_), .A2(new_n370_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n385_), .A2(KEYINPUT27), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n337_), .A2(new_n341_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n344_), .A2(new_n346_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n366_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n450_), .A2(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(KEYINPUT27), .B1(new_n384_), .B2(new_n385_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT107), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n454_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(KEYINPUT107), .B1(new_n417_), .B2(new_n418_), .ZN(new_n458_));
  OAI211_X1 g257(.A(new_n448_), .B(new_n449_), .C1(new_n457_), .C2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT108), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n417_), .A2(KEYINPUT107), .A3(new_n418_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n456_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n414_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n464_), .A2(KEYINPUT108), .A3(new_n449_), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n422_), .A2(new_n447_), .B1(new_n461_), .B2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G29gat), .B(G36gat), .ZN(new_n467_));
  OR2_X1    g266(.A1(new_n467_), .A2(KEYINPUT78), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(KEYINPUT78), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G43gat), .B(G50gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n468_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT15), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n473_), .A2(KEYINPUT15), .A3(new_n474_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G15gat), .B(G22gat), .ZN(new_n480_));
  INV_X1    g279(.A(G1gat), .ZN(new_n481_));
  INV_X1    g280(.A(G8gat), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT14), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n480_), .A2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G1gat), .B(G8gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n479_), .A2(new_n486_), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n475_), .A2(new_n486_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G229gat), .A2(G233gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n475_), .B(new_n486_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n489_), .ZN(new_n492_));
  AND3_X1   g291(.A1(new_n491_), .A2(KEYINPUT83), .A3(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(KEYINPUT83), .B1(new_n491_), .B2(new_n492_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n490_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G113gat), .B(G141gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G169gat), .B(G197gat), .ZN(new_n497_));
  XOR2_X1   g296(.A(new_n496_), .B(new_n497_), .Z(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n495_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n495_), .A2(new_n499_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n466_), .A2(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(G85gat), .B(G92gat), .Z(new_n505_));
  NOR2_X1   g304(.A1(G99gat), .A2(G106gat), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT7), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G99gat), .A2(G106gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT6), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT6), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n511_), .A2(G99gat), .A3(G106gat), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n505_), .B1(new_n508_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT8), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(KEYINPUT65), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n510_), .A2(new_n512_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT65), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n508_), .B1(new_n516_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT66), .ZN(new_n521_));
  OR2_X1    g320(.A1(new_n521_), .A2(KEYINPUT8), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(KEYINPUT8), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n505_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n515_), .B1(new_n520_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n516_), .A2(new_n519_), .ZN(new_n526_));
  XOR2_X1   g325(.A(KEYINPUT10), .B(G99gat), .Z(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n397_), .ZN(new_n528_));
  INV_X1    g327(.A(G85gat), .ZN(new_n529_));
  INV_X1    g328(.A(G92gat), .ZN(new_n530_));
  NOR3_X1   g329(.A1(new_n529_), .A2(new_n530_), .A3(KEYINPUT9), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n531_), .B1(new_n505_), .B2(KEYINPUT9), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n526_), .A2(new_n528_), .A3(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n525_), .A2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G57gat), .B(G64gat), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n535_), .A2(KEYINPUT11), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(KEYINPUT11), .ZN(new_n537_));
  XOR2_X1   g336(.A(G71gat), .B(G78gat), .Z(new_n538_));
  NAND3_X1  g337(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  OR2_X1    g338(.A1(new_n537_), .A2(new_n538_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n534_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT12), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n542_), .A2(KEYINPUT12), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT71), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n533_), .A2(new_n547_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n526_), .A2(KEYINPUT71), .A3(new_n528_), .A4(new_n532_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n548_), .A2(new_n525_), .A3(new_n549_), .ZN(new_n550_));
  AOI22_X1  g349(.A1(new_n543_), .A2(new_n544_), .B1(new_n546_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT72), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n525_), .A2(new_n541_), .A3(new_n533_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G230gat), .A2(G233gat), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n554_), .B(KEYINPUT64), .Z(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n552_), .B1(new_n553_), .B2(new_n556_), .ZN(new_n557_));
  AND3_X1   g356(.A1(new_n553_), .A2(new_n552_), .A3(new_n556_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n551_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G120gat), .B(G148gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G176gat), .B(G204gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(KEYINPUT73), .B(KEYINPUT5), .Z(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT69), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n543_), .B(new_n565_), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n553_), .A2(KEYINPUT67), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n553_), .A2(KEYINPUT67), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(KEYINPUT68), .A3(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT68), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n553_), .A2(KEYINPUT67), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n553_), .A2(KEYINPUT67), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n570_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n566_), .A2(new_n569_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT70), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n574_), .A2(new_n575_), .A3(new_n555_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n575_), .B1(new_n574_), .B2(new_n555_), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n559_), .B(new_n564_), .C1(new_n576_), .C2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n559_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n574_), .A2(new_n555_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT70), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n574_), .A2(new_n575_), .A3(new_n555_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n579_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n564_), .B(KEYINPUT74), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n578_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT75), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT13), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n586_), .A2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n559_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(new_n584_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(KEYINPUT75), .B(KEYINPUT13), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n592_), .A2(new_n578_), .A3(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n590_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n541_), .B(new_n486_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G231gat), .A2(G233gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(G127gat), .B(G155gat), .Z(new_n599_));
  XNOR2_X1  g398(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G183gat), .B(G211gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(KEYINPUT17), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n598_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n603_), .B(KEYINPUT17), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n606_), .B1(new_n598_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT80), .ZN(new_n609_));
  XNOR2_X1  g408(.A(KEYINPUT76), .B(KEYINPUT34), .ZN(new_n610_));
  AND2_X1   g409(.A1(G232gat), .A2(G233gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n612_), .A2(KEYINPUT35), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n613_), .B1(new_n479_), .B2(new_n550_), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n534_), .A2(new_n475_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n612_), .A2(KEYINPUT35), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT77), .Z(new_n618_));
  NAND2_X1  g417(.A1(new_n479_), .A2(new_n550_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n618_), .B1(new_n619_), .B2(KEYINPUT79), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n616_), .A2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G190gat), .B(G218gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G134gat), .B(G162gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n624_), .A2(KEYINPUT36), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT79), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n626_), .B1(new_n479_), .B2(new_n550_), .ZN(new_n627_));
  OAI211_X1 g426(.A(new_n614_), .B(new_n615_), .C1(new_n627_), .C2(new_n618_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n621_), .A2(new_n625_), .A3(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n624_), .B(KEYINPUT36), .Z(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n632_), .B1(new_n621_), .B2(new_n628_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n630_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT37), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n609_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  OAI211_X1 g435(.A(KEYINPUT80), .B(KEYINPUT37), .C1(new_n630_), .C2(new_n633_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT81), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n634_), .A2(new_n639_), .A3(new_n635_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n633_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n641_), .A2(new_n635_), .A3(new_n629_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT81), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n638_), .A2(new_n644_), .ZN(new_n645_));
  AND4_X1   g444(.A1(new_n504_), .A2(new_n595_), .A3(new_n608_), .A4(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n420_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n646_), .A2(new_n481_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT38), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n466_), .A2(new_n634_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n608_), .ZN(new_n652_));
  AOI211_X1 g451(.A(new_n503_), .B(new_n652_), .C1(new_n590_), .C2(new_n594_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(G1gat), .B1(new_n654_), .B2(new_n420_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n648_), .A2(new_n649_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n650_), .A2(new_n655_), .A3(new_n656_), .ZN(G1324gat));
  NAND2_X1  g456(.A1(new_n462_), .A2(new_n463_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n646_), .A2(new_n482_), .A3(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(G8gat), .B1(new_n654_), .B2(new_n658_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT109), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT39), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT109), .ZN(new_n664_));
  OAI211_X1 g463(.A(new_n664_), .B(G8gat), .C1(new_n654_), .C2(new_n658_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n662_), .A2(new_n663_), .A3(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n663_), .B1(new_n662_), .B2(new_n665_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n660_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT40), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  OAI211_X1 g469(.A(KEYINPUT40), .B(new_n660_), .C1(new_n666_), .C2(new_n667_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1325gat));
  INV_X1    g471(.A(G15gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n646_), .A2(new_n673_), .A3(new_n446_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT110), .Z(new_n675_));
  OAI21_X1  g474(.A(G15gat), .B1(new_n654_), .B2(new_n447_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT41), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n676_), .A2(KEYINPUT41), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n675_), .A2(new_n677_), .A3(new_n678_), .ZN(G1326gat));
  OAI21_X1  g478(.A(G22gat), .B1(new_n654_), .B2(new_n448_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT42), .ZN(new_n681_));
  INV_X1    g480(.A(G22gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n646_), .A2(new_n682_), .A3(new_n414_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(G1327gat));
  NAND2_X1  g483(.A1(new_n461_), .A2(new_n465_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n421_), .A2(new_n419_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n414_), .B1(new_n371_), .B2(new_n392_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n447_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n645_), .B1(new_n685_), .B2(new_n688_), .ZN(new_n689_));
  OAI211_X1 g488(.A(KEYINPUT112), .B(KEYINPUT43), .C1(new_n689_), .C2(KEYINPUT111), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n590_), .A2(new_n594_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n691_), .A2(new_n503_), .A3(new_n608_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT112), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n459_), .A2(new_n460_), .ZN(new_n694_));
  AOI21_X1  g493(.A(KEYINPUT108), .B1(new_n464_), .B2(new_n449_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n688_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n645_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT111), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n693_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n701_), .B1(new_n689_), .B2(KEYINPUT112), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n690_), .B(new_n692_), .C1(new_n700_), .C2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(KEYINPUT43), .B1(new_n698_), .B2(new_n693_), .ZN(new_n706_));
  OAI21_X1  g505(.A(KEYINPUT112), .B1(new_n689_), .B2(KEYINPUT111), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n708_), .A2(KEYINPUT44), .A3(new_n690_), .A4(new_n692_), .ZN(new_n709_));
  AND4_X1   g508(.A1(G29gat), .A2(new_n705_), .A3(new_n647_), .A4(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n634_), .A2(new_n652_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n691_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n504_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(G29gat), .B1(new_n714_), .B2(new_n647_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n710_), .A2(new_n715_), .ZN(G1328gat));
  NAND3_X1  g515(.A1(new_n705_), .A2(new_n659_), .A3(new_n709_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(G36gat), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n713_), .A2(G36gat), .A3(new_n658_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT45), .Z(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT46), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n718_), .A2(new_n720_), .A3(KEYINPUT46), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(G1329gat));
  NAND4_X1  g524(.A1(new_n705_), .A2(new_n709_), .A3(G43gat), .A4(new_n446_), .ZN(new_n726_));
  INV_X1    g525(.A(G43gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n727_), .B1(new_n713_), .B2(new_n447_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT47), .ZN(G1330gat));
  AND4_X1   g529(.A1(G50gat), .A2(new_n705_), .A3(new_n414_), .A4(new_n709_), .ZN(new_n731_));
  AOI21_X1  g530(.A(G50gat), .B1(new_n714_), .B2(new_n414_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1331gat));
  NAND4_X1  g532(.A1(new_n651_), .A2(new_n503_), .A3(new_n691_), .A4(new_n608_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT113), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n735_), .A2(G57gat), .A3(new_n647_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n736_), .A2(KEYINPUT114), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n736_), .A2(KEYINPUT114), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n595_), .A2(new_n697_), .A3(new_n652_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n466_), .A2(new_n502_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(G57gat), .B1(new_n742_), .B2(new_n647_), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n737_), .A2(new_n738_), .A3(new_n743_), .ZN(G1332gat));
  OR3_X1    g543(.A1(new_n741_), .A2(G64gat), .A3(new_n658_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n735_), .A2(new_n659_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(KEYINPUT115), .B(KEYINPUT48), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n746_), .A2(G64gat), .A3(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n746_), .B2(G64gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n745_), .B1(new_n748_), .B2(new_n749_), .ZN(G1333gat));
  NAND3_X1  g549(.A1(new_n742_), .A2(new_n424_), .A3(new_n446_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT49), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n735_), .A2(new_n446_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n753_), .B2(G71gat), .ZN(new_n754_));
  AOI211_X1 g553(.A(KEYINPUT49), .B(new_n424_), .C1(new_n735_), .C2(new_n446_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(G1334gat));
  INV_X1    g555(.A(KEYINPUT50), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n735_), .A2(new_n414_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n758_), .B2(G78gat), .ZN(new_n759_));
  AOI211_X1 g558(.A(KEYINPUT50), .B(new_n395_), .C1(new_n735_), .C2(new_n414_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n414_), .A2(new_n395_), .ZN(new_n761_));
  XOR2_X1   g560(.A(new_n761_), .B(KEYINPUT116), .Z(new_n762_));
  OAI22_X1  g561(.A1(new_n759_), .A2(new_n760_), .B1(new_n741_), .B2(new_n762_), .ZN(G1335gat));
  NOR4_X1   g562(.A1(new_n466_), .A2(new_n595_), .A3(new_n502_), .A4(new_n711_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n764_), .A2(new_n529_), .A3(new_n647_), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n595_), .A2(new_n502_), .A3(new_n608_), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n690_), .B(new_n766_), .C1(new_n700_), .C2(new_n702_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT117), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT117), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n708_), .A2(new_n769_), .A3(new_n690_), .A4(new_n766_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n420_), .B1(new_n768_), .B2(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n765_), .B1(new_n771_), .B2(new_n529_), .ZN(G1336gat));
  NAND3_X1  g571(.A1(new_n764_), .A2(new_n530_), .A3(new_n659_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n658_), .B1(new_n768_), .B2(new_n770_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(new_n774_), .B2(new_n530_), .ZN(G1337gat));
  NAND3_X1  g574(.A1(new_n764_), .A2(new_n446_), .A3(new_n527_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n447_), .B1(new_n768_), .B2(new_n770_), .ZN(new_n777_));
  INV_X1    g576(.A(G99gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n776_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT51), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n781_), .B(new_n776_), .C1(new_n777_), .C2(new_n778_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(G1338gat));
  NAND3_X1  g582(.A1(new_n764_), .A2(new_n397_), .A3(new_n414_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n708_), .A2(new_n414_), .A3(new_n690_), .A4(new_n766_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n785_), .A2(new_n786_), .A3(G106gat), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n785_), .B2(G106gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n784_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT53), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n791_), .B(new_n784_), .C1(new_n787_), .C2(new_n788_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(G1339gat));
  OAI21_X1  g592(.A(KEYINPUT118), .B1(new_n502_), .B2(new_n652_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT118), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n500_), .A2(new_n608_), .A3(new_n795_), .A4(new_n501_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n797_), .B1(new_n638_), .B2(new_n644_), .ZN(new_n798_));
  AOI211_X1 g597(.A(KEYINPUT119), .B(KEYINPUT54), .C1(new_n595_), .C2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n595_), .A2(new_n798_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT119), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n800_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n595_), .A2(KEYINPUT119), .A3(new_n798_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n799_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT121), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n559_), .A2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n551_), .A2(new_n568_), .A3(new_n567_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n555_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n551_), .B(KEYINPUT55), .C1(new_n557_), .C2(new_n558_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n808_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n584_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT56), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n812_), .A2(KEYINPUT56), .A3(new_n584_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n487_), .A2(new_n488_), .A3(new_n492_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n498_), .B1(new_n491_), .B2(new_n489_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  OR2_X1    g619(.A1(new_n820_), .A2(KEYINPUT120), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(KEYINPUT120), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n500_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n578_), .A2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n806_), .B1(new_n817_), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT58), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT58), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n806_), .B(new_n827_), .C1(new_n817_), .C2(new_n824_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n826_), .A2(new_n697_), .A3(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n815_), .A2(new_n816_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n503_), .B1(new_n583_), .B2(new_n564_), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n831_), .A2(new_n832_), .B1(new_n586_), .B2(new_n823_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n830_), .B1(new_n833_), .B2(new_n634_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n586_), .A2(new_n823_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n831_), .A2(new_n502_), .A3(new_n578_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n634_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(KEYINPUT57), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n829_), .A2(new_n834_), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n652_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n805_), .A2(new_n840_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n464_), .A2(new_n446_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n841_), .A2(new_n647_), .A3(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(G113gat), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(new_n845_), .A3(new_n502_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT59), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT122), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n841_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n843_), .A2(new_n847_), .A3(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n420_), .B1(new_n805_), .B2(new_n840_), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT122), .B1(new_n805_), .B2(new_n840_), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n851_), .B(new_n842_), .C1(new_n852_), .C2(KEYINPUT59), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n503_), .B1(new_n850_), .B2(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n846_), .B1(new_n854_), .B2(new_n845_), .ZN(G1340gat));
  INV_X1    g654(.A(G120gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n856_), .B1(new_n595_), .B2(KEYINPUT60), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n844_), .B(new_n857_), .C1(KEYINPUT60), .C2(new_n856_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n595_), .B1(new_n850_), .B2(new_n853_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n859_), .B2(new_n856_), .ZN(G1341gat));
  AOI21_X1  g659(.A(G127gat), .B1(new_n844_), .B2(new_n608_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n850_), .A2(new_n853_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT123), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(G127gat), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n608_), .A2(KEYINPUT123), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(G127gat), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n861_), .B1(new_n862_), .B2(new_n866_), .ZN(G1342gat));
  INV_X1    g666(.A(G134gat), .ZN(new_n868_));
  INV_X1    g667(.A(new_n634_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n843_), .B2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(KEYINPUT124), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT124), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n872_), .B(new_n868_), .C1(new_n843_), .C2(new_n869_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n645_), .A2(new_n868_), .ZN(new_n874_));
  AOI22_X1  g673(.A1(new_n871_), .A2(new_n873_), .B1(new_n862_), .B2(new_n874_), .ZN(G1343gat));
  NOR3_X1   g674(.A1(new_n659_), .A2(new_n448_), .A3(new_n446_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n851_), .A2(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(new_n503_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(new_n222_), .ZN(G1344gat));
  NOR2_X1   g678(.A1(new_n877_), .A2(new_n595_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(new_n223_), .ZN(G1345gat));
  NAND3_X1  g680(.A1(new_n851_), .A2(new_n608_), .A3(new_n876_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT61), .B(G155gat), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1346gat));
  OAI21_X1  g683(.A(G162gat), .B1(new_n877_), .B2(new_n645_), .ZN(new_n885_));
  OR2_X1    g684(.A1(new_n869_), .A2(G162gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n877_), .B2(new_n886_), .ZN(G1347gat));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n448_), .A2(new_n449_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n837_), .B(new_n830_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n608_), .B1(new_n891_), .B2(new_n829_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n801_), .A2(new_n802_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n893_), .A2(KEYINPUT54), .A3(new_n804_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n799_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n659_), .B(new_n890_), .C1(new_n892_), .C2(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n503_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n888_), .B1(new_n898_), .B2(new_n284_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n898_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n900_));
  OAI211_X1 g699(.A(KEYINPUT62), .B(G169gat), .C1(new_n897_), .C2(new_n503_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n899_), .A2(new_n900_), .A3(new_n901_), .ZN(G1348gat));
  NOR2_X1   g701(.A1(new_n897_), .A2(new_n595_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(new_n286_), .ZN(G1349gat));
  OAI21_X1  g703(.A(KEYINPUT126), .B1(new_n897_), .B2(new_n652_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n658_), .B1(new_n805_), .B2(new_n840_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT126), .ZN(new_n907_));
  NAND4_X1  g706(.A1(new_n906_), .A2(new_n907_), .A3(new_n608_), .A4(new_n890_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n905_), .A2(new_n278_), .A3(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n327_), .ZN(new_n910_));
  NAND4_X1  g709(.A1(new_n906_), .A2(new_n910_), .A3(new_n608_), .A4(new_n890_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(KEYINPUT125), .ZN(new_n912_));
  INV_X1    g711(.A(new_n897_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT125), .ZN(new_n914_));
  NAND4_X1  g713(.A1(new_n913_), .A2(new_n914_), .A3(new_n910_), .A4(new_n608_), .ZN(new_n915_));
  AND3_X1   g714(.A1(new_n909_), .A2(new_n912_), .A3(new_n915_), .ZN(G1350gat));
  OAI21_X1  g715(.A(G190gat), .B1(new_n897_), .B2(new_n645_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n634_), .A2(new_n326_), .A3(new_n328_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n897_), .B2(new_n918_), .ZN(G1351gat));
  NOR2_X1   g718(.A1(new_n421_), .A2(new_n446_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n906_), .A2(new_n502_), .A3(new_n920_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g721(.A1(new_n906_), .A2(new_n920_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n923_), .A2(new_n595_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n924_), .B(new_n925_), .ZN(G1353gat));
  XNOR2_X1  g725(.A(KEYINPUT63), .B(G211gat), .ZN(new_n927_));
  OR2_X1    g726(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n906_), .A2(new_n608_), .A3(new_n920_), .ZN(new_n929_));
  MUX2_X1   g728(.A(new_n927_), .B(new_n928_), .S(new_n929_), .Z(G1354gat));
  OAI21_X1  g729(.A(G218gat), .B1(new_n923_), .B2(new_n645_), .ZN(new_n931_));
  OR2_X1    g730(.A1(new_n869_), .A2(G218gat), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n923_), .B2(new_n932_), .ZN(G1355gat));
endmodule


