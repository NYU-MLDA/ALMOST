//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 1 0 0 0 0 0 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 0 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n818_, new_n819_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n834_,
    new_n835_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n883_, new_n884_, new_n885_, new_n887_, new_n888_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT31), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT83), .ZN(new_n206_));
  NOR2_X1   g005(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(G169gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT80), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n209_), .B1(new_n210_), .B2(KEYINPUT23), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(KEYINPUT23), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G183gat), .A3(G190gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n211_), .B1(new_n215_), .B2(new_n209_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n208_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT26), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT78), .B1(new_n219_), .B2(G190gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT25), .B(G183gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(KEYINPUT26), .B(G190gat), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n220_), .B(new_n221_), .C1(new_n222_), .C2(KEYINPUT78), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n226_));
  OR3_X1    g025(.A1(new_n225_), .A2(new_n226_), .A3(KEYINPUT79), .ZN(new_n227_));
  NOR3_X1   g026(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n228_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT79), .B1(new_n225_), .B2(new_n226_), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n223_), .A2(new_n227_), .A3(new_n229_), .A4(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n218_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT30), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT82), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n234_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G227gat), .A2(G233gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT81), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G71gat), .B(G99gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(G15gat), .B(G43gat), .Z(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n235_), .A2(new_n236_), .A3(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n236_), .A2(new_n242_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n206_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n205_), .B1(new_n245_), .B2(KEYINPUT84), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT83), .B1(new_n205_), .B2(KEYINPUT84), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n243_), .A2(new_n247_), .A3(new_n244_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  OR2_X1    g049(.A1(G155gat), .A2(G162gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G155gat), .A2(G162gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G141gat), .A2(G148gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT2), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n256_));
  INV_X1    g055(.A(G141gat), .ZN(new_n257_));
  INV_X1    g056(.A(G148gat), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n256_), .A2(new_n257_), .A3(new_n258_), .A4(KEYINPUT85), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT85), .ZN(new_n260_));
  OAI22_X1  g059(.A1(new_n260_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n251_), .B(new_n252_), .C1(new_n255_), .C2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n257_), .A2(new_n258_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n252_), .A2(KEYINPUT1), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(new_n251_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n252_), .A2(KEYINPUT1), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n264_), .B(new_n253_), .C1(new_n266_), .C2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n204_), .A2(new_n263_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n204_), .B1(new_n263_), .B2(new_n268_), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT97), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G225gat), .A2(G233gat), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n263_), .A2(new_n268_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n204_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT97), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(new_n278_), .A3(new_n269_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n272_), .A2(new_n274_), .A3(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n277_), .A2(KEYINPUT4), .A3(new_n269_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n271_), .A2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n281_), .A2(new_n273_), .A3(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G1gat), .B(G29gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(G85gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT0), .B(G57gat), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n286_), .B(new_n287_), .Z(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  AND3_X1   g088(.A1(new_n280_), .A2(new_n284_), .A3(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n273_), .B1(new_n281_), .B2(new_n283_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n274_), .B1(new_n277_), .B2(new_n269_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n288_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(KEYINPUT96), .A2(KEYINPUT33), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n288_), .B(new_n294_), .C1(new_n291_), .C2(new_n292_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n290_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n215_), .B1(G183gat), .B2(G190gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(new_n208_), .ZN(new_n300_));
  INV_X1    g099(.A(G183gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT25), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT25), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(G183gat), .ZN(new_n304_));
  AND3_X1   g103(.A1(new_n302_), .A2(new_n304_), .A3(KEYINPUT92), .ZN(new_n305_));
  AOI21_X1  g104(.A(KEYINPUT92), .B1(new_n302_), .B2(new_n304_), .ZN(new_n306_));
  XOR2_X1   g105(.A(KEYINPUT26), .B(G190gat), .Z(new_n307_));
  NOR3_X1   g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n226_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n228_), .B1(new_n309_), .B2(new_n224_), .ZN(new_n310_));
  AOI21_X1  g109(.A(KEYINPUT80), .B1(new_n212_), .B2(new_n214_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n310_), .B1(new_n311_), .B2(new_n211_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n300_), .B1(new_n308_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(G211gat), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n314_), .A2(G218gat), .ZN(new_n315_));
  INV_X1    g114(.A(G218gat), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n316_), .A2(G211gat), .ZN(new_n317_));
  NOR2_X1   g116(.A1(G197gat), .A2(G204gat), .ZN(new_n318_));
  AND2_X1   g117(.A1(G197gat), .A2(G204gat), .ZN(new_n319_));
  OAI22_X1  g118(.A1(new_n315_), .A2(new_n317_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G211gat), .B(G218gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT87), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n322_), .B1(new_n319_), .B2(new_n318_), .ZN(new_n323_));
  AOI22_X1  g122(.A1(new_n320_), .A2(KEYINPUT21), .B1(new_n321_), .B2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n323_), .A2(KEYINPUT21), .A3(new_n321_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT94), .B1(new_n313_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G226gat), .A2(G233gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(KEYINPUT19), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT20), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n328_), .A2(new_n332_), .ZN(new_n333_));
  OR3_X1    g132(.A1(new_n313_), .A2(new_n327_), .A3(KEYINPUT94), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT93), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT88), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n336_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT21), .ZN(new_n338_));
  INV_X1    g137(.A(new_n321_), .ZN(new_n339_));
  OR2_X1    g138(.A1(new_n319_), .A2(new_n318_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n338_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n323_), .A2(new_n321_), .ZN(new_n342_));
  OAI211_X1 g141(.A(KEYINPUT88), .B(new_n325_), .C1(new_n341_), .C2(new_n342_), .ZN(new_n343_));
  AOI221_X4 g142(.A(new_n335_), .B1(new_n218_), .B2(new_n231_), .C1(new_n337_), .C2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n337_), .A2(new_n343_), .ZN(new_n345_));
  AOI21_X1  g144(.A(KEYINPUT93), .B1(new_n345_), .B2(new_n232_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n333_), .B(new_n334_), .C1(new_n344_), .C2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n331_), .B1(new_n313_), .B2(new_n327_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n348_), .B1(new_n232_), .B2(new_n345_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n330_), .B(KEYINPUT91), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  XOR2_X1   g150(.A(G8gat), .B(G36gat), .Z(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT18), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G64gat), .B(G92gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n347_), .A2(KEYINPUT95), .A3(new_n351_), .A4(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n344_), .A2(new_n346_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n334_), .A2(new_n328_), .A3(new_n332_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n351_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n355_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n351_), .B(new_n355_), .C1(new_n357_), .C2(new_n358_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT95), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n298_), .A2(new_n356_), .A3(new_n361_), .A4(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT98), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n355_), .B1(new_n347_), .B2(new_n351_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n368_), .B1(new_n363_), .B2(new_n362_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n369_), .A2(KEYINPUT98), .A3(new_n356_), .A4(new_n298_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n355_), .A2(KEYINPUT32), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n359_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n327_), .ZN(new_n374_));
  OR2_X1    g173(.A1(new_n308_), .A2(new_n312_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n374_), .A2(new_n375_), .A3(new_n300_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT20), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n330_), .B1(new_n357_), .B2(new_n377_), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n349_), .A2(new_n350_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n373_), .B1(new_n380_), .B2(new_n372_), .ZN(new_n381_));
  OR3_X1    g180(.A1(new_n291_), .A2(new_n288_), .A3(new_n292_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n382_), .A2(KEYINPUT99), .A3(new_n293_), .ZN(new_n383_));
  OR4_X1    g182(.A1(KEYINPUT99), .A2(new_n291_), .A3(new_n288_), .A4(new_n292_), .ZN(new_n384_));
  AND2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n381_), .A2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n367_), .A2(new_n370_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n275_), .A2(KEYINPUT29), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT86), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G228gat), .A2(G233gat), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n275_), .A2(KEYINPUT86), .A3(KEYINPUT29), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n390_), .A2(new_n391_), .A3(new_n392_), .A4(new_n345_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n388_), .A2(new_n327_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n394_), .A2(G228gat), .A3(G233gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT90), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT90), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n393_), .A2(new_n398_), .A3(new_n395_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G78gat), .B(G106gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT89), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT28), .B1(new_n275_), .B2(KEYINPUT29), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NOR3_X1   g203(.A1(new_n275_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G22gat), .B(G50gat), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NOR3_X1   g206(.A1(new_n404_), .A2(new_n405_), .A3(new_n407_), .ZN(new_n408_));
  OR3_X1    g207(.A1(new_n275_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n406_), .B1(new_n409_), .B2(new_n403_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n402_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n407_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n409_), .A2(new_n403_), .A3(new_n406_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n402_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n412_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n411_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n400_), .A2(new_n416_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n397_), .A2(new_n411_), .A3(new_n399_), .A4(new_n415_), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n387_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n417_), .A2(new_n418_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n383_), .A2(new_n384_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n364_), .A2(new_n356_), .A3(new_n361_), .ZN(new_n425_));
  XOR2_X1   g224(.A(KEYINPUT100), .B(KEYINPUT27), .Z(new_n426_));
  NAND2_X1  g225(.A1(new_n380_), .A2(new_n360_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n362_), .A2(KEYINPUT27), .ZN(new_n428_));
  AOI22_X1  g227(.A1(new_n425_), .A2(new_n426_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n424_), .A2(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n250_), .B1(new_n420_), .B2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n246_), .A2(new_n248_), .A3(new_n422_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT101), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n425_), .A2(new_n426_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n427_), .A2(new_n428_), .ZN(new_n436_));
  AND4_X1   g235(.A1(new_n434_), .A2(new_n435_), .A3(new_n419_), .A4(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n434_), .B1(new_n429_), .B2(new_n419_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n433_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT102), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n435_), .A2(new_n419_), .A3(new_n436_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT101), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n429_), .A2(new_n434_), .A3(new_n419_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT102), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n444_), .A2(new_n445_), .A3(new_n433_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n431_), .B1(new_n440_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(G1gat), .ZN(new_n448_));
  INV_X1    g247(.A(G8gat), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT14), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT73), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  OAI211_X1 g251(.A(KEYINPUT73), .B(KEYINPUT14), .C1(new_n448_), .C2(new_n449_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G15gat), .B(G22gat), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT74), .ZN(new_n456_));
  XOR2_X1   g255(.A(G1gat), .B(G8gat), .Z(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G29gat), .B(G36gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G43gat), .B(G50gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  XOR2_X1   g260(.A(new_n461_), .B(KEYINPUT76), .Z(new_n462_));
  XNOR2_X1  g261(.A(new_n458_), .B(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G229gat), .A2(G233gat), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n461_), .B(KEYINPUT15), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  OR2_X1    g267(.A1(new_n458_), .A2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n465_), .B1(new_n458_), .B2(new_n462_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G113gat), .B(G141gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(KEYINPUT77), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G169gat), .B(G197gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n466_), .A2(new_n471_), .A3(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n475_), .B1(new_n466_), .B2(new_n471_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n447_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT72), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G232gat), .A2(G233gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT34), .ZN(new_n482_));
  NAND3_X1  g281(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT66), .B(G92gat), .ZN(new_n484_));
  INV_X1    g283(.A(G85gat), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  OAI22_X1  g285(.A1(KEYINPUT65), .A2(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n487_), .B1(KEYINPUT65), .B2(KEYINPUT9), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n483_), .B1(new_n486_), .B2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT6), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n490_), .B1(G99gat), .B2(G106gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G99gat), .A2(G106gat), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n492_), .A2(KEYINPUT6), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(KEYINPUT10), .B(G99gat), .Z(new_n495_));
  XOR2_X1   g294(.A(KEYINPUT64), .B(G106gat), .Z(new_n496_));
  AOI21_X1  g295(.A(new_n494_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n489_), .A2(new_n497_), .ZN(new_n498_));
  OR3_X1    g297(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n499_), .B(new_n500_), .C1(new_n491_), .C2(new_n493_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT8), .ZN(new_n502_));
  XOR2_X1   g301(.A(G85gat), .B(G92gat), .Z(new_n503_));
  NAND3_X1  g302(.A1(new_n501_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n502_), .B1(new_n501_), .B2(new_n503_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n498_), .B(KEYINPUT67), .C1(new_n505_), .C2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n501_), .A2(new_n503_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT8), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(new_n504_), .ZN(new_n511_));
  AOI21_X1  g310(.A(KEYINPUT67), .B1(new_n511_), .B2(new_n498_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n508_), .A2(new_n512_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n513_), .A2(new_n461_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n498_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n467_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT69), .ZN(new_n517_));
  OAI211_X1 g316(.A(KEYINPUT35), .B(new_n482_), .C1(new_n514_), .C2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n513_), .A2(new_n461_), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n482_), .B(KEYINPUT35), .Z(new_n520_));
  NAND3_X1  g319(.A1(new_n519_), .A2(new_n516_), .A3(new_n520_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n518_), .A2(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(G190gat), .B(G218gat), .Z(new_n523_));
  XNOR2_X1  g322(.A(G134gat), .B(G162gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT36), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n480_), .B1(new_n522_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n518_), .A2(new_n521_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n529_), .A2(KEYINPUT72), .A3(new_n526_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT36), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n525_), .A2(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n533_), .B(KEYINPUT70), .Z(new_n534_));
  NAND3_X1  g333(.A1(new_n518_), .A2(new_n521_), .A3(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT71), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n531_), .A2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT37), .B1(new_n522_), .B2(new_n527_), .ZN(new_n538_));
  OAI22_X1  g337(.A1(new_n537_), .A2(KEYINPUT37), .B1(new_n536_), .B2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G57gat), .B(G64gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT11), .ZN(new_n541_));
  XOR2_X1   g340(.A(G71gat), .B(G78gat), .Z(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n540_), .A2(KEYINPUT11), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n541_), .A2(new_n542_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n548_), .B1(new_n508_), .B2(new_n512_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT67), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n515_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n551_), .A2(new_n507_), .A3(new_n547_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n549_), .A2(KEYINPUT68), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G230gat), .A2(G233gat), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n553_), .B(new_n555_), .C1(KEYINPUT68), .C2(new_n552_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT12), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n548_), .A2(KEYINPUT12), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  AOI22_X1  g358(.A1(new_n549_), .A2(new_n557_), .B1(new_n559_), .B2(new_n515_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n555_), .B1(new_n513_), .B2(new_n547_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n556_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G120gat), .B(G148gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT5), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G176gat), .B(G204gat), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n565_), .B(new_n566_), .Z(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n563_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n556_), .A2(new_n562_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(new_n567_), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n569_), .A2(KEYINPUT13), .A3(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(KEYINPUT13), .B1(new_n569_), .B2(new_n571_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G231gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n547_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(new_n458_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT75), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G127gat), .B(G155gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT16), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G183gat), .B(G211gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT17), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n579_), .B(new_n584_), .ZN(new_n585_));
  OR3_X1    g384(.A1(new_n578_), .A2(KEYINPUT17), .A3(new_n583_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NOR3_X1   g387(.A1(new_n539_), .A2(new_n575_), .A3(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n479_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n590_), .A2(new_n448_), .A3(new_n385_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT38), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n478_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n574_), .A2(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n595_), .A2(new_n588_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT103), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT71), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n535_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n535_), .A2(new_n598_), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n528_), .B(new_n530_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT104), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n447_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n597_), .A2(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(G1gat), .B1(new_n606_), .B2(new_n422_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n591_), .A2(new_n592_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n593_), .A2(new_n607_), .A3(new_n608_), .ZN(G1324gat));
  INV_X1    g408(.A(new_n429_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n590_), .A2(new_n449_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT39), .ZN(new_n612_));
  INV_X1    g411(.A(new_n606_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n610_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n612_), .B1(new_n614_), .B2(G8gat), .ZN(new_n615_));
  AOI211_X1 g414(.A(KEYINPUT39), .B(new_n449_), .C1(new_n613_), .C2(new_n610_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n611_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g417(.A(G15gat), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n590_), .A2(new_n619_), .A3(new_n250_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n613_), .A2(new_n250_), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n621_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n622_));
  AOI21_X1  g421(.A(KEYINPUT41), .B1(new_n621_), .B2(G15gat), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n620_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT105), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(G1326gat));
  OAI21_X1  g425(.A(G22gat), .B1(new_n606_), .B2(new_n419_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT42), .ZN(new_n628_));
  INV_X1    g427(.A(G22gat), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n590_), .A2(new_n629_), .A3(new_n421_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(G1327gat));
  NOR2_X1   g430(.A1(new_n602_), .A2(new_n587_), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n479_), .A2(new_n574_), .A3(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(G29gat), .B1(new_n633_), .B2(new_n385_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n595_), .A2(new_n587_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n601_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n538_), .B1(new_n636_), .B2(new_n599_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT37), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n638_), .B2(new_n602_), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n447_), .A2(KEYINPUT43), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT43), .ZN(new_n641_));
  AOI22_X1  g440(.A1(new_n365_), .A2(new_n366_), .B1(new_n381_), .B2(new_n385_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n421_), .B1(new_n642_), .B2(new_n370_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n430_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n249_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n445_), .B1(new_n444_), .B2(new_n433_), .ZN(new_n646_));
  AOI211_X1 g445(.A(KEYINPUT102), .B(new_n432_), .C1(new_n442_), .C2(new_n443_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n645_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n641_), .B1(new_n648_), .B2(new_n539_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n635_), .B1(new_n640_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT44), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  OAI211_X1 g451(.A(KEYINPUT44), .B(new_n635_), .C1(new_n640_), .C2(new_n649_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n385_), .A2(G29gat), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n634_), .B1(new_n655_), .B2(new_n656_), .ZN(G1328gat));
  INV_X1    g456(.A(G36gat), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n633_), .A2(new_n658_), .A3(new_n610_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT45), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n652_), .A2(new_n610_), .A3(new_n653_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n661_), .A2(KEYINPUT106), .A3(G36gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT106), .B1(new_n661_), .B2(G36gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n660_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT46), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  OAI211_X1 g465(.A(KEYINPUT46), .B(new_n660_), .C1(new_n662_), .C2(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1329gat));
  NAND2_X1  g467(.A1(new_n250_), .A2(G43gat), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n633_), .A2(new_n250_), .ZN(new_n670_));
  OAI22_X1  g469(.A1(new_n654_), .A2(new_n669_), .B1(G43gat), .B2(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n671_), .B(new_n672_), .Z(G1330gat));
  AOI21_X1  g472(.A(G50gat), .B1(new_n633_), .B2(new_n421_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n421_), .A2(G50gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n655_), .B2(new_n675_), .ZN(G1331gat));
  NAND3_X1  g475(.A1(new_n639_), .A2(new_n575_), .A3(new_n587_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT108), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n447_), .A2(new_n594_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(G57gat), .B1(new_n681_), .B2(new_n385_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n575_), .A2(new_n478_), .ZN(new_n683_));
  NOR4_X1   g482(.A1(new_n447_), .A2(new_n604_), .A3(new_n588_), .A4(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(G57gat), .A3(new_n385_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT109), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n685_), .A2(new_n686_), .ZN(new_n688_));
  NOR3_X1   g487(.A1(new_n682_), .A2(new_n687_), .A3(new_n688_), .ZN(G1332gat));
  INV_X1    g488(.A(G64gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n690_), .B1(new_n684_), .B2(new_n610_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT48), .Z(new_n692_));
  NAND3_X1  g491(.A1(new_n681_), .A2(new_n690_), .A3(new_n610_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1333gat));
  INV_X1    g493(.A(G71gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n695_), .B1(new_n684_), .B2(new_n250_), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT49), .Z(new_n697_));
  NAND3_X1  g496(.A1(new_n681_), .A2(new_n695_), .A3(new_n250_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(G1334gat));
  INV_X1    g498(.A(G78gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n700_), .B1(new_n684_), .B2(new_n421_), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT50), .Z(new_n702_));
  NAND3_X1  g501(.A1(new_n681_), .A2(new_n700_), .A3(new_n421_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1335gat));
  NAND3_X1  g503(.A1(new_n679_), .A2(new_n575_), .A3(new_n632_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT110), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n706_), .A2(new_n485_), .A3(new_n385_), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n640_), .A2(new_n649_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n683_), .A2(new_n587_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(G85gat), .B1(new_n710_), .B2(new_n422_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n707_), .A2(new_n711_), .ZN(G1336gat));
  AOI21_X1  g511(.A(G92gat), .B1(new_n706_), .B2(new_n610_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n429_), .A2(new_n484_), .ZN(new_n714_));
  XOR2_X1   g513(.A(new_n714_), .B(KEYINPUT111), .Z(new_n715_));
  NOR2_X1   g514(.A1(new_n710_), .A2(new_n715_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n713_), .A2(new_n716_), .ZN(G1337gat));
  OAI21_X1  g516(.A(G99gat), .B1(new_n710_), .B2(new_n249_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n250_), .A2(new_n495_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n706_), .A2(KEYINPUT112), .A3(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT112), .B1(new_n706_), .B2(new_n720_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n718_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT51), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT51), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n725_), .B(new_n718_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1338gat));
  NAND3_X1  g526(.A1(new_n706_), .A2(new_n421_), .A3(new_n496_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n708_), .A2(new_n421_), .A3(new_n709_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT52), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n729_), .A2(new_n730_), .A3(G106gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n729_), .B2(G106gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g533(.A1(new_n444_), .A2(new_n250_), .A3(new_n385_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n478_), .B1(new_n563_), .B2(new_n568_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n549_), .A2(new_n557_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n559_), .A2(new_n515_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n561_), .A2(new_n737_), .A3(KEYINPUT55), .A4(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(KEYINPUT114), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT114), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n560_), .A2(new_n741_), .A3(KEYINPUT55), .A4(new_n561_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT55), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n547_), .B1(new_n551_), .B2(new_n507_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n738_), .B1(new_n744_), .B2(KEYINPUT12), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n552_), .A2(new_n554_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n743_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n552_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n555_), .B1(new_n745_), .B2(new_n748_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n740_), .A2(new_n742_), .A3(new_n747_), .A4(new_n749_), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n750_), .A2(KEYINPUT115), .A3(KEYINPUT56), .A4(new_n567_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(KEYINPUT56), .A3(new_n567_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT115), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(KEYINPUT56), .B1(new_n750_), .B2(new_n567_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n736_), .B(new_n751_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n569_), .A2(new_n571_), .ZN(new_n757_));
  AOI22_X1  g556(.A1(new_n463_), .A2(new_n465_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n475_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n464_), .B1(new_n458_), .B2(new_n462_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n469_), .ZN(new_n761_));
  AOI22_X1  g560(.A1(new_n758_), .A2(new_n475_), .B1(new_n759_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n757_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n756_), .A2(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(KEYINPUT57), .B1(new_n764_), .B2(new_n602_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT57), .ZN(new_n766_));
  AOI211_X1 g565(.A(new_n766_), .B(new_n537_), .C1(new_n756_), .C2(new_n763_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n765_), .A2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n750_), .A2(new_n567_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT56), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT116), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n772_), .A3(new_n752_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n569_), .A2(new_n762_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n774_), .B1(new_n755_), .B2(KEYINPUT116), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT58), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT117), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n778_), .A2(new_n779_), .A3(new_n539_), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT58), .B1(new_n773_), .B2(new_n775_), .ZN(new_n781_));
  OAI21_X1  g580(.A(KEYINPUT117), .B1(new_n781_), .B2(new_n639_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n773_), .A2(new_n775_), .A3(KEYINPUT58), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n780_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n768_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n588_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n589_), .A2(KEYINPUT113), .A3(new_n787_), .A4(new_n478_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT113), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n639_), .A2(new_n478_), .A3(new_n574_), .A4(new_n587_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n789_), .B1(new_n790_), .B2(KEYINPUT54), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(KEYINPUT54), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n788_), .A2(new_n791_), .A3(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n735_), .B1(new_n786_), .B2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(G113gat), .B1(new_n794_), .B2(new_n594_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n587_), .B1(new_n768_), .B2(new_n784_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT119), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  AOI211_X1 g597(.A(KEYINPUT119), .B(new_n587_), .C1(new_n768_), .C2(new_n784_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n793_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n735_), .A2(KEYINPUT59), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n735_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n788_), .A2(new_n791_), .A3(new_n792_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n803_), .B1(new_n804_), .B2(new_n796_), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n805_), .A2(KEYINPUT118), .A3(KEYINPUT59), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT118), .B1(new_n805_), .B2(KEYINPUT59), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n802_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n594_), .A2(G113gat), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(KEYINPUT120), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n795_), .B1(new_n809_), .B2(new_n811_), .ZN(G1340gat));
  OAI21_X1  g611(.A(G120gat), .B1(new_n808_), .B2(new_n574_), .ZN(new_n813_));
  INV_X1    g612(.A(G120gat), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n574_), .B2(KEYINPUT60), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n794_), .B(new_n815_), .C1(KEYINPUT60), .C2(new_n814_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n813_), .A2(new_n816_), .ZN(G1341gat));
  OAI21_X1  g616(.A(G127gat), .B1(new_n808_), .B2(new_n588_), .ZN(new_n818_));
  OR3_X1    g617(.A1(new_n805_), .A2(G127gat), .A3(new_n588_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(G1342gat));
  INV_X1    g619(.A(G134gat), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n821_), .B1(new_n805_), .B2(new_n603_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT121), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n822_), .B(new_n823_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n639_), .A2(new_n821_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n824_), .B1(new_n809_), .B2(new_n825_), .ZN(G1343gat));
  NAND2_X1  g625(.A1(new_n786_), .A2(new_n793_), .ZN(new_n827_));
  NOR4_X1   g626(.A1(new_n250_), .A2(new_n610_), .A3(new_n422_), .A4(new_n419_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n594_), .ZN(new_n831_));
  XNOR2_X1  g630(.A(KEYINPUT122), .B(G141gat), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n831_), .B(new_n832_), .ZN(G1344gat));
  NAND2_X1  g632(.A1(new_n830_), .A2(new_n575_), .ZN(new_n834_));
  XOR2_X1   g633(.A(KEYINPUT123), .B(G148gat), .Z(new_n835_));
  XNOR2_X1  g634(.A(new_n834_), .B(new_n835_), .ZN(G1345gat));
  OR3_X1    g635(.A1(new_n829_), .A2(KEYINPUT124), .A3(new_n588_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT124), .B1(new_n829_), .B2(new_n588_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(KEYINPUT61), .B(G155gat), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n837_), .A2(new_n838_), .A3(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n839_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n840_), .A2(new_n841_), .ZN(G1346gat));
  OAI211_X1 g641(.A(new_n604_), .B(new_n828_), .C1(new_n804_), .C2(new_n796_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT125), .ZN(new_n844_));
  INV_X1    g643(.A(G162gat), .ZN(new_n845_));
  AND3_X1   g644(.A1(new_n843_), .A2(new_n844_), .A3(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n844_), .B1(new_n843_), .B2(new_n845_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n539_), .A2(G162gat), .ZN(new_n848_));
  OAI22_X1  g647(.A1(new_n846_), .A2(new_n847_), .B1(new_n829_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT126), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  OAI221_X1 g650(.A(KEYINPUT126), .B1(new_n829_), .B2(new_n848_), .C1(new_n846_), .C2(new_n847_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1347gat));
  INV_X1    g652(.A(KEYINPUT22), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n432_), .A2(new_n429_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n856_), .A2(new_n421_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n800_), .A2(new_n854_), .A3(new_n594_), .A4(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(G169gat), .ZN(new_n859_));
  AND3_X1   g658(.A1(new_n858_), .A2(KEYINPUT62), .A3(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(KEYINPUT62), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT62), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n800_), .A2(new_n862_), .A3(new_n594_), .A4(new_n857_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n863_), .A2(G169gat), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n860_), .B1(new_n861_), .B2(new_n864_), .ZN(G1348gat));
  NAND3_X1  g664(.A1(new_n800_), .A2(new_n575_), .A3(new_n857_), .ZN(new_n866_));
  INV_X1    g665(.A(G176gat), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT127), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n866_), .A2(KEYINPUT127), .A3(new_n867_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n421_), .B1(new_n786_), .B2(new_n793_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n574_), .A2(new_n856_), .A3(new_n867_), .ZN(new_n873_));
  AOI22_X1  g672(.A1(new_n870_), .A2(new_n871_), .B1(new_n872_), .B2(new_n873_), .ZN(G1349gat));
  NOR2_X1   g673(.A1(new_n856_), .A2(new_n588_), .ZN(new_n875_));
  AOI21_X1  g674(.A(G183gat), .B1(new_n872_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n800_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n857_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n305_), .A2(new_n306_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n587_), .A2(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n876_), .B1(new_n879_), .B2(new_n881_), .ZN(G1350gat));
  NAND3_X1  g681(.A1(new_n879_), .A2(new_n222_), .A3(new_n604_), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n877_), .A2(new_n639_), .A3(new_n878_), .ZN(new_n884_));
  INV_X1    g683(.A(G190gat), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n883_), .B1(new_n884_), .B2(new_n885_), .ZN(G1351gat));
  AND4_X1   g685(.A1(new_n249_), .A2(new_n827_), .A3(new_n424_), .A4(new_n610_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n594_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n575_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g690(.A(KEYINPUT63), .B(G211gat), .C1(new_n887_), .C2(new_n587_), .ZN(new_n892_));
  XOR2_X1   g691(.A(KEYINPUT63), .B(G211gat), .Z(new_n893_));
  AND3_X1   g692(.A1(new_n887_), .A2(new_n587_), .A3(new_n893_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n892_), .A2(new_n894_), .ZN(G1354gat));
  NAND3_X1  g694(.A1(new_n887_), .A2(new_n316_), .A3(new_n604_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n887_), .A2(new_n539_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n896_), .B1(new_n898_), .B2(new_n316_), .ZN(G1355gat));
endmodule


