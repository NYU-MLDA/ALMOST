//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 1 1 1 1 0 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 1 1 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n741_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n822_, new_n823_, new_n825_, new_n826_,
    new_n827_, new_n829_, new_n830_, new_n831_, new_n832_, new_n834_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n859_, new_n860_, new_n862_, new_n863_, new_n864_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_;
  INV_X1    g000(.A(KEYINPUT64), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G99gat), .A2(G106gat), .ZN(new_n203_));
  AOI21_X1  g002(.A(new_n202_), .B1(new_n203_), .B2(KEYINPUT65), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT7), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT6), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT7), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n208_), .B1(new_n203_), .B2(new_n202_), .ZN(new_n209_));
  OAI211_X1 g008(.A(new_n205_), .B(new_n207_), .C1(new_n204_), .C2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT66), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT8), .ZN(new_n212_));
  XOR2_X1   g011(.A(G85gat), .B(G92gat), .Z(new_n213_));
  NAND3_X1  g012(.A1(new_n210_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n211_), .A2(KEYINPUT8), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n214_), .A2(new_n215_), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT69), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n214_), .A2(new_n215_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT69), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(new_n221_), .A3(new_n216_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n213_), .A2(KEYINPUT9), .ZN(new_n223_));
  XOR2_X1   g022(.A(KEYINPUT10), .B(G99gat), .Z(new_n224_));
  INV_X1    g023(.A(G106gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT9), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(G85gat), .A3(G92gat), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n223_), .A2(new_n226_), .A3(new_n207_), .A4(new_n228_), .ZN(new_n229_));
  XOR2_X1   g028(.A(new_n229_), .B(KEYINPUT70), .Z(new_n230_));
  NAND3_X1  g029(.A1(new_n219_), .A2(new_n222_), .A3(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G29gat), .B(G36gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(G50gat), .ZN(new_n233_));
  XOR2_X1   g032(.A(KEYINPUT73), .B(G43gat), .Z(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT15), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n231_), .A2(new_n236_), .ZN(new_n237_));
  AND3_X1   g036(.A1(new_n220_), .A2(new_n216_), .A3(new_n229_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(new_n235_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G232gat), .A2(G233gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT34), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n237_), .B(new_n239_), .C1(KEYINPUT35), .C2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(KEYINPUT35), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n243_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G190gat), .B(G218gat), .ZN(new_n247_));
  INV_X1    g046(.A(G162gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT74), .B(G134gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n246_), .B1(KEYINPUT36), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT37), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n251_), .B(KEYINPUT36), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n244_), .A2(new_n254_), .A3(new_n245_), .ZN(new_n255_));
  AND3_X1   g054(.A1(new_n252_), .A2(new_n253_), .A3(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n253_), .B1(new_n252_), .B2(new_n255_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G231gat), .A2(G233gat), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G183gat), .B(G211gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G127gat), .B(G155gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT17), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT77), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G15gat), .B(G22gat), .ZN(new_n269_));
  INV_X1    g068(.A(G1gat), .ZN(new_n270_));
  INV_X1    g069(.A(G8gat), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT14), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n269_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G1gat), .B(G8gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n273_), .B(new_n274_), .Z(new_n275_));
  XNOR2_X1  g074(.A(new_n268_), .B(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT75), .ZN(new_n277_));
  INV_X1    g076(.A(new_n275_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n268_), .B(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT75), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n260_), .B1(new_n277_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT67), .B(G71gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(G78gat), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n285_), .A2(KEYINPUT11), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G57gat), .B(G64gat), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n285_), .A2(KEYINPUT11), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n287_), .B1(new_n286_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n277_), .A2(new_n281_), .A3(new_n260_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n283_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n288_), .A2(new_n290_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n292_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n294_), .B1(new_n295_), .B2(new_n282_), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n265_), .A2(KEYINPUT17), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n293_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT78), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n293_), .A2(new_n296_), .A3(KEYINPUT78), .A4(new_n297_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n258_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT79), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n231_), .A2(KEYINPUT12), .A3(new_n291_), .ZN(new_n305_));
  AND2_X1   g104(.A1(G230gat), .A2(G233gat), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n306_), .B1(new_n238_), .B2(new_n294_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n220_), .A2(new_n216_), .A3(new_n229_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(new_n291_), .ZN(new_n309_));
  XOR2_X1   g108(.A(KEYINPUT71), .B(KEYINPUT12), .Z(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n305_), .A2(new_n307_), .A3(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G230gat), .A2(G233gat), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT68), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n238_), .A2(new_n294_), .A3(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT68), .B1(new_n308_), .B2(new_n291_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n314_), .B1(new_n318_), .B2(new_n309_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G176gat), .B(G204gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G120gat), .B(G148gat), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n322_), .B(new_n323_), .Z(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  OR3_X1    g124(.A1(new_n313_), .A2(new_n319_), .A3(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n325_), .B1(new_n313_), .B2(new_n319_), .ZN(new_n327_));
  AND3_X1   g126(.A1(new_n326_), .A2(KEYINPUT13), .A3(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(KEYINPUT13), .B1(new_n326_), .B2(new_n327_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G169gat), .B(G197gat), .ZN(new_n331_));
  INV_X1    g130(.A(G141gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT81), .B(G113gat), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n333_), .B(new_n334_), .Z(new_n335_));
  XNOR2_X1  g134(.A(new_n235_), .B(KEYINPUT80), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n275_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n236_), .A2(new_n278_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G229gat), .A2(G233gat), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT80), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n235_), .B(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n278_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n339_), .B1(new_n337_), .B2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n335_), .B1(new_n340_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n337_), .A2(new_n343_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n339_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n335_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n348_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n345_), .A2(new_n351_), .A3(KEYINPUT82), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT82), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n353_), .B(new_n335_), .C1(new_n340_), .C2(new_n344_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n330_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT3), .ZN(new_n361_));
  INV_X1    g160(.A(G148gat), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n361_), .A2(new_n332_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G141gat), .A2(G148gat), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT2), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n363_), .A2(new_n366_), .A3(new_n367_), .A4(new_n368_), .ZN(new_n369_));
  AND2_X1   g168(.A1(G155gat), .A2(G162gat), .ZN(new_n370_));
  NOR2_X1   g169(.A1(G155gat), .A2(G162gat), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n369_), .A2(new_n372_), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n370_), .A2(KEYINPUT1), .B1(new_n332_), .B2(new_n362_), .ZN(new_n374_));
  OR2_X1    g173(.A1(G155gat), .A2(G162gat), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT1), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G155gat), .A2(G162gat), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n374_), .A2(new_n378_), .A3(new_n364_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT29), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n373_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT93), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT93), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n373_), .A2(new_n379_), .A3(new_n383_), .A4(new_n380_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G22gat), .B(G50gat), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n382_), .A2(new_n384_), .A3(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n386_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n360_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n382_), .A2(new_n384_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n385_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n382_), .A2(new_n384_), .A3(new_n386_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(new_n359_), .A3(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n389_), .A2(new_n393_), .A3(KEYINPUT95), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G78gat), .B(G106gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G211gat), .B(G218gat), .ZN(new_n397_));
  INV_X1    g196(.A(G197gat), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n398_), .A2(G204gat), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n397_), .B(KEYINPUT21), .C1(KEYINPUT94), .C2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G197gat), .B(G204gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n397_), .A2(KEYINPUT21), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n399_), .A2(KEYINPUT94), .ZN(new_n404_));
  INV_X1    g203(.A(new_n401_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n404_), .A2(new_n405_), .A3(KEYINPUT21), .A4(new_n397_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n402_), .A2(new_n403_), .A3(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n373_), .A2(new_n379_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n407_), .B1(KEYINPUT29), .B2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G228gat), .A2(G233gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n395_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n389_), .A2(new_n393_), .A3(new_n412_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n396_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n411_), .B1(new_n396_), .B2(new_n413_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G113gat), .B(G120gat), .ZN(new_n418_));
  INV_X1    g217(.A(G134gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(G127gat), .ZN(new_n420_));
  INV_X1    g219(.A(G127gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(G134gat), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT90), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n420_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n423_), .B1(new_n420_), .B2(new_n422_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n418_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n421_), .A2(G134gat), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n419_), .A2(G127gat), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT90), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n418_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n420_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n429_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n426_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n364_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n434_), .B1(new_n372_), .B2(new_n376_), .ZN(new_n435_));
  AOI22_X1  g234(.A1(new_n435_), .A2(new_n374_), .B1(new_n369_), .B2(new_n372_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n433_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n408_), .A2(new_n432_), .A3(new_n426_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(KEYINPUT97), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT97), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n408_), .A2(new_n440_), .A3(new_n432_), .A4(new_n426_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n439_), .A2(KEYINPUT4), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT4), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n438_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G225gat), .A2(G233gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT98), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n445_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n439_), .A2(new_n441_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n446_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT100), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G57gat), .B(G85gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G1gat), .B(G29gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT100), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n450_), .A2(new_n458_), .A3(new_n446_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n449_), .A2(new_n452_), .A3(new_n457_), .A4(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT33), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n460_), .A2(KEYINPUT101), .A3(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n461_), .B1(new_n460_), .B2(KEYINPUT101), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G169gat), .A2(G176gat), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT85), .B1(G169gat), .B2(G176gat), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NOR3_X1   g265(.A1(KEYINPUT85), .A2(G169gat), .A3(G176gat), .ZN(new_n467_));
  OAI211_X1 g266(.A(KEYINPUT24), .B(new_n464_), .C1(new_n466_), .C2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT26), .B(G190gat), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT25), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(G183gat), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT84), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n470_), .A2(KEYINPUT84), .A3(G183gat), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n469_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(G183gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT25), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT83), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n476_), .A2(KEYINPUT83), .A3(KEYINPUT25), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n468_), .B1(new_n475_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT86), .ZN(new_n483_));
  INV_X1    g282(.A(G190gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT23), .B1(new_n476_), .B2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT23), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n486_), .A2(G183gat), .A3(G190gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n467_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(new_n465_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n488_), .B1(new_n490_), .B2(KEYINPUT24), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT87), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT87), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n493_), .B(new_n488_), .C1(new_n490_), .C2(KEYINPUT24), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT86), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n468_), .B(new_n495_), .C1(new_n475_), .C2(new_n481_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n483_), .A2(new_n492_), .A3(new_n494_), .A4(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n488_), .B1(G183gat), .B2(G190gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT22), .B(G169gat), .ZN(new_n499_));
  INV_X1    g298(.A(G176gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n498_), .A2(new_n501_), .A3(new_n464_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n407_), .B1(new_n497_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n407_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n471_), .A2(new_n477_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(new_n469_), .ZN(new_n507_));
  OR3_X1    g306(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n507_), .A2(new_n488_), .A3(new_n468_), .A4(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n502_), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT20), .B1(new_n504_), .B2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G226gat), .A2(G233gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  OR3_X1    g313(.A1(new_n503_), .A2(new_n511_), .A3(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G8gat), .B(G36gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(G92gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT18), .B(G64gat), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n517_), .B(new_n518_), .Z(new_n519_));
  NAND3_X1  g318(.A1(new_n497_), .A2(new_n502_), .A3(new_n407_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT20), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n521_), .B1(new_n504_), .B2(new_n510_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n514_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n515_), .A2(new_n519_), .A3(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n445_), .A2(new_n446_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n457_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n450_), .A2(new_n448_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n526_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n519_), .ZN(new_n530_));
  NOR3_X1   g329(.A1(new_n503_), .A2(new_n511_), .A3(new_n514_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n514_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n532_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n530_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n525_), .A2(new_n529_), .A3(new_n534_), .ZN(new_n535_));
  NOR3_X1   g334(.A1(new_n462_), .A2(new_n463_), .A3(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n519_), .A2(KEYINPUT32), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n514_), .B1(new_n503_), .B2(new_n511_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n520_), .A2(new_n532_), .A3(new_n522_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n537_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n515_), .A2(new_n524_), .A3(new_n537_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n452_), .A2(new_n459_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n447_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n527_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  AOI211_X1 g343(.A(new_n540_), .B(new_n541_), .C1(new_n544_), .C2(new_n460_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n417_), .B1(new_n536_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT102), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n525_), .A2(new_n534_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT27), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT104), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n548_), .A2(KEYINPUT104), .A3(new_n549_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n459_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n458_), .B1(new_n450_), .B2(new_n446_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n457_), .B1(new_n557_), .B2(new_n449_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n460_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n538_), .A2(new_n539_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(new_n530_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n562_), .A2(new_n525_), .A3(KEYINPUT27), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT103), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n562_), .A2(new_n525_), .A3(KEYINPUT103), .A4(KEYINPUT27), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n554_), .A2(new_n560_), .A3(new_n567_), .A4(new_n416_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n460_), .A2(KEYINPUT101), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT33), .ZN(new_n570_));
  AND3_X1   g369(.A1(new_n525_), .A2(new_n529_), .A3(new_n534_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n460_), .A2(KEYINPUT101), .A3(new_n461_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n570_), .A2(new_n571_), .A3(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n541_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n540_), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n574_), .B(new_n575_), .C1(new_n558_), .C2(new_n559_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT102), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n577_), .A2(new_n578_), .A3(new_n417_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n547_), .A2(new_n568_), .A3(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n433_), .B(KEYINPUT91), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT88), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n497_), .A2(new_n502_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n582_), .A2(new_n584_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT89), .B(KEYINPUT30), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n586_), .A2(new_n587_), .A3(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n589_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G15gat), .B(G43gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT31), .ZN(new_n593_));
  XOR2_X1   g392(.A(G71gat), .B(G99gat), .Z(new_n594_));
  XOR2_X1   g393(.A(new_n593_), .B(new_n594_), .Z(new_n595_));
  NAND2_X1  g394(.A1(G227gat), .A2(G233gat), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n595_), .B(new_n596_), .Z(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  OR3_X1    g397(.A1(new_n590_), .A2(new_n591_), .A3(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n598_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n580_), .A2(new_n601_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n554_), .A2(new_n417_), .A3(new_n560_), .A4(new_n567_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n603_), .A2(new_n601_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n602_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n304_), .A2(new_n358_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n560_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n608_), .A2(new_n270_), .A3(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT38), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n252_), .A2(new_n255_), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(KEYINPUT105), .Z(new_n613_));
  AND2_X1   g412(.A1(new_n606_), .A2(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n614_), .A2(new_n358_), .A3(new_n302_), .ZN(new_n615_));
  OAI21_X1  g414(.A(G1gat), .B1(new_n615_), .B2(new_n560_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n611_), .A2(new_n616_), .ZN(G1324gat));
  AND2_X1   g416(.A1(new_n554_), .A2(new_n567_), .ZN(new_n618_));
  OAI21_X1  g417(.A(G8gat), .B1(new_n615_), .B2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT39), .ZN(new_n620_));
  INV_X1    g419(.A(new_n618_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n608_), .A2(new_n271_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(G1325gat));
  OR3_X1    g424(.A1(new_n607_), .A2(G15gat), .A3(new_n601_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G15gat), .B1(new_n615_), .B2(new_n601_), .ZN(new_n627_));
  XOR2_X1   g426(.A(KEYINPUT107), .B(KEYINPUT41), .Z(new_n628_));
  AND2_X1   g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n627_), .A2(new_n628_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n626_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT108), .Z(G1326gat));
  OAI21_X1  g431(.A(G22gat), .B1(new_n615_), .B2(new_n417_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT42), .ZN(new_n634_));
  OR3_X1    g433(.A1(new_n607_), .A2(G22gat), .A3(new_n417_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT109), .ZN(G1327gat));
  NAND2_X1  g436(.A1(new_n606_), .A2(new_n612_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n357_), .A2(new_n302_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n638_), .A2(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(G29gat), .B1(new_n641_), .B2(new_n609_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT113), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n643_), .B1(KEYINPUT112), .B2(KEYINPUT44), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n644_), .B1(new_n643_), .B2(KEYINPUT44), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT43), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT110), .B1(new_n602_), .B2(new_n605_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT110), .ZN(new_n648_));
  AOI211_X1 g447(.A(new_n648_), .B(new_n604_), .C1(new_n580_), .C2(new_n601_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n647_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT111), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n256_), .A2(new_n257_), .A3(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n612_), .A2(KEYINPUT37), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n252_), .A2(new_n253_), .A3(new_n255_), .ZN(new_n654_));
  AOI21_X1  g453(.A(KEYINPUT111), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n652_), .A2(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n646_), .B1(new_n650_), .B2(new_n656_), .ZN(new_n657_));
  AOI211_X1 g456(.A(KEYINPUT43), .B(new_n258_), .C1(new_n602_), .C2(new_n605_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n639_), .B(new_n645_), .C1(new_n657_), .C2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n601_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n578_), .B1(new_n577_), .B2(new_n417_), .ZN(new_n661_));
  AOI211_X1 g460(.A(KEYINPUT102), .B(new_n416_), .C1(new_n573_), .C2(new_n576_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n660_), .B1(new_n663_), .B2(new_n568_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n648_), .B1(new_n664_), .B2(new_n604_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n602_), .A2(KEYINPUT110), .A3(new_n605_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n665_), .A2(new_n656_), .A3(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n658_), .B1(new_n667_), .B2(KEYINPUT43), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n644_), .B1(new_n668_), .B2(new_n640_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n659_), .A2(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n609_), .A2(G29gat), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n642_), .B1(new_n670_), .B2(new_n671_), .ZN(G1328gat));
  NAND3_X1  g471(.A1(new_n659_), .A2(new_n669_), .A3(new_n621_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(G36gat), .ZN(new_n674_));
  INV_X1    g473(.A(G36gat), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n641_), .A2(new_n675_), .A3(new_n621_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT45), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n676_), .B(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n674_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT114), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT46), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n678_), .B1(new_n673_), .B2(G36gat), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT46), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n683_), .A2(KEYINPUT114), .A3(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n682_), .A2(new_n685_), .ZN(G1329gat));
  NAND3_X1  g485(.A1(new_n670_), .A2(G43gat), .A3(new_n660_), .ZN(new_n687_));
  AOI21_X1  g486(.A(G43gat), .B1(new_n641_), .B2(new_n660_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT115), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT47), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT47), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n687_), .A2(new_n692_), .A3(new_n689_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1330gat));
  INV_X1    g493(.A(G50gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n641_), .A2(new_n695_), .A3(new_n416_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n670_), .A2(new_n416_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n696_), .B1(new_n697_), .B2(new_n695_), .ZN(G1331gat));
  NOR2_X1   g497(.A1(new_n330_), .A2(new_n356_), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n304_), .A2(new_n606_), .A3(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(G57gat), .B1(new_n700_), .B2(new_n609_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n614_), .A2(new_n699_), .A3(new_n302_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT116), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT116), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n614_), .A2(new_n699_), .A3(new_n704_), .A4(new_n302_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n609_), .A2(G57gat), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n701_), .B1(new_n706_), .B2(new_n707_), .ZN(G1332gat));
  INV_X1    g507(.A(G64gat), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n700_), .A2(new_n709_), .A3(new_n621_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n703_), .A2(new_n621_), .A3(new_n705_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT48), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n711_), .A2(new_n712_), .A3(G64gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n711_), .B2(G64gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n710_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT117), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n715_), .B(new_n716_), .ZN(G1333gat));
  INV_X1    g516(.A(G71gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n700_), .A2(new_n718_), .A3(new_n660_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT49), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n706_), .A2(new_n660_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n721_), .B2(G71gat), .ZN(new_n722_));
  AOI211_X1 g521(.A(KEYINPUT49), .B(new_n718_), .C1(new_n706_), .C2(new_n660_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n719_), .B1(new_n722_), .B2(new_n723_), .ZN(G1334gat));
  INV_X1    g523(.A(G78gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n700_), .A2(new_n725_), .A3(new_n416_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n706_), .A2(new_n416_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(G78gat), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n728_), .A2(KEYINPUT50), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n728_), .A2(KEYINPUT50), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n726_), .B1(new_n729_), .B2(new_n730_), .ZN(G1335gat));
  INV_X1    g530(.A(new_n302_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n699_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n638_), .A2(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(G85gat), .B1(new_n734_), .B2(new_n609_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n668_), .A2(new_n733_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n609_), .A2(G85gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n735_), .B1(new_n736_), .B2(new_n737_), .ZN(G1336gat));
  AOI21_X1  g537(.A(G92gat), .B1(new_n734_), .B2(new_n621_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n621_), .A2(G92gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n736_), .B2(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT118), .ZN(G1337gat));
  NAND3_X1  g541(.A1(new_n734_), .A2(new_n224_), .A3(new_n660_), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n668_), .A2(new_n601_), .A3(new_n733_), .ZN(new_n744_));
  INV_X1    g543(.A(G99gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n743_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g546(.A1(new_n734_), .A2(new_n225_), .A3(new_n416_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n736_), .A2(new_n416_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(new_n751_), .A3(G106gat), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n668_), .A2(new_n417_), .A3(new_n733_), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT52), .B1(new_n753_), .B2(new_n225_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n749_), .B1(new_n752_), .B2(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n755_), .B(new_n757_), .ZN(G1339gat));
  NAND3_X1  g557(.A1(new_n318_), .A2(new_n305_), .A3(new_n311_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(new_n306_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT55), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n312_), .A2(new_n761_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n305_), .A2(new_n307_), .A3(KEYINPUT55), .A4(new_n311_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n760_), .A2(new_n762_), .A3(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n325_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT56), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT56), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n764_), .A2(new_n767_), .A3(new_n325_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n766_), .A2(new_n356_), .A3(new_n326_), .A4(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n337_), .A2(new_n338_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT120), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n337_), .A2(new_n338_), .A3(KEYINPUT120), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n772_), .A2(new_n347_), .A3(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n350_), .B1(new_n346_), .B2(new_n339_), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n774_), .A2(KEYINPUT121), .A3(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT121), .B1(new_n774_), .B2(new_n775_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n351_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n776_), .A2(new_n777_), .A3(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n326_), .A2(new_n327_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n612_), .B1(new_n769_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT57), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n782_), .B(new_n783_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n779_), .A2(new_n766_), .A3(new_n326_), .A4(new_n768_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT122), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT58), .ZN(new_n787_));
  INV_X1    g586(.A(new_n258_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT58), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n785_), .A2(KEYINPUT122), .A3(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n787_), .A2(new_n788_), .A3(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n302_), .B1(new_n784_), .B2(new_n791_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n258_), .A2(new_n302_), .A3(new_n330_), .A4(new_n355_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n793_), .B(new_n794_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n792_), .A2(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n621_), .A2(new_n560_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  NOR4_X1   g597(.A1(new_n796_), .A2(new_n601_), .A3(new_n416_), .A4(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(G113gat), .B1(new_n799_), .B2(new_n356_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(KEYINPUT123), .A3(KEYINPUT59), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n787_), .A2(new_n788_), .A3(new_n790_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n782_), .B(KEYINPUT57), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n732_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n793_), .B(KEYINPUT54), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n416_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n806_), .A2(KEYINPUT123), .A3(new_n660_), .A4(new_n797_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT59), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n355_), .B1(new_n801_), .B2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n800_), .B1(new_n810_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g610(.A(new_n330_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT60), .ZN(new_n813_));
  AOI21_X1  g612(.A(G120gat), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT124), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT124), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n816_), .B1(new_n813_), .B2(G120gat), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n799_), .B(new_n815_), .C1(new_n814_), .C2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n330_), .B1(new_n801_), .B2(new_n809_), .ZN(new_n819_));
  INV_X1    g618(.A(G120gat), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n818_), .B1(new_n819_), .B2(new_n820_), .ZN(G1341gat));
  AOI21_X1  g620(.A(G127gat), .B1(new_n799_), .B2(new_n302_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n732_), .B1(new_n801_), .B2(new_n809_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n823_), .B2(G127gat), .ZN(G1342gat));
  INV_X1    g623(.A(new_n613_), .ZN(new_n825_));
  AOI21_X1  g624(.A(G134gat), .B1(new_n799_), .B2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n258_), .B1(new_n801_), .B2(new_n809_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n826_), .B1(new_n827_), .B2(G134gat), .ZN(G1343gat));
  NOR2_X1   g627(.A1(new_n796_), .A2(new_n798_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n660_), .A2(new_n417_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n831_), .A2(new_n355_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(new_n332_), .ZN(G1344gat));
  NOR2_X1   g632(.A1(new_n831_), .A2(new_n330_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n834_), .B(new_n362_), .ZN(G1345gat));
  NOR2_X1   g634(.A1(new_n831_), .A2(new_n732_), .ZN(new_n836_));
  XOR2_X1   g635(.A(KEYINPUT61), .B(G155gat), .Z(new_n837_));
  XNOR2_X1  g636(.A(new_n836_), .B(new_n837_), .ZN(G1346gat));
  INV_X1    g637(.A(new_n831_), .ZN(new_n839_));
  AOI21_X1  g638(.A(G162gat), .B1(new_n839_), .B2(new_n825_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n652_), .A2(new_n655_), .A3(new_n248_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n840_), .B1(new_n839_), .B2(new_n841_), .ZN(G1347gat));
  INV_X1    g641(.A(KEYINPUT125), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n618_), .A2(new_n601_), .A3(new_n609_), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n417_), .B(new_n844_), .C1(new_n792_), .C2(new_n795_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n843_), .B1(new_n845_), .B2(new_n355_), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n806_), .A2(KEYINPUT125), .A3(new_n356_), .A4(new_n844_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(new_n847_), .A3(G169gat), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT126), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n846_), .A2(new_n847_), .A3(KEYINPUT126), .A4(G169gat), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n850_), .A2(KEYINPUT62), .A3(new_n851_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n806_), .A2(new_n356_), .A3(new_n499_), .A4(new_n844_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT62), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n848_), .A2(new_n849_), .A3(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n852_), .A2(new_n853_), .A3(new_n855_), .ZN(G1348gat));
  NOR2_X1   g655(.A1(new_n845_), .A2(new_n330_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(new_n500_), .ZN(G1349gat));
  NOR2_X1   g657(.A1(new_n845_), .A2(new_n732_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(G183gat), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n860_), .B1(new_n505_), .B2(new_n859_), .ZN(G1350gat));
  OAI21_X1  g660(.A(G190gat), .B1(new_n845_), .B2(new_n258_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n825_), .A2(new_n469_), .ZN(new_n863_));
  XOR2_X1   g662(.A(new_n863_), .B(KEYINPUT127), .Z(new_n864_));
  OAI21_X1  g663(.A(new_n862_), .B1(new_n845_), .B2(new_n864_), .ZN(G1351gat));
  NOR2_X1   g664(.A1(new_n796_), .A2(new_n609_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n660_), .A2(new_n618_), .A3(new_n417_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n355_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(new_n398_), .ZN(G1352gat));
  INV_X1    g669(.A(new_n868_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n812_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g672(.A1(new_n868_), .A2(new_n732_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n875_));
  AND2_X1   g674(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n874_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n877_), .B1(new_n874_), .B2(new_n875_), .ZN(G1354gat));
  AND3_X1   g677(.A1(new_n871_), .A2(G218gat), .A3(new_n788_), .ZN(new_n879_));
  AOI21_X1  g678(.A(G218gat), .B1(new_n871_), .B2(new_n825_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1355gat));
endmodule


