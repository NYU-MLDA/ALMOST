//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 1 0 0 0 0 0 0 0 0 0 0 1 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_;
  INV_X1    g000(.A(G169gat), .ZN(new_n202_));
  INV_X1    g001(.A(G176gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n204_), .A2(KEYINPUT24), .A3(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT25), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT81), .B1(new_n207_), .B2(G183gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT81), .ZN(new_n209_));
  INV_X1    g008(.A(G183gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(new_n210_), .A3(KEYINPUT25), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n208_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n207_), .A2(G183gat), .ZN(new_n213_));
  INV_X1    g012(.A(G190gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT26), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT26), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(G190gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n213_), .A2(new_n215_), .A3(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n206_), .B1(new_n212_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT82), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  OR2_X1    g020(.A1(new_n204_), .A2(KEYINPUT24), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n223_));
  AND2_X1   g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT84), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT23), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT83), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT83), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT23), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n227_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT84), .ZN(new_n231_));
  INV_X1    g030(.A(new_n224_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n224_), .A2(new_n226_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n225_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  OAI211_X1 g034(.A(KEYINPUT82), .B(new_n206_), .C1(new_n212_), .C2(new_n218_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n221_), .A2(new_n222_), .A3(new_n235_), .A4(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n224_), .A2(KEYINPUT23), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n238_), .B1(new_n224_), .B2(new_n230_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(G183gat), .A2(G190gat), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n202_), .A2(KEYINPUT22), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT22), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(G169gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(new_n245_), .A3(new_n203_), .ZN(new_n246_));
  AOI22_X1  g045(.A1(new_n246_), .A2(KEYINPUT85), .B1(G169gat), .B2(G176gat), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n242_), .B(new_n247_), .C1(KEYINPUT85), .C2(new_n246_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n237_), .A2(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(KEYINPUT86), .B(G43gat), .Z(new_n250_));
  XNOR2_X1  g049(.A(G71gat), .B(G99gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n249_), .A2(new_n252_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n249_), .A2(new_n252_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(G134gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(G127gat), .ZN(new_n257_));
  INV_X1    g056(.A(G127gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(G134gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT87), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n257_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n260_), .B1(new_n257_), .B2(new_n259_), .ZN(new_n263_));
  INV_X1    g062(.A(G120gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(G113gat), .ZN(new_n265_));
  INV_X1    g064(.A(G113gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(G120gat), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n265_), .A2(new_n267_), .A3(KEYINPUT88), .ZN(new_n268_));
  AOI21_X1  g067(.A(KEYINPUT88), .B1(new_n265_), .B2(new_n267_), .ZN(new_n269_));
  OAI22_X1  g068(.A1(new_n262_), .A2(new_n263_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n258_), .A2(G134gat), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n256_), .A2(G127gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT87), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT88), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n266_), .A2(G120gat), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n264_), .A2(G113gat), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n274_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n265_), .A2(new_n267_), .A3(KEYINPUT88), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n273_), .A2(new_n277_), .A3(new_n261_), .A4(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT89), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n270_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  AOI22_X1  g080(.A1(new_n261_), .A2(new_n273_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT89), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n255_), .A2(new_n284_), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n283_), .B(new_n281_), .C1(new_n254_), .C2(new_n253_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G227gat), .A2(G233gat), .ZN(new_n287_));
  INV_X1    g086(.A(G15gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT30), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT31), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n285_), .A2(new_n286_), .A3(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n291_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(G204gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G197gat), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n296_), .A2(KEYINPUT93), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(KEYINPUT93), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n295_), .A2(G197gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT94), .B(KEYINPUT21), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n297_), .A2(new_n298_), .A3(new_n299_), .A4(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(G211gat), .B(G218gat), .Z(new_n302_));
  NAND2_X1  g101(.A1(new_n299_), .A2(new_n296_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n302_), .B1(new_n303_), .B2(KEYINPUT21), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n302_), .A2(KEYINPUT21), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n297_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n301_), .A2(new_n304_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT3), .ZN(new_n308_));
  INV_X1    g107(.A(G141gat), .ZN(new_n309_));
  INV_X1    g108(.A(G148gat), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n308_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G141gat), .A2(G148gat), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT2), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n311_), .A2(new_n314_), .A3(new_n315_), .A4(new_n316_), .ZN(new_n317_));
  OR2_X1    g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G155gat), .A2(G162gat), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n317_), .A2(KEYINPUT91), .A3(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(KEYINPUT91), .B1(new_n317_), .B2(new_n320_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT90), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n323_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT90), .B1(G141gat), .B2(G148gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT1), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n318_), .A2(new_n327_), .A3(new_n319_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n329_), .A2(new_n312_), .ZN(new_n330_));
  AND3_X1   g129(.A1(new_n326_), .A2(new_n328_), .A3(new_n330_), .ZN(new_n331_));
  OR3_X1    g130(.A1(new_n321_), .A2(new_n322_), .A3(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n307_), .B1(new_n332_), .B2(KEYINPUT29), .ZN(new_n333_));
  XOR2_X1   g132(.A(G22gat), .B(G50gat), .Z(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  XOR2_X1   g135(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n337_));
  OR3_X1    g136(.A1(new_n332_), .A2(KEYINPUT29), .A3(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G228gat), .A2(G233gat), .ZN(new_n339_));
  INV_X1    g138(.A(G78gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(G106gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n337_), .B1(new_n332_), .B2(KEYINPUT29), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n338_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n344_), .B1(new_n338_), .B2(new_n345_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n336_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n348_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n350_), .A2(new_n335_), .A3(new_n346_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G1gat), .B(G29gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(G85gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT0), .B(G57gat), .ZN(new_n356_));
  XOR2_X1   g155(.A(new_n355_), .B(new_n356_), .Z(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT4), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n284_), .A2(new_n332_), .ZN(new_n360_));
  AND4_X1   g159(.A1(new_n261_), .A2(new_n273_), .A3(new_n277_), .A4(new_n278_), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT101), .B1(new_n361_), .B2(new_n282_), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n321_), .A2(new_n322_), .A3(new_n331_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT101), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n270_), .A2(new_n279_), .A3(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n362_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n360_), .A2(new_n366_), .A3(KEYINPUT102), .ZN(new_n367_));
  AND3_X1   g166(.A1(new_n270_), .A2(new_n364_), .A3(new_n279_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n364_), .B1(new_n270_), .B2(new_n279_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT102), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(new_n371_), .A3(new_n363_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n359_), .B1(new_n367_), .B2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G225gat), .A2(G233gat), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n360_), .A2(KEYINPUT4), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n373_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n367_), .A2(new_n372_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(new_n374_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n358_), .B1(new_n376_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n374_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n375_), .ZN(new_n382_));
  AND4_X1   g181(.A1(new_n371_), .A2(new_n362_), .A3(new_n363_), .A4(new_n365_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n371_), .B1(new_n370_), .B2(new_n363_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n383_), .B1(new_n384_), .B2(new_n360_), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n381_), .B(new_n382_), .C1(new_n385_), .C2(new_n359_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(new_n357_), .A3(new_n378_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT104), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n380_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  OAI211_X1 g188(.A(KEYINPUT104), .B(new_n358_), .C1(new_n376_), .C2(new_n379_), .ZN(new_n390_));
  AOI211_X1 g189(.A(new_n294_), .B(new_n353_), .C1(new_n389_), .C2(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(G8gat), .B(G36gat), .Z(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G64gat), .B(G92gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G226gat), .A2(G233gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT19), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n237_), .A2(new_n248_), .A3(new_n307_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT20), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT95), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n215_), .A2(new_n217_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT96), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT25), .B(G183gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n408_), .A2(new_n222_), .A3(new_n206_), .A4(new_n239_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT98), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n224_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n234_), .B1(new_n411_), .B2(new_n231_), .ZN(new_n412_));
  NOR3_X1   g211(.A1(new_n223_), .A2(KEYINPUT84), .A3(new_n224_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n410_), .B(new_n241_), .C1(new_n412_), .C2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT97), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n246_), .A2(new_n415_), .A3(new_n205_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n415_), .B1(new_n246_), .B2(new_n205_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n414_), .A2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n410_), .B1(new_n235_), .B2(new_n241_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n409_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n307_), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n402_), .A2(new_n403_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n401_), .A2(KEYINPUT95), .A3(KEYINPUT20), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n400_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n241_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT98), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n427_), .A2(new_n414_), .A3(new_n418_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n428_), .A2(new_n307_), .A3(new_n409_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n249_), .A2(new_n422_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n429_), .A2(new_n430_), .A3(KEYINPUT20), .A4(new_n400_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n397_), .B1(new_n425_), .B2(new_n432_), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n401_), .A2(KEYINPUT95), .A3(KEYINPUT20), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT95), .B1(new_n401_), .B2(KEYINPUT20), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n307_), .B1(new_n428_), .B2(new_n409_), .ZN(new_n436_));
  NOR3_X1   g235(.A1(new_n434_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n396_), .B(new_n431_), .C1(new_n437_), .C2(new_n400_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n433_), .A2(KEYINPUT100), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT27), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n425_), .A2(new_n432_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT100), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n441_), .A2(new_n442_), .A3(new_n396_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n439_), .A2(new_n440_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT105), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n423_), .A2(new_n400_), .A3(new_n424_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n429_), .A2(new_n430_), .A3(KEYINPUT20), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n399_), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  OAI211_X1 g248(.A(KEYINPUT27), .B(new_n438_), .C1(new_n449_), .C2(new_n396_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n444_), .A2(new_n445_), .A3(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n445_), .B1(new_n444_), .B2(new_n450_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n391_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT106), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT106), .ZN(new_n455_));
  OAI211_X1 g254(.A(new_n455_), .B(new_n391_), .C1(new_n451_), .C2(new_n452_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n396_), .A2(KEYINPUT32), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n457_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n458_), .B1(new_n441_), .B2(new_n457_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n389_), .A2(new_n390_), .A3(new_n459_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n439_), .A2(new_n443_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT33), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n387_), .A2(new_n462_), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n386_), .A2(KEYINPUT33), .A3(new_n357_), .A4(new_n378_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n374_), .B1(new_n367_), .B2(new_n372_), .ZN(new_n465_));
  OR3_X1    g264(.A1(new_n465_), .A2(KEYINPUT103), .A3(new_n357_), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT103), .B1(new_n465_), .B2(new_n357_), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n374_), .B(new_n382_), .C1(new_n385_), .C2(new_n359_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n463_), .A2(new_n464_), .A3(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n460_), .B1(new_n461_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n352_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n389_), .A2(new_n390_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n473_), .A2(new_n444_), .A3(new_n353_), .A4(new_n450_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  AOI22_X1  g274(.A1(new_n454_), .A2(new_n456_), .B1(new_n475_), .B2(new_n294_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n477_));
  INV_X1    g276(.A(G99gat), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n478_), .A2(new_n342_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n477_), .B(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(G85gat), .A2(G92gat), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT9), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G85gat), .A2(G92gat), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n484_), .A2(KEYINPUT64), .A3(new_n483_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT64), .B1(new_n484_), .B2(new_n483_), .ZN(new_n486_));
  OAI221_X1 g285(.A(new_n482_), .B1(new_n483_), .B2(new_n484_), .C1(new_n485_), .C2(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(KEYINPUT10), .B(G99gat), .Z(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n342_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n480_), .A2(new_n487_), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT8), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT66), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n480_), .A2(new_n492_), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n477_), .A2(new_n479_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n477_), .A2(new_n479_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n494_), .A2(KEYINPUT66), .A3(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(G99gat), .A2(G106gat), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT7), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT67), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n497_), .B(KEYINPUT7), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT67), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n493_), .A2(new_n496_), .A3(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n482_), .A2(new_n484_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n491_), .B1(new_n505_), .B2(new_n507_), .ZN(new_n508_));
  AOI211_X1 g307(.A(KEYINPUT8), .B(new_n506_), .C1(new_n480_), .C2(new_n502_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n490_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G29gat), .B(G36gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G43gat), .B(G50gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT15), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n510_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G232gat), .A2(G233gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT34), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT35), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n513_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n515_), .B(new_n520_), .C1(new_n521_), .C2(new_n510_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n518_), .A2(new_n519_), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n523_), .ZN(new_n525_));
  XOR2_X1   g324(.A(G190gat), .B(G218gat), .Z(new_n526_));
  XNOR2_X1  g325(.A(G134gat), .B(G162gat), .ZN(new_n527_));
  OR2_X1    g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n527_), .ZN(new_n529_));
  AOI21_X1  g328(.A(KEYINPUT36), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT71), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n524_), .A2(new_n525_), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n528_), .A2(KEYINPUT36), .A3(new_n529_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n534_), .A2(new_n530_), .ZN(new_n535_));
  XOR2_X1   g334(.A(new_n535_), .B(KEYINPUT72), .Z(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n537_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n533_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G120gat), .B(G148gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT5), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G176gat), .B(G204gat), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n541_), .B(new_n542_), .Z(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT68), .B(G71gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(new_n340_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G57gat), .B(G64gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT11), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n545_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n546_), .B(KEYINPUT11), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n549_), .B1(new_n550_), .B2(new_n545_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n510_), .A2(new_n552_), .ZN(new_n553_));
  OAI211_X1 g352(.A(new_n490_), .B(new_n551_), .C1(new_n508_), .C2(new_n509_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G230gat), .A2(G233gat), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT69), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n555_), .A2(KEYINPUT69), .A3(new_n557_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n553_), .A2(KEYINPUT12), .A3(new_n554_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT12), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n510_), .A2(new_n564_), .A3(new_n552_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n557_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n543_), .B1(new_n562_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n563_), .A2(new_n565_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(new_n556_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n543_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n569_), .A2(new_n560_), .A3(new_n561_), .A4(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n567_), .A2(KEYINPUT13), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(KEYINPUT13), .B1(new_n567_), .B2(new_n571_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n288_), .A2(G22gat), .ZN(new_n576_));
  INV_X1    g375(.A(G22gat), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(G15gat), .ZN(new_n578_));
  INV_X1    g377(.A(G1gat), .ZN(new_n579_));
  INV_X1    g378(.A(G8gat), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT14), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT75), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n576_), .B(new_n578_), .C1(new_n581_), .C2(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n583_), .B1(new_n582_), .B2(new_n581_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G1gat), .B(G8gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT78), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n584_), .B(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n587_), .B(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(new_n513_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n587_), .B(new_n588_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(new_n521_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(G229gat), .A3(G233gat), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n592_), .A2(new_n514_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G229gat), .A2(G233gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT79), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n591_), .A2(new_n596_), .A3(new_n598_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n595_), .A2(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(G113gat), .B(G141gat), .Z(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT80), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G169gat), .B(G197gat), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n602_), .B(new_n603_), .Z(new_n604_));
  OR2_X1    g403(.A1(new_n600_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n595_), .A2(new_n599_), .A3(new_n604_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n575_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(G231gat), .A2(G233gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n590_), .B(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(new_n551_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT17), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G127gat), .B(G155gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT16), .ZN(new_n614_));
  XOR2_X1   g413(.A(G183gat), .B(G211gat), .Z(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n611_), .B1(new_n612_), .B2(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n610_), .B(new_n552_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n616_), .B(new_n612_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n617_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NOR4_X1   g421(.A1(new_n476_), .A2(new_n539_), .A3(new_n608_), .A4(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n473_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(G1gat), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT38), .ZN(new_n627_));
  INV_X1    g426(.A(new_n607_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n476_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT70), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n630_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n574_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(KEYINPUT70), .A3(new_n572_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n524_), .A2(new_n525_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n536_), .B(KEYINPUT73), .Z(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(new_n532_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT37), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT37), .ZN(new_n641_));
  AOI21_X1  g440(.A(KEYINPUT74), .B1(new_n539_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT74), .ZN(new_n643_));
  NOR4_X1   g442(.A1(new_n533_), .A2(new_n538_), .A3(new_n643_), .A4(KEYINPUT37), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n640_), .B1(new_n642_), .B2(new_n644_), .ZN(new_n645_));
  AND4_X1   g444(.A1(new_n629_), .A2(new_n635_), .A3(new_n645_), .A4(new_n621_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n646_), .A2(new_n579_), .A3(new_n624_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(new_n627_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n648_), .A2(KEYINPUT107), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n648_), .A2(KEYINPUT107), .ZN(new_n650_));
  OAI221_X1 g449(.A(new_n626_), .B1(new_n627_), .B2(new_n647_), .C1(new_n649_), .C2(new_n650_), .ZN(G1324gat));
  NAND2_X1  g450(.A1(new_n444_), .A2(new_n450_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(KEYINPUT105), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n444_), .A2(new_n445_), .A3(new_n450_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n646_), .A2(new_n580_), .A3(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT39), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n623_), .A2(new_n656_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n659_), .B2(G8gat), .ZN(new_n660_));
  AOI211_X1 g459(.A(KEYINPUT39), .B(new_n580_), .C1(new_n623_), .C2(new_n656_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n657_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n662_), .B(new_n663_), .Z(G1325gat));
  INV_X1    g463(.A(new_n294_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n288_), .B1(new_n623_), .B2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT41), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n646_), .A2(new_n288_), .A3(new_n665_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1326gat));
  AOI21_X1  g468(.A(new_n577_), .B1(new_n623_), .B2(new_n353_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(KEYINPUT109), .B(KEYINPUT42), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n670_), .B(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n646_), .A2(new_n577_), .A3(new_n353_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1327gat));
  NAND2_X1  g473(.A1(new_n622_), .A2(new_n539_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n632_), .A2(new_n572_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n629_), .A2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(G29gat), .B1(new_n678_), .B2(new_n624_), .ZN(new_n679_));
  OAI21_X1  g478(.A(KEYINPUT43), .B1(new_n476_), .B2(new_n645_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n439_), .A2(new_n443_), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n681_), .A2(new_n463_), .A3(new_n464_), .A4(new_n469_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n353_), .B1(new_n682_), .B2(new_n460_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n474_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n294_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n455_), .B1(new_n655_), .B2(new_n391_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n456_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n685_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n689_));
  INV_X1    g488(.A(new_n645_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n688_), .A2(new_n689_), .A3(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n680_), .A2(new_n691_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n608_), .A2(new_n621_), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n692_), .A2(KEYINPUT44), .A3(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(KEYINPUT44), .B1(new_n692_), .B2(new_n693_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n624_), .A2(G29gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n679_), .B1(new_n696_), .B2(new_n697_), .ZN(G1328gat));
  INV_X1    g497(.A(KEYINPUT112), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT46), .ZN(new_n700_));
  INV_X1    g499(.A(G36gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n701_), .B1(new_n696_), .B2(new_n656_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n655_), .A2(G36gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n629_), .A2(new_n677_), .A3(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT111), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n629_), .A2(KEYINPUT111), .A3(new_n677_), .A4(new_n703_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  XOR2_X1   g507(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n706_), .A2(new_n709_), .A3(new_n707_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n699_), .B(new_n700_), .C1(new_n702_), .C2(new_n713_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n711_), .A2(new_n712_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n699_), .A2(new_n700_), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n694_), .A2(new_n695_), .A3(new_n655_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n715_), .B(new_n716_), .C1(new_n701_), .C2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n714_), .A2(new_n718_), .ZN(G1329gat));
  AOI21_X1  g518(.A(G43gat), .B1(new_n678_), .B2(new_n665_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n665_), .A2(G43gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n696_), .B2(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n722_), .B(new_n723_), .ZN(G1330gat));
  AOI21_X1  g523(.A(G50gat), .B1(new_n678_), .B2(new_n353_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n353_), .A2(G50gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n696_), .B2(new_n726_), .ZN(G1331gat));
  NAND2_X1  g526(.A1(new_n454_), .A2(new_n456_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n607_), .B1(new_n728_), .B2(new_n685_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n729_), .A2(new_n676_), .A3(new_n645_), .A4(new_n621_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(G57gat), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n731_), .A2(new_n732_), .A3(new_n624_), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n533_), .A2(new_n538_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n622_), .A2(new_n607_), .ZN(new_n735_));
  AND4_X1   g534(.A1(new_n688_), .A2(new_n634_), .A3(new_n734_), .A4(new_n735_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n736_), .A2(new_n624_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n733_), .B1(new_n732_), .B2(new_n737_), .ZN(G1332gat));
  INV_X1    g537(.A(G64gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n736_), .B2(new_n656_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(KEYINPUT114), .B(KEYINPUT48), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n740_), .B(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n731_), .A2(new_n739_), .A3(new_n656_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1333gat));
  INV_X1    g543(.A(G71gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n736_), .B2(new_n665_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT49), .Z(new_n747_));
  NAND3_X1  g546(.A1(new_n731_), .A2(new_n745_), .A3(new_n665_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1334gat));
  NAND3_X1  g548(.A1(new_n731_), .A2(new_n340_), .A3(new_n353_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n736_), .A2(new_n353_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n752_), .B2(G78gat), .ZN(new_n753_));
  AOI211_X1 g552(.A(KEYINPUT50), .B(new_n340_), .C1(new_n736_), .C2(new_n353_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n750_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT115), .Z(G1335gat));
  NAND3_X1  g555(.A1(new_n676_), .A2(new_n628_), .A3(new_n622_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n757_), .B1(new_n680_), .B2(new_n691_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(G85gat), .B1(new_n759_), .B2(new_n473_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT116), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n675_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n729_), .B2(new_n762_), .ZN(new_n763_));
  AND4_X1   g562(.A1(new_n761_), .A2(new_n688_), .A3(new_n628_), .A4(new_n762_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  OR2_X1    g564(.A1(new_n473_), .A2(G85gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n760_), .B1(new_n765_), .B2(new_n766_), .ZN(G1336gat));
  OAI21_X1  g566(.A(new_n656_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n768_));
  INV_X1    g567(.A(G92gat), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n656_), .A2(G92gat), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT117), .ZN(new_n771_));
  AOI22_X1  g570(.A1(new_n768_), .A2(new_n769_), .B1(new_n758_), .B2(new_n771_), .ZN(G1337gat));
  NAND2_X1  g571(.A1(new_n665_), .A2(new_n488_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n774_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n775_));
  AOI211_X1 g574(.A(new_n294_), .B(new_n757_), .C1(new_n680_), .C2(new_n691_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(new_n478_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n778_), .A2(KEYINPUT120), .A3(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT120), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n781_), .B1(new_n777_), .B2(KEYINPUT51), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT119), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n779_), .B1(new_n777_), .B2(KEYINPUT118), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT118), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n775_), .B(new_n786_), .C1(new_n776_), .C2(new_n478_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n784_), .B1(new_n785_), .B2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n478_), .B1(new_n758_), .B2(new_n665_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n688_), .A2(new_n628_), .A3(new_n762_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT116), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n729_), .A2(new_n761_), .A3(new_n762_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n773_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(KEYINPUT118), .B1(new_n789_), .B2(new_n793_), .ZN(new_n794_));
  AND4_X1   g593(.A1(new_n784_), .A2(new_n794_), .A3(KEYINPUT51), .A4(new_n787_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n783_), .B1(new_n788_), .B2(new_n795_), .ZN(G1338gat));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n758_), .A2(new_n353_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n797_), .B1(new_n798_), .B2(G106gat), .ZN(new_n799_));
  AOI211_X1 g598(.A(KEYINPUT52), .B(new_n342_), .C1(new_n758_), .C2(new_n353_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n353_), .A2(new_n342_), .ZN(new_n801_));
  OAI22_X1  g600(.A1(new_n799_), .A2(new_n800_), .B1(new_n765_), .B2(new_n801_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g602(.A1(new_n735_), .A2(new_n575_), .ZN(new_n804_));
  OAI21_X1  g603(.A(KEYINPUT121), .B1(new_n690_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT121), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n645_), .A2(new_n806_), .A3(new_n575_), .A4(new_n735_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n805_), .A2(KEYINPUT54), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n805_), .A2(new_n807_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n563_), .A2(new_n557_), .A3(new_n565_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n569_), .A2(KEYINPUT55), .A3(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n570_), .B1(new_n566_), .B2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT56), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT123), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n813_), .A2(KEYINPUT56), .A3(new_n815_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n818_), .A2(new_n819_), .A3(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n598_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n591_), .A2(new_n596_), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n604_), .B1(new_n594_), .B2(new_n598_), .ZN(new_n824_));
  AOI22_X1  g623(.A1(new_n600_), .A2(new_n604_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n816_), .A2(KEYINPUT123), .A3(new_n817_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n821_), .A2(new_n571_), .A3(new_n825_), .A4(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT58), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n645_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  OR2_X1    g628(.A1(new_n827_), .A2(new_n828_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT122), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n818_), .A2(new_n831_), .A3(new_n820_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n816_), .A2(KEYINPUT122), .A3(new_n817_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n832_), .A2(new_n607_), .A3(new_n571_), .A4(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n567_), .A2(new_n571_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n825_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n734_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT57), .ZN(new_n839_));
  AOI22_X1  g638(.A1(new_n829_), .A2(new_n830_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n837_), .A2(KEYINPUT57), .A3(new_n734_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n808_), .B(new_n811_), .C1(new_n842_), .C2(new_n621_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT124), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n656_), .A2(new_n294_), .A3(new_n473_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n843_), .A2(new_n844_), .A3(new_n352_), .A4(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n811_), .A2(new_n808_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n621_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n352_), .B(new_n845_), .C1(new_n847_), .C2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT124), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n846_), .A2(new_n850_), .A3(new_n266_), .A4(new_n607_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n843_), .A2(KEYINPUT59), .A3(new_n352_), .A4(new_n845_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n849_), .A2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n628_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n851_), .B1(new_n855_), .B2(new_n266_), .ZN(G1340gat));
  OR2_X1    g655(.A1(new_n264_), .A2(KEYINPUT60), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n264_), .B1(new_n575_), .B2(KEYINPUT60), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n846_), .A2(new_n850_), .A3(new_n857_), .A4(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n635_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n860_), .B2(new_n264_), .ZN(G1341gat));
  NAND4_X1  g660(.A1(new_n846_), .A2(new_n850_), .A3(new_n258_), .A4(new_n621_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n622_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n863_), .B2(new_n258_), .ZN(G1342gat));
  NAND4_X1  g663(.A1(new_n846_), .A2(new_n850_), .A3(new_n256_), .A4(new_n539_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n645_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(new_n256_), .ZN(G1343gat));
  NOR2_X1   g666(.A1(new_n665_), .A2(new_n352_), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n655_), .A2(new_n624_), .A3(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n843_), .A2(new_n607_), .A3(new_n869_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g670(.A1(new_n843_), .A2(new_n634_), .A3(new_n869_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g672(.A1(new_n843_), .A2(new_n621_), .A3(new_n869_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(KEYINPUT61), .B(G155gat), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1346gat));
  AND4_X1   g675(.A1(G162gat), .A2(new_n843_), .A3(new_n690_), .A4(new_n869_), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n539_), .B(new_n869_), .C1(new_n847_), .C2(new_n848_), .ZN(new_n878_));
  INV_X1    g677(.A(G162gat), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT125), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n878_), .A2(KEYINPUT125), .A3(new_n879_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n877_), .B1(new_n882_), .B2(new_n883_), .ZN(G1347gat));
  INV_X1    g683(.A(KEYINPUT62), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n624_), .A2(new_n294_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n656_), .A2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n352_), .B(new_n888_), .C1(new_n847_), .C2(new_n848_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n889_), .A2(new_n628_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n885_), .B1(new_n890_), .B2(new_n202_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n890_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n892_));
  OAI211_X1 g691(.A(KEYINPUT62), .B(G169gat), .C1(new_n889_), .C2(new_n628_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n891_), .A2(new_n892_), .A3(new_n893_), .ZN(G1348gat));
  NAND3_X1  g693(.A1(new_n843_), .A2(KEYINPUT126), .A3(new_n352_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT126), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n847_), .A2(new_n848_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n897_), .B2(new_n353_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n635_), .A2(new_n203_), .A3(new_n887_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n895_), .A2(new_n898_), .A3(new_n899_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n203_), .B1(new_n889_), .B2(new_n575_), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n900_), .A2(new_n901_), .ZN(G1349gat));
  NOR3_X1   g701(.A1(new_n889_), .A2(new_n407_), .A3(new_n622_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n895_), .A2(new_n898_), .A3(new_n621_), .A4(new_n888_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n903_), .B1(new_n904_), .B2(new_n210_), .ZN(G1350gat));
  OAI21_X1  g704(.A(G190gat), .B1(new_n889_), .B2(new_n645_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n539_), .A2(new_n406_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n889_), .B2(new_n907_), .ZN(G1351gat));
  NAND3_X1  g707(.A1(new_n656_), .A2(new_n473_), .A3(new_n868_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n897_), .A2(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n607_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G197gat), .ZN(G1352gat));
  NOR3_X1   g711(.A1(new_n897_), .A2(new_n635_), .A3(new_n909_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(KEYINPUT127), .B(G204gat), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n913_), .B(new_n914_), .ZN(G1353gat));
  NOR3_X1   g714(.A1(new_n897_), .A2(new_n622_), .A3(new_n909_), .ZN(new_n916_));
  OR2_X1    g715(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  XOR2_X1   g717(.A(KEYINPUT63), .B(G211gat), .Z(new_n919_));
  AOI21_X1  g718(.A(new_n918_), .B1(new_n916_), .B2(new_n919_), .ZN(G1354gat));
  INV_X1    g719(.A(G218gat), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n910_), .A2(new_n921_), .A3(new_n539_), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n897_), .A2(new_n645_), .A3(new_n909_), .ZN(new_n923_));
  OAI21_X1  g722(.A(new_n922_), .B1(new_n921_), .B2(new_n923_), .ZN(G1355gat));
endmodule


