//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 1 0 1 1 1 1 1 0 1 0 1 0 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0 1 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n606_, new_n607_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n791_, new_n792_, new_n793_, new_n794_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n823_, new_n824_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n845_, new_n846_, new_n847_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n888_;
  XNOR2_X1  g000(.A(G85gat), .B(G92gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT9), .ZN(new_n204_));
  XOR2_X1   g003(.A(KEYINPUT10), .B(G99gat), .Z(new_n205_));
  INV_X1    g004(.A(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G85gat), .ZN(new_n208_));
  INV_X1    g007(.A(G92gat), .ZN(new_n209_));
  OR3_X1    g008(.A1(new_n208_), .A2(new_n209_), .A3(KEYINPUT9), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT6), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n204_), .A2(new_n207_), .A3(new_n210_), .A4(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n212_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT66), .ZN(new_n215_));
  INV_X1    g014(.A(G99gat), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n215_), .A2(new_n216_), .A3(new_n206_), .A4(KEYINPUT7), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT7), .ZN(new_n218_));
  OAI22_X1  g017(.A1(new_n218_), .A2(KEYINPUT66), .B1(G99gat), .B2(G106gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n215_), .A2(KEYINPUT7), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n217_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT67), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT67), .ZN(new_n223_));
  OAI211_X1 g022(.A(new_n217_), .B(new_n223_), .C1(new_n219_), .C2(new_n220_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n214_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n225_));
  OAI211_X1 g024(.A(KEYINPUT68), .B(KEYINPUT8), .C1(new_n225_), .C2(new_n202_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n221_), .A2(new_n212_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT8), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n228_), .A3(new_n203_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n226_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n224_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n216_), .A2(new_n206_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n215_), .A2(KEYINPUT7), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n218_), .A2(KEYINPUT66), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n223_), .B1(new_n235_), .B2(new_n217_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n212_), .B1(new_n231_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(new_n203_), .ZN(new_n238_));
  AOI21_X1  g037(.A(KEYINPUT68), .B1(new_n238_), .B2(KEYINPUT8), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n213_), .B1(new_n230_), .B2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G29gat), .B(G36gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT70), .ZN(new_n242_));
  XOR2_X1   g041(.A(G43gat), .B(G50gat), .Z(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT71), .B(KEYINPUT15), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT35), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G232gat), .A2(G233gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT34), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  AOI22_X1  g049(.A1(new_n240_), .A2(new_n246_), .B1(new_n247_), .B2(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n247_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT8), .B1(new_n225_), .B2(new_n202_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(new_n226_), .A3(new_n229_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(new_n244_), .A3(new_n213_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n251_), .A2(new_n253_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT73), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n251_), .A2(KEYINPUT73), .A3(new_n253_), .A4(new_n258_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n251_), .A2(new_n258_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(new_n252_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT72), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n253_), .B1(new_n251_), .B2(new_n258_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT72), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n263_), .A2(new_n267_), .A3(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(G190gat), .B(G218gat), .Z(new_n271_));
  XNOR2_X1  g070(.A(G134gat), .B(G162gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT36), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n270_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n273_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n276_), .A2(KEYINPUT36), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n263_), .A2(new_n267_), .A3(new_n269_), .A4(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n275_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(G176gat), .ZN(new_n281_));
  INV_X1    g080(.A(G169gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(KEYINPUT85), .B1(new_n282_), .B2(KEYINPUT22), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT22), .B(G169gat), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n281_), .B(new_n283_), .C1(new_n284_), .C2(KEYINPUT85), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT86), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT23), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n290_), .B1(G183gat), .B2(G190gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n285_), .A2(new_n286_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n287_), .A2(new_n288_), .A3(new_n291_), .A4(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT84), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n296_), .A2(KEYINPUT24), .A3(new_n288_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n294_), .B(KEYINPUT84), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT24), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT25), .B(G183gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT26), .B(G190gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n297_), .A2(new_n300_), .A3(new_n303_), .A4(new_n290_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n293_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT30), .ZN(new_n306_));
  XOR2_X1   g105(.A(G71gat), .B(G99gat), .Z(new_n307_));
  NAND2_X1  g106(.A1(G227gat), .A2(G233gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G15gat), .B(G43gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT87), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n309_), .B(new_n311_), .Z(new_n312_));
  AND2_X1   g111(.A1(new_n306_), .A2(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n306_), .A2(new_n312_), .ZN(new_n314_));
  OR3_X1    g113(.A1(new_n313_), .A2(new_n314_), .A3(KEYINPUT31), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT31), .B1(new_n313_), .B2(new_n314_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G127gat), .B(G134gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G113gat), .B(G120gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n317_), .A2(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT89), .ZN(new_n324_));
  AOI21_X1  g123(.A(KEYINPUT1), .B1(G155gat), .B2(G162gat), .ZN(new_n325_));
  AND3_X1   g124(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n324_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G141gat), .A2(G148gat), .ZN(new_n328_));
  NOR2_X1   g127(.A1(G141gat), .A2(G148gat), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT88), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n327_), .A2(new_n328_), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n329_), .B(KEYINPUT3), .Z(new_n334_));
  XOR2_X1   g133(.A(new_n328_), .B(KEYINPUT2), .Z(new_n335_));
  OAI211_X1 g134(.A(new_n324_), .B(new_n333_), .C1(new_n334_), .C2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n332_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(new_n320_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n337_), .A2(new_n321_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(KEYINPUT4), .A3(new_n340_), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n340_), .A2(KEYINPUT4), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G225gat), .A2(G233gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n341_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n345_));
  XOR2_X1   g144(.A(G1gat), .B(G29gat), .Z(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT0), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(G57gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(new_n208_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n339_), .A2(new_n340_), .A3(new_n343_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n345_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT98), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT98), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n345_), .A2(new_n350_), .A3(new_n354_), .A4(new_n351_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n345_), .A2(new_n351_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n349_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n353_), .A2(new_n355_), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n315_), .A2(new_n320_), .A3(new_n316_), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n322_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(G22gat), .B(G50gat), .Z(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT29), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n364_), .B1(new_n332_), .B2(new_n336_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  XOR2_X1   g165(.A(G197gat), .B(G204gat), .Z(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT21), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT90), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G211gat), .B(G218gat), .ZN(new_n370_));
  OR3_X1    g169(.A1(new_n368_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n369_), .B1(new_n368_), .B2(new_n370_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n368_), .A2(new_n370_), .ZN(new_n374_));
  OR2_X1    g173(.A1(new_n367_), .A2(KEYINPUT21), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n373_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G228gat), .A2(G233gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT91), .ZN(new_n379_));
  OR2_X1    g178(.A1(new_n378_), .A2(KEYINPUT91), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n366_), .A2(new_n377_), .A3(new_n379_), .A4(new_n380_), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n371_), .A2(new_n372_), .B1(new_n375_), .B2(new_n374_), .ZN(new_n382_));
  OAI211_X1 g181(.A(KEYINPUT91), .B(new_n378_), .C1(new_n382_), .C2(new_n365_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G78gat), .B(G106gat), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n381_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n384_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n363_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n387_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n389_), .A2(new_n385_), .A3(new_n362_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n338_), .A2(new_n364_), .ZN(new_n392_));
  XOR2_X1   g191(.A(new_n392_), .B(KEYINPUT28), .Z(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n391_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n388_), .A2(new_n390_), .A3(new_n393_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT27), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n284_), .A2(new_n281_), .ZN(new_n399_));
  XOR2_X1   g198(.A(new_n288_), .B(KEYINPUT92), .Z(new_n400_));
  NAND3_X1  g199(.A1(new_n291_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n304_), .A2(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT93), .B1(new_n377_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n305_), .A2(new_n377_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n402_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT93), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(new_n382_), .A3(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G226gat), .A2(G233gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT19), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT20), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n403_), .A2(new_n404_), .A3(new_n407_), .A4(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n305_), .A2(new_n382_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n405_), .A2(new_n377_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n410_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n409_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n412_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G8gat), .B(G36gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT18), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G64gat), .B(G92gat), .ZN(new_n420_));
  XOR2_X1   g219(.A(new_n419_), .B(new_n420_), .Z(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n417_), .A2(new_n422_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n412_), .B(new_n421_), .C1(new_n415_), .C2(new_n416_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n424_), .A2(KEYINPUT27), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n415_), .A2(new_n416_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n402_), .B(KEYINPUT96), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n382_), .ZN(new_n429_));
  XOR2_X1   g228(.A(KEYINPUT95), .B(KEYINPUT20), .Z(new_n430_));
  AOI21_X1  g229(.A(new_n430_), .B1(new_n305_), .B2(new_n377_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n416_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n422_), .B1(new_n427_), .B2(new_n432_), .ZN(new_n433_));
  AOI22_X1  g232(.A1(new_n398_), .A2(new_n425_), .B1(new_n426_), .B2(new_n433_), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n397_), .A2(new_n434_), .A3(KEYINPUT99), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT99), .B1(new_n397_), .B2(new_n434_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n361_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT33), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n352_), .A2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n339_), .A2(new_n340_), .A3(new_n344_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(new_n349_), .A3(new_n441_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n345_), .A2(new_n350_), .A3(KEYINPUT33), .A4(new_n351_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n439_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT94), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n444_), .A2(new_n445_), .A3(new_n424_), .A4(new_n423_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n421_), .A2(KEYINPUT32), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n447_), .B1(new_n427_), .B2(new_n432_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT97), .ZN(new_n449_));
  OR2_X1    g248(.A1(new_n417_), .A2(new_n447_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT97), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n451_), .B(new_n447_), .C1(new_n427_), .C2(new_n432_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n449_), .A2(new_n358_), .A3(new_n450_), .A4(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n439_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT94), .B1(new_n454_), .B2(new_n425_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n446_), .A2(new_n453_), .A3(new_n397_), .A4(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n434_), .A2(new_n359_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n397_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n322_), .A2(new_n360_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n456_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n280_), .B1(new_n437_), .B2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT102), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G57gat), .B(G64gat), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n464_), .A2(KEYINPUT11), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(KEYINPUT11), .ZN(new_n466_));
  XOR2_X1   g265(.A(G71gat), .B(G78gat), .Z(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  OR2_X1    g267(.A1(new_n466_), .A2(new_n467_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n213_), .B(new_n470_), .C1(new_n230_), .C2(new_n239_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G230gat), .A2(G233gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n471_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT69), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT69), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n471_), .A2(new_n477_), .A3(new_n474_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  AOI211_X1 g278(.A(KEYINPUT12), .B(new_n470_), .C1(new_n257_), .C2(new_n213_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT12), .ZN(new_n481_));
  INV_X1    g280(.A(new_n470_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n481_), .B1(new_n240_), .B2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n480_), .A2(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n479_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n240_), .A2(new_n482_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n474_), .B1(new_n486_), .B2(new_n471_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G120gat), .B(G148gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT5), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G176gat), .B(G204gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n489_), .B(new_n490_), .Z(new_n491_));
  OR3_X1    g290(.A1(new_n485_), .A2(new_n487_), .A3(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n491_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n494_), .A2(KEYINPUT13), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(KEYINPUT13), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  XOR2_X1   g297(.A(KEYINPUT76), .B(G8gat), .Z(new_n499_));
  INV_X1    g298(.A(G1gat), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT14), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G15gat), .B(G22gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G1gat), .B(G8gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT82), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(new_n507_), .A3(new_n244_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n244_), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT82), .B1(new_n509_), .B2(new_n505_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n511_), .B1(new_n506_), .B2(new_n244_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G229gat), .A2(G233gat), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n246_), .A2(new_n505_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT83), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n246_), .A2(KEYINPUT83), .A3(new_n505_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(new_n518_), .A3(new_n511_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n514_), .B1(new_n519_), .B2(new_n513_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G113gat), .B(G141gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G169gat), .B(G197gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n520_), .B(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n498_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G231gat), .A2(G233gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n470_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(new_n505_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n529_), .A2(KEYINPUT79), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G127gat), .B(G155gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT16), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT77), .ZN(new_n533_));
  XOR2_X1   g332(.A(G183gat), .B(G211gat), .Z(new_n534_));
  XOR2_X1   g333(.A(new_n534_), .B(KEYINPUT78), .Z(new_n535_));
  XNOR2_X1  g334(.A(new_n533_), .B(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT17), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n530_), .A2(new_n538_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n536_), .A2(new_n537_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n530_), .A2(new_n538_), .B1(new_n529_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n463_), .B1(new_n526_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n542_), .ZN(new_n544_));
  NOR4_X1   g343(.A1(new_n498_), .A2(KEYINPUT102), .A3(new_n525_), .A4(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n462_), .B1(new_n543_), .B2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(G1gat), .B1(new_n546_), .B2(new_n359_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT75), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n548_), .B1(new_n279_), .B2(KEYINPUT37), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT74), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n278_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n268_), .B(new_n266_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n552_), .A2(KEYINPUT74), .A3(new_n263_), .A4(new_n277_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n551_), .A2(new_n553_), .A3(new_n275_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(KEYINPUT37), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT37), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n275_), .A2(KEYINPUT75), .A3(new_n556_), .A4(new_n278_), .ZN(new_n557_));
  AND3_X1   g356(.A1(new_n549_), .A2(new_n555_), .A3(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n542_), .B(KEYINPUT80), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(new_n497_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT81), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n561_), .A2(KEYINPUT81), .A3(new_n497_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n437_), .A2(new_n461_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n525_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n566_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT100), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n566_), .A2(KEYINPUT100), .A3(new_n570_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n359_), .A2(G1gat), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT101), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT38), .ZN(new_n579_));
  AOI21_X1  g378(.A(KEYINPUT100), .B1(new_n566_), .B2(new_n570_), .ZN(new_n580_));
  AOI211_X1 g379(.A(new_n572_), .B(new_n569_), .C1(new_n564_), .C2(new_n565_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n582_), .A2(KEYINPUT101), .A3(new_n575_), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n578_), .A2(new_n579_), .A3(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n579_), .B1(new_n578_), .B2(new_n583_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n547_), .B1(new_n584_), .B2(new_n585_), .ZN(G1324gat));
  OAI21_X1  g385(.A(G8gat), .B1(new_n546_), .B2(new_n434_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT39), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT103), .ZN(new_n589_));
  INV_X1    g388(.A(new_n434_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(new_n499_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n589_), .B1(new_n582_), .B2(new_n592_), .ZN(new_n593_));
  NOR4_X1   g392(.A1(new_n580_), .A2(new_n581_), .A3(KEYINPUT103), .A4(new_n591_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n588_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT40), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  OAI211_X1 g396(.A(KEYINPUT40), .B(new_n588_), .C1(new_n593_), .C2(new_n594_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(G1325gat));
  OAI21_X1  g398(.A(G15gat), .B1(new_n546_), .B2(new_n460_), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n600_), .B(KEYINPUT41), .Z(new_n601_));
  INV_X1    g400(.A(new_n582_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n460_), .A2(G15gat), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n601_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT104), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n601_), .B(KEYINPUT104), .C1(new_n602_), .C2(new_n603_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(G1326gat));
  OR3_X1    g407(.A1(new_n602_), .A2(G22gat), .A3(new_n397_), .ZN(new_n609_));
  OAI21_X1  g408(.A(G22gat), .B1(new_n546_), .B2(new_n397_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n610_), .A2(KEYINPUT42), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(KEYINPUT42), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n609_), .B1(new_n611_), .B2(new_n612_), .ZN(G1327gat));
  NOR2_X1   g412(.A1(new_n279_), .A2(new_n559_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n526_), .A2(new_n567_), .A3(new_n614_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n615_), .A2(KEYINPUT107), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(KEYINPUT107), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(G29gat), .B1(new_n618_), .B2(new_n358_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n567_), .A2(new_n555_), .A3(new_n549_), .A4(new_n557_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT105), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n549_), .A2(new_n555_), .A3(new_n621_), .A4(new_n557_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n620_), .A2(KEYINPUT43), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT43), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n558_), .B(new_n567_), .C1(new_n621_), .C2(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n559_), .B1(new_n623_), .B2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(new_n526_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT44), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n629_), .A2(G29gat), .A3(new_n358_), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT106), .B1(new_n627_), .B2(new_n628_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT106), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n626_), .A2(new_n632_), .A3(KEYINPUT44), .A4(new_n526_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n619_), .B1(new_n630_), .B2(new_n634_), .ZN(G1328gat));
  INV_X1    g434(.A(G36gat), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n616_), .A2(new_n636_), .A3(new_n590_), .A4(new_n617_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT45), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n629_), .A2(new_n590_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n639_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n638_), .B1(new_n640_), .B2(new_n636_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT46), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  OAI211_X1 g442(.A(KEYINPUT46), .B(new_n638_), .C1(new_n640_), .C2(new_n636_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(G1329gat));
  INV_X1    g444(.A(new_n460_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n618_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(G43gat), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n634_), .A2(new_n629_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n646_), .A2(G43gat), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n649_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g452(.A(G50gat), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n618_), .A2(new_n654_), .A3(new_n458_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT108), .ZN(new_n656_));
  AOI22_X1  g455(.A1(new_n631_), .A2(new_n633_), .B1(new_n628_), .B2(new_n627_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(new_n458_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n656_), .B1(new_n658_), .B2(G50gat), .ZN(new_n659_));
  AOI211_X1 g458(.A(KEYINPUT108), .B(new_n654_), .C1(new_n657_), .C2(new_n458_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n655_), .B1(new_n659_), .B2(new_n660_), .ZN(G1331gat));
  NOR2_X1   g460(.A1(new_n497_), .A2(new_n568_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n662_), .A2(new_n462_), .A3(new_n559_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G57gat), .B1(new_n663_), .B2(new_n359_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n662_), .A2(new_n567_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(new_n561_), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n359_), .A2(G57gat), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n664_), .B1(new_n666_), .B2(new_n667_), .ZN(G1332gat));
  OAI21_X1  g467(.A(G64gat), .B1(new_n663_), .B2(new_n434_), .ZN(new_n669_));
  XOR2_X1   g468(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n434_), .A2(G64gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(new_n666_), .B2(new_n672_), .ZN(G1333gat));
  OAI21_X1  g472(.A(G71gat), .B1(new_n663_), .B2(new_n460_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT49), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n460_), .A2(G71gat), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n666_), .B2(new_n676_), .ZN(G1334gat));
  OAI21_X1  g476(.A(G78gat), .B1(new_n663_), .B2(new_n397_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT50), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n397_), .A2(G78gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n679_), .B1(new_n666_), .B2(new_n680_), .ZN(G1335gat));
  NAND2_X1  g480(.A1(new_n665_), .A2(new_n614_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n683_), .A2(new_n208_), .A3(new_n358_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n626_), .A2(new_n662_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT110), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT110), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n626_), .A2(new_n687_), .A3(new_n662_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n359_), .B1(new_n686_), .B2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n684_), .B1(new_n689_), .B2(new_n208_), .ZN(G1336gat));
  NAND3_X1  g489(.A1(new_n683_), .A2(new_n209_), .A3(new_n590_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n434_), .B1(new_n686_), .B2(new_n688_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n691_), .B1(new_n692_), .B2(new_n209_), .ZN(G1337gat));
  INV_X1    g492(.A(KEYINPUT112), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n683_), .A2(new_n205_), .A3(new_n646_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n460_), .B1(new_n686_), .B2(new_n688_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(new_n696_), .B2(new_n216_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n694_), .B1(new_n697_), .B2(KEYINPUT51), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n696_), .A2(new_n216_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT51), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n699_), .A2(KEYINPUT112), .A3(new_n700_), .A4(new_n695_), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n697_), .A2(KEYINPUT111), .A3(KEYINPUT51), .ZN(new_n702_));
  AOI21_X1  g501(.A(KEYINPUT111), .B1(new_n697_), .B2(KEYINPUT51), .ZN(new_n703_));
  OAI211_X1 g502(.A(new_n698_), .B(new_n701_), .C1(new_n702_), .C2(new_n703_), .ZN(G1338gat));
  NAND3_X1  g503(.A1(new_n683_), .A2(new_n206_), .A3(new_n458_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n626_), .A2(new_n458_), .A3(new_n662_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT52), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n706_), .A2(new_n707_), .A3(G106gat), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n707_), .B1(new_n706_), .B2(G106gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n705_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g511(.A(KEYINPUT59), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n646_), .B(new_n358_), .C1(new_n435_), .C2(new_n436_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n561_), .A2(new_n525_), .A3(new_n497_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT54), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n716_), .B(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n524_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n719_), .B1(new_n513_), .B2(new_n519_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n720_), .B1(new_n520_), .B2(new_n523_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n485_), .A2(new_n487_), .A3(new_n491_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT55), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n724_), .B1(new_n479_), .B2(new_n484_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n486_), .A2(KEYINPUT12), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n240_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND4_X1  g527(.A1(new_n728_), .A2(KEYINPUT55), .A3(new_n476_), .A4(new_n478_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n471_), .B1(new_n480_), .B2(new_n483_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n474_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n725_), .A2(new_n729_), .A3(new_n732_), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n733_), .A2(KEYINPUT56), .A3(new_n491_), .ZN(new_n734_));
  AOI21_X1  g533(.A(KEYINPUT56), .B1(new_n733_), .B2(new_n491_), .ZN(new_n735_));
  OAI211_X1 g534(.A(KEYINPUT58), .B(new_n723_), .C1(new_n734_), .C2(new_n735_), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n555_), .A2(new_n549_), .A3(new_n736_), .A4(new_n557_), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n734_), .A2(new_n735_), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT58), .B1(new_n738_), .B2(new_n723_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n737_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT57), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n525_), .A2(new_n722_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n735_), .A2(KEYINPUT113), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT113), .ZN(new_n745_));
  AOI211_X1 g544(.A(new_n745_), .B(KEYINPUT56), .C1(new_n733_), .C2(new_n491_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n733_), .A2(KEYINPUT56), .A3(new_n491_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT114), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n733_), .A2(KEYINPUT114), .A3(KEYINPUT56), .A4(new_n491_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n743_), .B1(new_n747_), .B2(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n721_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n741_), .B(new_n279_), .C1(new_n753_), .C2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n491_), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n476_), .B(new_n478_), .C1(new_n483_), .C2(new_n480_), .ZN(new_n757_));
  AOI22_X1  g556(.A1(new_n757_), .A2(new_n724_), .B1(new_n731_), .B2(new_n730_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n756_), .B1(new_n758_), .B2(new_n729_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n745_), .B1(new_n759_), .B2(KEYINPUT56), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n733_), .A2(new_n491_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT56), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n761_), .A2(KEYINPUT113), .A3(new_n762_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n760_), .A2(new_n763_), .A3(new_n750_), .A4(new_n751_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n754_), .B1(new_n764_), .B2(new_n742_), .ZN(new_n765_));
  OAI21_X1  g564(.A(KEYINPUT57), .B1(new_n765_), .B2(new_n280_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n740_), .B1(new_n755_), .B2(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n767_), .A2(new_n559_), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n713_), .B(new_n715_), .C1(new_n718_), .C2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n755_), .A2(new_n766_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n740_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT115), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT115), .ZN(new_n773_));
  AOI211_X1 g572(.A(new_n773_), .B(new_n740_), .C1(new_n755_), .C2(new_n766_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n544_), .B1(new_n772_), .B2(new_n774_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n716_), .B(KEYINPUT54), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n714_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n769_), .B1(new_n777_), .B2(new_n713_), .ZN(new_n778_));
  OAI21_X1  g577(.A(G113gat), .B1(new_n778_), .B2(new_n525_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n775_), .A2(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n715_), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n525_), .A2(G113gat), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n779_), .B1(new_n781_), .B2(new_n782_), .ZN(G1340gat));
  XOR2_X1   g582(.A(KEYINPUT116), .B(G120gat), .Z(new_n784_));
  NOR2_X1   g583(.A1(new_n497_), .A2(new_n784_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n780_), .B(new_n715_), .C1(KEYINPUT60), .C2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n498_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n784_), .B1(new_n787_), .B2(new_n778_), .ZN(new_n788_));
  OR2_X1    g587(.A1(new_n786_), .A2(KEYINPUT60), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(G1341gat));
  AOI21_X1  g589(.A(G127gat), .B1(new_n777_), .B2(new_n559_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n778_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(KEYINPUT117), .B(G127gat), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n544_), .A2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n791_), .B1(new_n792_), .B2(new_n794_), .ZN(G1342gat));
  NAND2_X1  g594(.A1(new_n558_), .A2(G134gat), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT118), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n769_), .B(new_n797_), .C1(new_n777_), .C2(new_n713_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n764_), .A2(new_n742_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n754_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n741_), .B1(new_n801_), .B2(new_n279_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n765_), .A2(KEYINPUT57), .A3(new_n280_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n771_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n773_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n767_), .A2(KEYINPUT115), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n542_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n280_), .B(new_n715_), .C1(new_n807_), .C2(new_n718_), .ZN(new_n808_));
  INV_X1    g607(.A(G134gat), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n798_), .A2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT119), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT119), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n798_), .A2(new_n813_), .A3(new_n810_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(G1343gat));
  NOR2_X1   g614(.A1(new_n807_), .A2(new_n718_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n646_), .A2(new_n397_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n817_), .A2(new_n358_), .A3(new_n434_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(KEYINPUT120), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n816_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n568_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n498_), .ZN(new_n823_));
  XOR2_X1   g622(.A(KEYINPUT121), .B(G148gat), .Z(new_n824_));
  XNOR2_X1  g623(.A(new_n823_), .B(new_n824_), .ZN(G1345gat));
  NAND2_X1  g624(.A1(new_n820_), .A2(new_n559_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(KEYINPUT61), .B(G155gat), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n826_), .B(new_n827_), .ZN(G1346gat));
  INV_X1    g627(.A(new_n820_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n558_), .ZN(new_n830_));
  OAI21_X1  g629(.A(G162gat), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(G162gat), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n820_), .A2(new_n832_), .A3(new_n280_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(G1347gat));
  NAND2_X1  g633(.A1(new_n361_), .A2(new_n590_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n835_), .A2(new_n458_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n836_), .B1(new_n718_), .B2(new_n768_), .ZN(new_n837_));
  OAI21_X1  g636(.A(G169gat), .B1(new_n837_), .B2(new_n525_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT62), .ZN(new_n839_));
  OR2_X1    g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n839_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n837_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n842_), .A2(new_n568_), .A3(new_n284_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n840_), .A2(new_n841_), .A3(new_n843_), .ZN(G1348gat));
  AOI21_X1  g643(.A(G176gat), .B1(new_n842_), .B2(new_n498_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n816_), .A2(new_n458_), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n497_), .A2(new_n281_), .A3(new_n835_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n845_), .B1(new_n846_), .B2(new_n847_), .ZN(G1349gat));
  NOR2_X1   g647(.A1(new_n544_), .A2(new_n301_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n836_), .B(new_n849_), .C1(new_n718_), .C2(new_n768_), .ZN(new_n850_));
  XOR2_X1   g649(.A(new_n850_), .B(KEYINPUT122), .Z(new_n851_));
  INV_X1    g650(.A(new_n835_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n780_), .A2(new_n397_), .A3(new_n559_), .A4(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT123), .ZN(new_n855_));
  AOI21_X1  g654(.A(G183gat), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n853_), .A2(KEYINPUT123), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n851_), .B1(new_n856_), .B2(new_n857_), .ZN(G1350gat));
  OAI21_X1  g657(.A(G190gat), .B1(new_n837_), .B2(new_n830_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n280_), .A2(new_n302_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n837_), .B2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT124), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n861_), .B(new_n862_), .ZN(G1351gat));
  INV_X1    g662(.A(new_n817_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n864_), .A2(new_n358_), .A3(new_n434_), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n568_), .B(new_n865_), .C1(new_n807_), .C2(new_n718_), .ZN(new_n866_));
  INV_X1    g665(.A(G197gat), .ZN(new_n867_));
  OAI21_X1  g666(.A(KEYINPUT125), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n865_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n869_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT125), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n870_), .A2(new_n871_), .A3(G197gat), .A4(new_n568_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n868_), .A2(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(G197gat), .B1(new_n870_), .B2(new_n568_), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n874_), .A2(KEYINPUT126), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(KEYINPUT126), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n873_), .B1(new_n875_), .B2(new_n876_), .ZN(G1352gat));
  NAND2_X1  g676(.A1(new_n870_), .A2(new_n498_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g678(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n542_), .A2(new_n880_), .ZN(new_n881_));
  XOR2_X1   g680(.A(new_n881_), .B(KEYINPUT127), .Z(new_n882_));
  NAND2_X1  g681(.A1(new_n870_), .A2(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n884_));
  XOR2_X1   g683(.A(new_n883_), .B(new_n884_), .Z(G1354gat));
  INV_X1    g684(.A(new_n870_), .ZN(new_n886_));
  OR3_X1    g685(.A1(new_n886_), .A2(G218gat), .A3(new_n279_), .ZN(new_n887_));
  OAI21_X1  g686(.A(G218gat), .B1(new_n886_), .B2(new_n830_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1355gat));
endmodule


