//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 1 0 0 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 1 0 1 0 0 1 1 0 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 1 1 1 1 1 1 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n771_, new_n772_, new_n773_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n932_, new_n933_, new_n934_, new_n935_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n948_, new_n949_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n957_, new_n958_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT23), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND3_X1  g003(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n205_));
  AND2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT24), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT24), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n211_), .A2(new_n207_), .ZN(new_n212_));
  AND3_X1   g011(.A1(new_n206_), .A2(new_n209_), .A3(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT26), .B(G190gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT76), .ZN(new_n215_));
  INV_X1    g014(.A(G183gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT25), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n216_), .A2(KEYINPUT25), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n214_), .B(new_n217_), .C1(new_n218_), .C2(new_n215_), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n204_), .B(new_n205_), .C1(G183gat), .C2(G190gat), .ZN(new_n220_));
  AND2_X1   g019(.A1(new_n220_), .A2(new_n210_), .ZN(new_n221_));
  INV_X1    g020(.A(G176gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT77), .ZN(new_n223_));
  INV_X1    g022(.A(G169gat), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n223_), .B1(new_n224_), .B2(KEYINPUT22), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT22), .B(G169gat), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n222_), .B(new_n225_), .C1(new_n226_), .C2(new_n223_), .ZN(new_n227_));
  AOI22_X1  g026(.A1(new_n213_), .A2(new_n219_), .B1(new_n221_), .B2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G227gat), .A2(G233gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(G15gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n228_), .B(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G71gat), .B(G99gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(G43gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT78), .B(KEYINPUT30), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n231_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n231_), .A2(new_n236_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G127gat), .B(G134gat), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  XOR2_X1   g040(.A(G113gat), .B(G120gat), .Z(new_n242_));
  INV_X1    g041(.A(KEYINPUT80), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(new_n242_), .A3(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G113gat), .B(G120gat), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT80), .B1(new_n240_), .B2(new_n245_), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n240_), .A2(new_n245_), .A3(KEYINPUT79), .ZN(new_n247_));
  AOI21_X1  g046(.A(KEYINPUT79), .B1(new_n240_), .B2(new_n245_), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n244_), .B(new_n246_), .C1(new_n247_), .C2(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(KEYINPUT81), .B(KEYINPUT31), .Z(new_n250_));
  XOR2_X1   g049(.A(new_n249_), .B(new_n250_), .Z(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n239_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n237_), .A2(new_n238_), .A3(new_n251_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT96), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT93), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n258_), .A2(KEYINPUT33), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G225gat), .A2(G233gat), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n249_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(G155gat), .A2(G162gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G155gat), .A2(G162gat), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n264_), .B1(KEYINPUT1), .B2(new_n265_), .ZN(new_n266_));
  OR2_X1    g065(.A1(new_n265_), .A2(KEYINPUT1), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G141gat), .A2(G148gat), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(G141gat), .A2(G148gat), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n268_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT3), .ZN(new_n274_));
  INV_X1    g073(.A(G141gat), .ZN(new_n275_));
  INV_X1    g074(.A(G148gat), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n274_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT2), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n269_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n277_), .A2(new_n279_), .A3(new_n280_), .A4(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT82), .ZN(new_n283_));
  XOR2_X1   g082(.A(G155gat), .B(G162gat), .Z(new_n284_));
  AND3_X1   g083(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n283_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n273_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT4), .B1(new_n263_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n240_), .B(new_n245_), .ZN(new_n290_));
  OAI211_X1 g089(.A(new_n273_), .B(new_n290_), .C1(new_n285_), .C2(new_n286_), .ZN(new_n291_));
  AOI211_X1 g090(.A(new_n270_), .B(new_n271_), .C1(new_n266_), .C2(new_n267_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n282_), .A2(new_n284_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT82), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n292_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n291_), .B1(new_n296_), .B2(new_n249_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT4), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n262_), .B(new_n289_), .C1(new_n298_), .C2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n261_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G1gat), .B(G29gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(G85gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT0), .B(G57gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n260_), .B1(new_n302_), .B2(new_n307_), .ZN(new_n308_));
  AOI211_X1 g107(.A(new_n306_), .B(new_n259_), .C1(new_n300_), .C2(new_n301_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(G8gat), .B(G36gat), .Z(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT18), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G64gat), .B(G92gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G226gat), .A2(G233gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT19), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT91), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT20), .ZN(new_n320_));
  INV_X1    g119(.A(G204gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(G197gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT85), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n321_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(KEYINPUT85), .A2(G204gat), .ZN(new_n325_));
  AOI21_X1  g124(.A(G197gat), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT86), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n322_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(G197gat), .ZN(new_n329_));
  AND2_X1   g128(.A1(KEYINPUT85), .A2(G204gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(KEYINPUT85), .A2(G204gat), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n327_), .B(new_n329_), .C1(new_n330_), .C2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT21), .B1(new_n328_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(G218gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(G211gat), .ZN(new_n336_));
  INV_X1    g135(.A(G211gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(G218gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n324_), .A2(KEYINPUT87), .A3(G197gat), .A4(new_n325_), .ZN(new_n340_));
  NOR3_X1   g139(.A1(new_n330_), .A2(new_n331_), .A3(new_n329_), .ZN(new_n341_));
  AOI21_X1  g140(.A(KEYINPUT87), .B1(new_n329_), .B2(G204gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n340_), .B1(new_n341_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT21), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n339_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n345_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n340_), .B(new_n347_), .C1(new_n341_), .C2(new_n343_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT88), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n324_), .A2(new_n325_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n342_), .B1(new_n351_), .B2(new_n329_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n352_), .A2(KEYINPUT88), .A3(new_n340_), .A4(new_n347_), .ZN(new_n353_));
  AOI22_X1  g152(.A1(new_n334_), .A2(new_n346_), .B1(new_n350_), .B2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n320_), .B1(new_n354_), .B2(new_n228_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n346_), .A2(new_n334_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n350_), .A2(new_n353_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n226_), .A2(new_n222_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n359_), .A2(new_n220_), .A3(new_n210_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT25), .B(G183gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n214_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n362_), .A2(new_n206_), .A3(new_n209_), .ZN(new_n363_));
  AND3_X1   g162(.A1(new_n210_), .A2(KEYINPUT92), .A3(KEYINPUT24), .ZN(new_n364_));
  AOI21_X1  g163(.A(KEYINPUT92), .B1(new_n210_), .B2(KEYINPUT24), .ZN(new_n365_));
  NOR3_X1   g164(.A1(new_n364_), .A2(new_n365_), .A3(new_n207_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n360_), .B1(new_n363_), .B2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n358_), .A2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n319_), .B1(new_n355_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n317_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n370_), .B1(new_n358_), .B2(new_n367_), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT20), .B1(new_n354_), .B2(new_n228_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n315_), .B1(new_n369_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n263_), .A2(new_n287_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n299_), .B1(new_n375_), .B2(new_n291_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n261_), .B1(new_n376_), .B2(new_n288_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n298_), .A2(KEYINPUT94), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT94), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n262_), .B1(new_n297_), .B2(new_n379_), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n377_), .B(new_n306_), .C1(new_n378_), .C2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n228_), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT20), .B1(new_n358_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n367_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n354_), .A2(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n318_), .B1(new_n383_), .B2(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n320_), .B1(new_n358_), .B2(new_n382_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n317_), .B1(new_n354_), .B2(new_n384_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n386_), .A2(new_n314_), .A3(new_n389_), .ZN(new_n390_));
  AND3_X1   g189(.A1(new_n374_), .A2(new_n381_), .A3(new_n390_), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n376_), .A2(new_n261_), .A3(new_n288_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n301_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n307_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n300_), .A2(new_n306_), .A3(new_n301_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n369_), .A2(new_n373_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n314_), .A2(KEYINPUT32), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n394_), .A2(new_n395_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT90), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n358_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n354_), .A2(KEYINPUT90), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT95), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n367_), .A2(new_n402_), .ZN(new_n403_));
  OAI211_X1 g202(.A(new_n360_), .B(KEYINPUT95), .C1(new_n363_), .C2(new_n366_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n400_), .A2(new_n401_), .A3(new_n403_), .A4(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n370_), .B1(new_n405_), .B2(new_n387_), .ZN(new_n406_));
  NOR3_X1   g205(.A1(new_n383_), .A2(new_n318_), .A3(new_n385_), .ZN(new_n407_));
  OAI211_X1 g206(.A(KEYINPUT32), .B(new_n314_), .C1(new_n406_), .C2(new_n407_), .ZN(new_n408_));
  AOI22_X1  g207(.A1(new_n310_), .A2(new_n391_), .B1(new_n398_), .B2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT29), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n296_), .A2(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(KEYINPUT83), .B(KEYINPUT28), .Z(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n411_), .B(new_n413_), .ZN(new_n414_));
  XOR2_X1   g213(.A(G22gat), .B(G50gat), .Z(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n414_), .B(new_n416_), .ZN(new_n417_));
  XOR2_X1   g216(.A(G78gat), .B(G106gat), .Z(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT89), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n420_), .B1(new_n296_), .B2(new_n410_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n287_), .A2(KEYINPUT89), .A3(KEYINPUT29), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n356_), .A2(KEYINPUT90), .A3(new_n357_), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT90), .B1(new_n356_), .B2(new_n357_), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n421_), .B(new_n422_), .C1(new_n423_), .C2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(G233gat), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n426_), .A2(KEYINPUT84), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(KEYINPUT84), .ZN(new_n428_));
  OAI21_X1  g227(.A(G228gat), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n425_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n287_), .A2(KEYINPUT29), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n358_), .A2(new_n429_), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n419_), .B1(new_n431_), .B2(new_n434_), .ZN(new_n435_));
  AOI211_X1 g234(.A(new_n418_), .B(new_n433_), .C1(new_n425_), .C2(new_n430_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n417_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n400_), .A2(new_n401_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n421_), .A2(new_n422_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n429_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n418_), .B1(new_n440_), .B2(new_n433_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n414_), .B(new_n415_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n431_), .A2(new_n419_), .A3(new_n434_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n441_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n437_), .A2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n257_), .B1(new_n409_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT98), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n403_), .A2(new_n404_), .ZN(new_n448_));
  NOR3_X1   g247(.A1(new_n423_), .A2(new_n424_), .A3(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n317_), .B1(new_n449_), .B2(new_n372_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n407_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n314_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n390_), .A2(KEYINPUT27), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n447_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n315_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n455_), .A2(KEYINPUT98), .A3(KEYINPUT27), .A4(new_n390_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT97), .ZN(new_n458_));
  NOR3_X1   g257(.A1(new_n392_), .A2(new_n307_), .A3(new_n393_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n306_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n458_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n394_), .A2(KEYINPUT97), .A3(new_n395_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT99), .B(KEYINPUT27), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n465_), .B1(new_n374_), .B2(new_n390_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n457_), .A2(new_n463_), .A3(new_n445_), .A4(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n394_), .A2(new_n259_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n460_), .A2(new_n260_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n374_), .A2(new_n381_), .A3(new_n390_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n386_), .A2(new_n389_), .A3(new_n397_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n473_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n397_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n475_));
  OAI22_X1  g274(.A1(new_n471_), .A2(new_n472_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n476_), .A2(KEYINPUT96), .A3(new_n444_), .A4(new_n437_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n446_), .A2(new_n468_), .A3(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n466_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n437_), .A2(new_n255_), .A3(new_n444_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n479_), .A2(new_n480_), .A3(new_n463_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT100), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT100), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n479_), .A2(new_n480_), .A3(new_n483_), .A4(new_n463_), .ZN(new_n484_));
  AOI22_X1  g283(.A1(new_n256_), .A2(new_n478_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G57gat), .B(G64gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT11), .ZN(new_n487_));
  XOR2_X1   g286(.A(G71gat), .B(G78gat), .Z(new_n488_));
  NOR2_X1   g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n487_), .A2(new_n488_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n486_), .A2(KEYINPUT11), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n489_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT12), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G99gat), .A2(G106gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT6), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT6), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n497_), .A2(G99gat), .A3(G106gat), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT65), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n496_), .A2(new_n498_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT65), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(G99gat), .A2(G106gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT7), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n500_), .A2(new_n503_), .A3(new_n505_), .ZN(new_n506_));
  XOR2_X1   g305(.A(G85gat), .B(G92gat), .Z(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n508_), .A2(KEYINPUT8), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n506_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT7), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n504_), .B(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n507_), .B1(new_n512_), .B2(new_n499_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT8), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n510_), .A2(new_n514_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n500_), .A2(new_n503_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT67), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT10), .B(G99gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT64), .B(G106gat), .ZN(new_n519_));
  OR2_X1    g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(G85gat), .ZN(new_n521_));
  INV_X1    g320(.A(G92gat), .ZN(new_n522_));
  NOR3_X1   g321(.A1(new_n521_), .A2(new_n522_), .A3(KEYINPUT9), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n523_), .B1(new_n507_), .B2(KEYINPUT9), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n516_), .A2(new_n517_), .A3(new_n520_), .A4(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n520_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n500_), .A2(new_n503_), .ZN(new_n527_));
  OAI21_X1  g326(.A(KEYINPUT67), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n515_), .A2(KEYINPUT66), .B1(new_n525_), .B2(new_n528_), .ZN(new_n529_));
  AOI22_X1  g328(.A1(new_n506_), .A2(new_n509_), .B1(new_n513_), .B2(KEYINPUT8), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT66), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n494_), .B1(new_n529_), .B2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n526_), .A2(new_n527_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n530_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n493_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n534_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n536_), .B1(new_n515_), .B2(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n537_), .B1(new_n539_), .B2(KEYINPUT12), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n533_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G230gat), .A2(G233gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n542_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n530_), .A2(new_n534_), .A3(new_n493_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n544_), .B1(new_n539_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(G120gat), .B(G148gat), .Z(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G176gat), .B(G204gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n547_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n552_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n543_), .A2(new_n546_), .A3(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n553_), .A2(KEYINPUT69), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT69), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n547_), .A2(new_n557_), .A3(new_n552_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT13), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n556_), .A2(KEYINPUT13), .A3(new_n558_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G29gat), .B(G36gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G43gat), .B(G50gat), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n566_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT15), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G15gat), .B(G22gat), .ZN(new_n571_));
  INV_X1    g370(.A(G1gat), .ZN(new_n572_));
  INV_X1    g371(.A(G8gat), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT14), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n571_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G1gat), .B(G8gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n570_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G229gat), .A2(G233gat), .ZN(new_n579_));
  INV_X1    g378(.A(new_n577_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(new_n569_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n578_), .A2(new_n579_), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n569_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n577_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n585_), .A2(G229gat), .A3(G233gat), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n582_), .A2(new_n586_), .ZN(new_n587_));
  XOR2_X1   g386(.A(G113gat), .B(G141gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT74), .ZN(new_n589_));
  XOR2_X1   g388(.A(G169gat), .B(G197gat), .Z(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n587_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n587_), .A2(new_n591_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT75), .ZN(new_n595_));
  NOR3_X1   g394(.A1(new_n485_), .A2(new_n564_), .A3(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G232gat), .A2(G233gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(KEYINPUT71), .B1(new_n535_), .B2(new_n569_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT71), .ZN(new_n601_));
  NOR4_X1   g400(.A1(new_n530_), .A2(new_n534_), .A3(new_n601_), .A4(new_n583_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n570_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n604_), .B1(new_n529_), .B2(new_n532_), .ZN(new_n605_));
  OAI211_X1 g404(.A(KEYINPUT35), .B(new_n599_), .C1(new_n603_), .C2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n602_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n515_), .A2(new_n538_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n601_), .B1(new_n608_), .B2(new_n583_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n515_), .A2(KEYINPUT66), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n525_), .A2(new_n528_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(new_n612_), .A3(new_n532_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n570_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n599_), .A2(KEYINPUT35), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n599_), .A2(KEYINPUT35), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n610_), .A2(new_n614_), .A3(new_n615_), .A4(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n606_), .A2(new_n617_), .A3(KEYINPUT73), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G190gat), .B(G218gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT72), .ZN(new_n620_));
  XOR2_X1   g419(.A(G134gat), .B(G162gat), .Z(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT36), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n618_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n624_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n606_), .A2(new_n617_), .A3(KEYINPUT73), .A4(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n606_), .A2(new_n617_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n622_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(KEYINPUT36), .A3(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n628_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT37), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT37), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n628_), .A2(new_n634_), .A3(new_n631_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n580_), .B(new_n493_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(G231gat), .A2(G233gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT17), .ZN(new_n640_));
  XOR2_X1   g439(.A(G127gat), .B(G155gat), .Z(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT16), .ZN(new_n642_));
  XNOR2_X1  g441(.A(G183gat), .B(G211gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(new_n644_));
  OR3_X1    g443(.A1(new_n639_), .A2(new_n640_), .A3(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(KEYINPUT17), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n639_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n636_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n596_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n463_), .B(KEYINPUT101), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT38), .ZN(new_n653_));
  AOI21_X1  g452(.A(G1gat), .B1(new_n653_), .B2(KEYINPUT102), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n651_), .A2(new_n652_), .A3(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n653_), .A2(KEYINPUT102), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n655_), .B(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n485_), .A2(new_n632_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n594_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n564_), .A2(new_n648_), .A3(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G1gat), .B1(new_n661_), .B2(new_n463_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT103), .Z(new_n663_));
  NAND2_X1  g462(.A1(new_n657_), .A2(new_n663_), .ZN(G1324gat));
  INV_X1    g463(.A(new_n479_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n651_), .A2(new_n573_), .A3(new_n665_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n661_), .A2(KEYINPUT104), .A3(new_n479_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n667_), .A2(new_n573_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT39), .ZN(new_n669_));
  OAI21_X1  g468(.A(KEYINPUT104), .B1(new_n661_), .B2(new_n479_), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n668_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n669_), .B1(new_n668_), .B2(new_n670_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n666_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT40), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  OAI211_X1 g474(.A(KEYINPUT40), .B(new_n666_), .C1(new_n671_), .C2(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1325gat));
  OAI21_X1  g476(.A(G15gat), .B1(new_n661_), .B2(new_n256_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT41), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n650_), .A2(G15gat), .A3(new_n256_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1326gat));
  INV_X1    g480(.A(new_n445_), .ZN(new_n682_));
  OAI21_X1  g481(.A(G22gat), .B1(new_n661_), .B2(new_n682_), .ZN(new_n683_));
  XOR2_X1   g482(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n684_));
  XNOR2_X1  g483(.A(new_n683_), .B(new_n684_), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n682_), .A2(G22gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n685_), .B1(new_n650_), .B2(new_n686_), .ZN(G1327gat));
  INV_X1    g486(.A(new_n632_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n648_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n596_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n463_), .ZN(new_n693_));
  AOI21_X1  g492(.A(G29gat), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT107), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n563_), .A2(new_n648_), .A3(new_n594_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n697_), .B1(new_n636_), .B2(KEYINPUT106), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n628_), .A2(new_n634_), .A3(new_n631_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n634_), .B1(new_n628_), .B2(new_n631_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n698_), .B1(new_n485_), .B2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n478_), .A2(new_n256_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n482_), .A2(new_n484_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT106), .ZN(new_n706_));
  OAI21_X1  g505(.A(KEYINPUT43), .B1(new_n701_), .B2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n705_), .A2(new_n636_), .A3(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n696_), .B1(new_n702_), .B2(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n695_), .B1(new_n709_), .B2(KEYINPUT44), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n485_), .A2(new_n698_), .A3(new_n701_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n707_), .B1(new_n705_), .B2(new_n636_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  OAI211_X1 g513(.A(KEYINPUT107), .B(new_n711_), .C1(new_n714_), .C2(new_n696_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n696_), .ZN(new_n716_));
  OAI211_X1 g515(.A(KEYINPUT44), .B(new_n716_), .C1(new_n712_), .C2(new_n713_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT108), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n709_), .A2(new_n719_), .A3(KEYINPUT44), .ZN(new_n720_));
  AOI22_X1  g519(.A1(new_n710_), .A2(new_n715_), .B1(new_n718_), .B2(new_n720_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n652_), .A2(G29gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n694_), .B1(new_n721_), .B2(new_n722_), .ZN(G1328gat));
  INV_X1    g522(.A(KEYINPUT46), .ZN(new_n724_));
  INV_X1    g523(.A(G36gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n721_), .B2(new_n665_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n692_), .A2(new_n725_), .A3(new_n665_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT45), .Z(new_n728_));
  OAI21_X1  g527(.A(new_n724_), .B1(new_n726_), .B2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n715_), .A2(new_n710_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n718_), .A2(new_n720_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n731_), .A3(new_n665_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(G36gat), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n727_), .B(KEYINPUT45), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n733_), .A2(KEYINPUT46), .A3(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n729_), .A2(new_n735_), .ZN(G1329gat));
  NAND4_X1  g535(.A1(new_n730_), .A2(new_n731_), .A3(G43gat), .A4(new_n255_), .ZN(new_n737_));
  INV_X1    g536(.A(G43gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n738_), .B1(new_n691_), .B2(new_n256_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT47), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT47), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n737_), .A2(new_n742_), .A3(new_n739_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1330gat));
  OR3_X1    g543(.A1(new_n691_), .A2(G50gat), .A3(new_n682_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n721_), .A2(new_n746_), .A3(new_n445_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(G50gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n746_), .B1(new_n721_), .B2(new_n445_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n745_), .B1(new_n748_), .B2(new_n749_), .ZN(G1331gat));
  NAND2_X1  g549(.A1(new_n595_), .A2(new_n689_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n705_), .A2(new_n688_), .A3(new_n564_), .A4(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(G57gat), .B1(new_n753_), .B2(new_n463_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n563_), .A2(new_n594_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n705_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n649_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT110), .ZN(new_n758_));
  INV_X1    g557(.A(new_n652_), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n759_), .A2(G57gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n754_), .B1(new_n758_), .B2(new_n760_), .ZN(G1332gat));
  OAI21_X1  g560(.A(G64gat), .B1(new_n753_), .B2(new_n479_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT48), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n479_), .A2(G64gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n758_), .B2(new_n764_), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT111), .Z(G1333gat));
  OAI21_X1  g565(.A(G71gat), .B1(new_n753_), .B2(new_n256_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT49), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n256_), .A2(G71gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n768_), .B1(new_n758_), .B2(new_n769_), .ZN(G1334gat));
  OAI21_X1  g569(.A(G78gat), .B1(new_n753_), .B2(new_n682_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT50), .ZN(new_n772_));
  OR2_X1    g571(.A1(new_n682_), .A2(G78gat), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n772_), .B1(new_n758_), .B2(new_n773_), .ZN(G1335gat));
  NAND2_X1  g573(.A1(new_n702_), .A2(new_n708_), .ZN(new_n775_));
  OR2_X1    g574(.A1(new_n775_), .A2(KEYINPUT112), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(KEYINPUT112), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n755_), .A2(new_n648_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n776_), .A2(new_n777_), .A3(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(G85gat), .B1(new_n780_), .B2(new_n463_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n756_), .A2(new_n690_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n652_), .A2(new_n521_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n781_), .B1(new_n782_), .B2(new_n783_), .ZN(G1336gat));
  OAI21_X1  g583(.A(G92gat), .B1(new_n780_), .B2(new_n479_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n665_), .A2(new_n522_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n785_), .B1(new_n782_), .B2(new_n786_), .ZN(G1337gat));
  OAI21_X1  g586(.A(G99gat), .B1(new_n780_), .B2(new_n256_), .ZN(new_n788_));
  OR3_X1    g587(.A1(new_n782_), .A2(new_n518_), .A3(new_n256_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT51), .ZN(G1338gat));
  OR3_X1    g590(.A1(new_n782_), .A2(new_n519_), .A3(new_n682_), .ZN(new_n792_));
  INV_X1    g591(.A(G106gat), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n778_), .A2(new_n682_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n775_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n795_), .A2(new_n796_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n792_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI21_X1  g599(.A(new_n591_), .B1(new_n585_), .B2(new_n579_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n578_), .A2(new_n581_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(new_n579_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n593_), .A2(new_n803_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n541_), .A2(KEYINPUT115), .A3(KEYINPUT55), .A4(new_n542_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n608_), .A2(new_n493_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT12), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n545_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n494_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n613_), .A2(new_n809_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n808_), .A2(new_n810_), .A3(KEYINPUT55), .A4(new_n542_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  XOR2_X1   g612(.A(KEYINPUT114), .B(KEYINPUT55), .Z(new_n814_));
  NAND2_X1  g613(.A1(new_n808_), .A2(new_n810_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n814_), .B1(new_n815_), .B2(new_n544_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n544_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n805_), .B(new_n813_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n818_), .A2(KEYINPUT56), .A3(new_n552_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT56), .B1(new_n818_), .B2(new_n552_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n555_), .B(new_n804_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT58), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  AOI22_X1  g622(.A1(new_n821_), .A2(new_n822_), .B1(new_n633_), .B2(new_n635_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n594_), .B(new_n555_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n556_), .A2(new_n558_), .A3(new_n804_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n632_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  AOI22_X1  g626(.A1(new_n823_), .A2(new_n824_), .B1(new_n827_), .B2(KEYINPUT57), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(KEYINPUT57), .B2(new_n827_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n648_), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n563_), .A2(KEYINPUT113), .A3(new_n752_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT113), .B1(new_n563_), .B2(new_n752_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n701_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT54), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n835_), .B(new_n701_), .C1(new_n831_), .C2(new_n832_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n830_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT59), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n652_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n840_));
  XOR2_X1   g639(.A(new_n840_), .B(KEYINPUT118), .Z(new_n841_));
  NAND3_X1  g640(.A1(new_n838_), .A2(new_n839_), .A3(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n841_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n827_), .A2(KEYINPUT116), .A3(KEYINPUT57), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT116), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n594_), .A2(new_n555_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n820_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n818_), .A2(KEYINPUT56), .A3(new_n552_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n846_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n826_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n688_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n845_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n828_), .B1(new_n844_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n828_), .B(KEYINPUT117), .C1(new_n844_), .C2(new_n853_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n856_), .A2(new_n648_), .A3(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n843_), .B1(new_n858_), .B2(new_n837_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n842_), .B1(new_n859_), .B2(new_n839_), .ZN(new_n860_));
  OAI21_X1  g659(.A(G113gat), .B1(new_n860_), .B2(new_n595_), .ZN(new_n861_));
  INV_X1    g660(.A(G113gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n859_), .A2(new_n862_), .A3(new_n594_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n863_), .ZN(G1340gat));
  XOR2_X1   g663(.A(KEYINPUT119), .B(G120gat), .Z(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n866_), .B1(new_n860_), .B2(new_n563_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n865_), .B1(new_n563_), .B2(KEYINPUT60), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n859_), .B(new_n868_), .C1(KEYINPUT60), .C2(new_n865_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n867_), .A2(new_n869_), .ZN(G1341gat));
  AND2_X1   g669(.A1(new_n689_), .A2(G127gat), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n842_), .B(new_n871_), .C1(new_n859_), .C2(new_n839_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n837_), .A2(new_n648_), .A3(new_n843_), .ZN(new_n873_));
  OR3_X1    g672(.A1(new_n873_), .A2(KEYINPUT120), .A3(G127gat), .ZN(new_n874_));
  OAI21_X1  g673(.A(KEYINPUT120), .B1(new_n873_), .B2(G127gat), .ZN(new_n875_));
  AND3_X1   g674(.A1(new_n872_), .A2(new_n874_), .A3(new_n875_), .ZN(G1342gat));
  NAND2_X1  g675(.A1(new_n636_), .A2(G134gat), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(KEYINPUT121), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n842_), .B(new_n878_), .C1(new_n859_), .C2(new_n839_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(G134gat), .B1(new_n859_), .B2(new_n632_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1343gat));
  NAND2_X1  g681(.A1(new_n858_), .A2(new_n837_), .ZN(new_n883_));
  NOR4_X1   g682(.A1(new_n759_), .A2(new_n255_), .A3(new_n682_), .A4(new_n665_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n883_), .A2(new_n594_), .A3(new_n884_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G141gat), .ZN(G1344gat));
  XNOR2_X1  g685(.A(KEYINPUT122), .B(G148gat), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n883_), .A2(new_n884_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n888_), .B2(new_n564_), .ZN(new_n889_));
  AND4_X1   g688(.A1(new_n564_), .A2(new_n883_), .A3(new_n884_), .A4(new_n887_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1345gat));
  NAND3_X1  g690(.A1(new_n883_), .A2(new_n689_), .A3(new_n884_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(KEYINPUT61), .B(G155gat), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n892_), .B(new_n893_), .ZN(G1346gat));
  NAND2_X1  g693(.A1(new_n888_), .A2(new_n632_), .ZN(new_n895_));
  INV_X1    g694(.A(G162gat), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n701_), .A2(new_n896_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(KEYINPUT123), .ZN(new_n898_));
  AOI22_X1  g697(.A1(new_n895_), .A2(new_n896_), .B1(new_n888_), .B2(new_n898_), .ZN(G1347gat));
  NOR3_X1   g698(.A1(new_n652_), .A2(new_n256_), .A3(new_n479_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  AOI211_X1 g700(.A(new_n445_), .B(new_n901_), .C1(new_n830_), .C2(new_n837_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n594_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(G169gat), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT62), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n903_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n902_), .A2(new_n226_), .A3(new_n594_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n906_), .A2(new_n907_), .A3(new_n908_), .ZN(G1348gat));
  AOI21_X1  g708(.A(G176gat), .B1(new_n902_), .B2(new_n564_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n445_), .B1(new_n858_), .B2(new_n837_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n901_), .A2(new_n222_), .A3(new_n563_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n910_), .B1(new_n911_), .B2(new_n912_), .ZN(G1349gat));
  NOR2_X1   g712(.A1(new_n901_), .A2(new_n648_), .ZN(new_n914_));
  AOI21_X1  g713(.A(G183gat), .B1(new_n911_), .B2(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n445_), .B1(new_n830_), .B2(new_n837_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n914_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n917_), .A2(new_n361_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n916_), .A2(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  OAI21_X1  g719(.A(KEYINPUT124), .B1(new_n915_), .B2(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT124), .ZN(new_n922_));
  AOI211_X1 g721(.A(new_n445_), .B(new_n917_), .C1(new_n858_), .C2(new_n837_), .ZN(new_n923_));
  OAI211_X1 g722(.A(new_n919_), .B(new_n922_), .C1(new_n923_), .C2(G183gat), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n921_), .A2(new_n924_), .ZN(G1350gat));
  INV_X1    g724(.A(KEYINPUT125), .ZN(new_n926_));
  INV_X1    g725(.A(G190gat), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n927_), .B1(new_n902_), .B2(new_n636_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n916_), .A2(new_n900_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n632_), .A2(new_n214_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n929_), .A2(new_n930_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n926_), .B1(new_n928_), .B2(new_n931_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n916_), .A2(new_n636_), .A3(new_n900_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(G190gat), .ZN(new_n934_));
  OAI211_X1 g733(.A(new_n934_), .B(KEYINPUT125), .C1(new_n929_), .C2(new_n930_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n932_), .A2(new_n935_), .ZN(G1351gat));
  NOR2_X1   g735(.A1(new_n682_), .A2(new_n693_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n937_), .A2(new_n256_), .A3(new_n665_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n938_), .B1(new_n858_), .B2(new_n837_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n939_), .A2(G197gat), .A3(new_n594_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(KEYINPUT126), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT126), .ZN(new_n942_));
  NAND4_X1  g741(.A1(new_n939_), .A2(new_n942_), .A3(G197gat), .A4(new_n594_), .ZN(new_n943_));
  INV_X1    g742(.A(new_n938_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n883_), .A2(new_n944_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n329_), .B1(new_n945_), .B2(new_n659_), .ZN(new_n946_));
  AND3_X1   g745(.A1(new_n941_), .A2(new_n943_), .A3(new_n946_), .ZN(G1352gat));
  AOI21_X1  g746(.A(G204gat), .B1(new_n939_), .B2(new_n564_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n945_), .A2(new_n563_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n948_), .B1(new_n949_), .B2(new_n351_), .ZN(G1353gat));
  NOR3_X1   g749(.A1(KEYINPUT127), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n951_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n939_), .A2(new_n689_), .A3(new_n952_), .ZN(new_n953_));
  OAI21_X1  g752(.A(KEYINPUT127), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n954_));
  INV_X1    g753(.A(new_n954_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n953_), .B(new_n955_), .ZN(G1354gat));
  OAI21_X1  g755(.A(G218gat), .B1(new_n945_), .B2(new_n701_), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n939_), .A2(new_n335_), .A3(new_n632_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n957_), .A2(new_n958_), .ZN(G1355gat));
endmodule


