//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n604_, new_n605_,
    new_n606_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n835_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n868_, new_n869_, new_n870_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT0), .B(G57gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  XOR2_X1   g004(.A(G141gat), .B(G148gat), .Z(new_n206_));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT1), .ZN(new_n208_));
  OR2_X1    g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n207_), .A2(KEYINPUT1), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n206_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT85), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n209_), .A2(new_n207_), .ZN(new_n214_));
  XOR2_X1   g013(.A(new_n214_), .B(KEYINPUT86), .Z(new_n215_));
  OR3_X1    g014(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT2), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n216_), .A2(new_n219_), .A3(new_n220_), .A4(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n215_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n213_), .A2(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(G127gat), .B(G134gat), .Z(new_n225_));
  XNOR2_X1  g024(.A(G113gat), .B(G120gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n225_), .B(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n224_), .B(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT4), .ZN(new_n229_));
  OR3_X1    g028(.A1(new_n228_), .A2(KEYINPUT93), .A3(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n224_), .A2(new_n229_), .A3(new_n227_), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT93), .B1(new_n228_), .B2(new_n229_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G225gat), .A2(G233gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT94), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n228_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n237_), .A2(new_n235_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n205_), .B1(new_n236_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT33), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(KEYINPUT95), .A3(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n238_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n205_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n240_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT95), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  OAI211_X1 g045(.A(KEYINPUT33), .B(new_n205_), .C1(new_n236_), .C2(new_n238_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT80), .B(KEYINPUT23), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G183gat), .A2(G190gat), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  MUX2_X1   g049(.A(KEYINPUT23), .B(new_n248_), .S(new_n250_), .Z(new_n251_));
  OAI21_X1  g050(.A(new_n251_), .B1(G183gat), .B2(G190gat), .ZN(new_n252_));
  NOR2_X1   g051(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(G169gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT25), .B(G183gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT26), .B(G190gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT24), .ZN(new_n258_));
  NOR2_X1   g057(.A1(G169gat), .A2(G176gat), .ZN(new_n259_));
  AOI22_X1  g058(.A1(new_n256_), .A2(new_n257_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  AND2_X1   g059(.A1(G169gat), .A2(G176gat), .ZN(new_n261_));
  OR3_X1    g060(.A1(new_n261_), .A2(new_n259_), .A3(new_n258_), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  OR3_X1    g062(.A1(new_n249_), .A2(KEYINPUT81), .A3(KEYINPUT23), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT81), .B1(new_n249_), .B2(KEYINPUT23), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n264_), .B(new_n265_), .C1(new_n250_), .C2(new_n248_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n263_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n255_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G197gat), .B(G204gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT88), .B(KEYINPUT21), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  OR2_X1    g070(.A1(new_n271_), .A2(KEYINPUT89), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(KEYINPUT89), .ZN(new_n273_));
  INV_X1    g072(.A(new_n269_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT21), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G211gat), .B(G218gat), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n272_), .A2(new_n273_), .A3(new_n275_), .A4(new_n276_), .ZN(new_n277_));
  OR2_X1    g076(.A1(new_n275_), .A2(new_n276_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n268_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT20), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n277_), .A2(new_n278_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n266_), .B1(G183gat), .B2(G190gat), .ZN(new_n284_));
  AOI22_X1  g083(.A1(new_n284_), .A2(new_n254_), .B1(new_n263_), .B2(new_n251_), .ZN(new_n285_));
  OR3_X1    g084(.A1(new_n283_), .A2(KEYINPUT91), .A3(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT91), .B1(new_n283_), .B2(new_n285_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n282_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G226gat), .A2(G233gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT19), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n283_), .A2(new_n285_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n268_), .A2(new_n279_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n292_), .A2(new_n293_), .A3(KEYINPUT20), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n294_), .A2(new_n290_), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n291_), .A2(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(G8gat), .B(G36gat), .Z(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G64gat), .B(G92gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n296_), .A2(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n205_), .B1(new_n237_), .B2(new_n235_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n303_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n291_), .A2(new_n295_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n301_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n302_), .A2(new_n304_), .A3(new_n307_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n241_), .A2(new_n246_), .A3(new_n247_), .A4(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n242_), .A2(new_n243_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n239_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n294_), .A2(new_n290_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n312_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(KEYINPUT32), .A3(new_n301_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT32), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n296_), .B1(new_n315_), .B2(new_n306_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n311_), .A2(new_n314_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n309_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G78gat), .B(G106gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G22gat), .B(G50gat), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n319_), .B(new_n320_), .Z(new_n321_));
  OR2_X1    g120(.A1(new_n224_), .A2(KEYINPUT29), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n322_), .B(KEYINPUT28), .Z(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(KEYINPUT87), .B1(new_n224_), .B2(KEYINPUT29), .ZN(new_n325_));
  AND2_X1   g124(.A1(G228gat), .A2(G233gat), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT90), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n224_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n325_), .A2(new_n326_), .A3(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n224_), .A2(new_n327_), .A3(KEYINPUT29), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n283_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n326_), .B1(new_n325_), .B2(new_n279_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n324_), .A2(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n323_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n321_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n334_), .A2(new_n335_), .A3(new_n321_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(KEYINPUT82), .B(G15gat), .Z(new_n341_));
  NAND2_X1  g140(.A1(G227gat), .A2(G233gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n268_), .B(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G71gat), .B(G99gat), .ZN(new_n345_));
  INV_X1    g144(.A(G43gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT30), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n344_), .B(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT84), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n227_), .B(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n352_), .A2(new_n354_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n350_), .A2(new_n351_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n355_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n340_), .A2(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n305_), .A2(new_n306_), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n361_), .A2(KEYINPUT97), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(KEYINPUT97), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT27), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n301_), .B(KEYINPUT96), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n364_), .B1(new_n313_), .B2(new_n365_), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n362_), .A2(new_n363_), .A3(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n302_), .A2(new_n307_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(new_n364_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT98), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT98), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n368_), .A2(new_n371_), .A3(new_n364_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n367_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n338_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n359_), .B1(new_n374_), .B2(new_n336_), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n352_), .A2(new_n354_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n352_), .A2(new_n354_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n376_), .B1(new_n357_), .B2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n378_), .A2(new_n338_), .A3(new_n337_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n311_), .B1(new_n375_), .B2(new_n379_), .ZN(new_n380_));
  AOI22_X1  g179(.A1(new_n318_), .A2(new_n360_), .B1(new_n373_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G232gat), .A2(G233gat), .ZN(new_n382_));
  XOR2_X1   g181(.A(new_n382_), .B(KEYINPUT34), .Z(new_n383_));
  XOR2_X1   g182(.A(KEYINPUT73), .B(KEYINPUT35), .Z(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT64), .ZN(new_n386_));
  OR2_X1    g185(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n387_));
  INV_X1    g186(.A(G106gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n387_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(G85gat), .ZN(new_n391_));
  INV_X1    g190(.A(G92gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G85gat), .A2(G92gat), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n393_), .A2(KEYINPUT9), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n390_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G99gat), .A2(G106gat), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT6), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT9), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(G85gat), .A3(G92gat), .ZN(new_n401_));
  NAND3_X1  g200(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n399_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n386_), .B1(new_n396_), .B2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n403_), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n405_), .A2(KEYINPUT64), .A3(new_n390_), .A4(new_n395_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n397_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT67), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n410_), .A2(KEYINPUT6), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n398_), .A2(KEYINPUT67), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n409_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n398_), .A2(KEYINPUT67), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(KEYINPUT6), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n415_), .A3(new_n397_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n413_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT65), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT7), .ZN(new_n419_));
  INV_X1    g218(.A(G99gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n388_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n418_), .B(new_n419_), .C1(new_n421_), .C2(KEYINPUT66), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n420_), .A2(new_n388_), .A3(KEYINPUT65), .ZN(new_n423_));
  NOR3_X1   g222(.A1(KEYINPUT66), .A2(G99gat), .A3(G106gat), .ZN(new_n424_));
  OAI211_X1 g223(.A(KEYINPUT7), .B(new_n423_), .C1(new_n424_), .C2(KEYINPUT65), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n417_), .B1(new_n422_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n393_), .A2(new_n394_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT8), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n399_), .A2(new_n402_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n429_), .B1(new_n425_), .B2(new_n422_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n427_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT8), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n430_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n408_), .B1(new_n428_), .B2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G29gat), .B(G36gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G43gat), .B(G50gat), .ZN(new_n438_));
  XOR2_X1   g237(.A(new_n437_), .B(new_n438_), .Z(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n437_), .B(new_n438_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n440_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n436_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n383_), .A2(new_n384_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n425_), .A2(new_n422_), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n414_), .A2(new_n415_), .A3(new_n397_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n397_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n449_), .A2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n432_), .B1(new_n453_), .B2(new_n431_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n407_), .B1(new_n454_), .B2(new_n434_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n442_), .A2(KEYINPUT15), .A3(new_n444_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT15), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n439_), .A2(new_n441_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n443_), .A2(new_n440_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n457_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n455_), .A2(new_n456_), .A3(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n385_), .B1(new_n448_), .B2(new_n461_), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n460_), .A2(new_n456_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n455_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n385_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n464_), .A2(new_n465_), .A3(new_n447_), .A4(new_n446_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G190gat), .B(G218gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G134gat), .B(G162gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n469_), .A2(KEYINPUT36), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n462_), .A2(new_n466_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(new_n469_), .B(KEYINPUT36), .Z(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n462_), .A2(new_n466_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT76), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n474_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n462_), .A2(new_n466_), .A3(KEYINPUT76), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n472_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G127gat), .B(G155gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT16), .ZN(new_n481_));
  XOR2_X1   g280(.A(G183gat), .B(G211gat), .Z(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT68), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G57gat), .B(G64gat), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n484_), .B1(new_n485_), .B2(KEYINPUT11), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n485_), .A2(KEYINPUT11), .ZN(new_n488_));
  XOR2_X1   g287(.A(G71gat), .B(G78gat), .Z(new_n489_));
  NAND3_X1  g288(.A1(new_n485_), .A2(new_n484_), .A3(KEYINPUT11), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .A4(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n489_), .B1(KEYINPUT11), .B2(new_n485_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n490_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n492_), .B1(new_n493_), .B2(new_n486_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n491_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G15gat), .B(G22gat), .ZN(new_n497_));
  INV_X1    g296(.A(G1gat), .ZN(new_n498_));
  INV_X1    g297(.A(G8gat), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT14), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G1gat), .B(G8gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n496_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n503_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n495_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(G231gat), .ZN(new_n508_));
  INV_X1    g307(.A(G233gat), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n507_), .B(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n483_), .B1(new_n512_), .B2(KEYINPUT77), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n483_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n513_), .B1(KEYINPUT17), .B2(new_n514_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n513_), .A2(KEYINPUT17), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NOR3_X1   g316(.A1(new_n381_), .A2(new_n479_), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT12), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n519_), .B1(new_n436_), .B2(new_n495_), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n407_), .B(new_n495_), .C1(new_n454_), .C2(new_n434_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G230gat), .A2(G233gat), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n455_), .A2(new_n496_), .A3(KEYINPUT12), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n520_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT69), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n436_), .A2(new_n495_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n521_), .ZN(new_n529_));
  OAI211_X1 g328(.A(G230gat), .B(G233gat), .C1(new_n528_), .C2(new_n529_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n520_), .A2(new_n523_), .A3(KEYINPUT69), .A4(new_n524_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n527_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  XOR2_X1   g331(.A(G120gat), .B(G148gat), .Z(new_n533_));
  XNOR2_X1  g332(.A(G176gat), .B(G204gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n535_), .B(new_n536_), .Z(new_n537_));
  NAND2_X1  g336(.A1(new_n532_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT71), .ZN(new_n539_));
  INV_X1    g338(.A(new_n537_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n527_), .A2(new_n530_), .A3(new_n531_), .A4(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n538_), .A2(new_n539_), .A3(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n532_), .A2(KEYINPUT71), .A3(new_n537_), .ZN(new_n543_));
  AOI21_X1  g342(.A(KEYINPUT13), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n542_), .A2(KEYINPUT13), .A3(new_n543_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT72), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n545_), .A2(KEYINPUT72), .A3(new_n546_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n463_), .A2(new_n503_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n445_), .A2(new_n505_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G229gat), .A2(G233gat), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n445_), .B(new_n503_), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n556_), .A2(new_n554_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G113gat), .B(G141gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G169gat), .B(G197gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n559_), .B(new_n560_), .Z(new_n561_));
  INV_X1    g360(.A(KEYINPUT79), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n558_), .B(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n551_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n518_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n311_), .ZN(new_n568_));
  OAI21_X1  g367(.A(G1gat), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n570_));
  NOR3_X1   g369(.A1(new_n381_), .A2(new_n551_), .A3(new_n565_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n475_), .A2(new_n473_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n572_), .A2(KEYINPUT37), .A3(new_n471_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n477_), .A2(new_n478_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(new_n471_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT37), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n574_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n517_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT78), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n571_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n583_), .A2(new_n498_), .A3(new_n311_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(new_n570_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n585_), .A2(KEYINPUT100), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n585_), .A2(KEYINPUT100), .ZN(new_n587_));
  OAI221_X1 g386(.A(new_n569_), .B1(new_n570_), .B2(new_n584_), .C1(new_n586_), .C2(new_n587_), .ZN(G1324gat));
  OAI21_X1  g387(.A(G8gat), .B1(new_n567_), .B2(new_n373_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT39), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT101), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n370_), .A2(new_n372_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n367_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(new_n499_), .ZN(new_n596_));
  OR3_X1    g395(.A1(new_n582_), .A2(new_n592_), .A3(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n592_), .B1(new_n582_), .B2(new_n596_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n589_), .A2(new_n590_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n591_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT40), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(G1325gat));
  OAI21_X1  g402(.A(G15gat), .B1(new_n567_), .B2(new_n378_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT41), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n582_), .A2(G15gat), .A3(new_n378_), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n605_), .A2(new_n606_), .ZN(G1326gat));
  OR3_X1    g406(.A1(new_n582_), .A2(G22gat), .A3(new_n339_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n518_), .A2(new_n566_), .A3(new_n340_), .ZN(new_n609_));
  XOR2_X1   g408(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n610_));
  AND3_X1   g409(.A1(new_n609_), .A2(G22gat), .A3(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n610_), .B1(new_n609_), .B2(G22gat), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n608_), .B1(new_n611_), .B2(new_n612_), .ZN(G1327gat));
  INV_X1    g412(.A(KEYINPUT44), .ZN(new_n614_));
  OAI21_X1  g413(.A(KEYINPUT43), .B1(new_n381_), .B2(new_n578_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n318_), .A2(new_n360_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n373_), .A2(new_n380_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT43), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n573_), .B1(new_n479_), .B2(KEYINPUT37), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n618_), .A2(new_n619_), .A3(new_n620_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n615_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n566_), .A2(new_n517_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n614_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n615_), .A2(new_n621_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n625_), .A2(KEYINPUT44), .A3(new_n517_), .A4(new_n566_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(G29gat), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n627_), .A2(new_n628_), .A3(new_n568_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n579_), .A2(new_n576_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n571_), .A2(new_n311_), .A3(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n629_), .B1(new_n628_), .B2(new_n631_), .ZN(G1328gat));
  NAND3_X1  g431(.A1(new_n624_), .A2(new_n595_), .A3(new_n626_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(G36gat), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n571_), .A2(new_n630_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n373_), .A2(G36gat), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT45), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n634_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT46), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n634_), .A2(KEYINPUT46), .A3(new_n639_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(G1329gat));
  OAI21_X1  g443(.A(new_n346_), .B1(new_n635_), .B2(new_n378_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n359_), .A2(G43gat), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n645_), .B1(new_n627_), .B2(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g447(.A(G50gat), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n627_), .A2(new_n649_), .A3(new_n339_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n571_), .A2(new_n340_), .A3(new_n630_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n649_), .B2(new_n651_), .ZN(G1331gat));
  INV_X1    g451(.A(KEYINPUT104), .ZN(new_n653_));
  OR3_X1    g452(.A1(new_n381_), .A2(KEYINPUT103), .A3(new_n564_), .ZN(new_n654_));
  OAI21_X1  g453(.A(KEYINPUT103), .B1(new_n381_), .B2(new_n564_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n551_), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n581_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n653_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n655_), .A2(new_n551_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n659_), .A2(KEYINPUT104), .A3(new_n581_), .A4(new_n654_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n568_), .A2(G57gat), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n658_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n565_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n618_), .A2(new_n576_), .A3(new_n551_), .A4(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G57gat), .B1(new_n665_), .B2(new_n568_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n662_), .A2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT105), .ZN(G1332gat));
  OAI21_X1  g467(.A(G64gat), .B1(new_n665_), .B2(new_n373_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT48), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n658_), .A2(new_n660_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n373_), .A2(G64gat), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT106), .Z(new_n673_));
  OAI21_X1  g472(.A(new_n670_), .B1(new_n671_), .B2(new_n673_), .ZN(G1333gat));
  INV_X1    g473(.A(G71gat), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n658_), .A2(new_n660_), .A3(new_n675_), .A4(new_n359_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G71gat), .B1(new_n665_), .B2(new_n378_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT49), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n679_), .B(new_n680_), .ZN(G1334gat));
  OAI21_X1  g480(.A(G78gat), .B1(new_n665_), .B2(new_n339_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT50), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n339_), .A2(G78gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n683_), .B1(new_n671_), .B2(new_n684_), .ZN(G1335gat));
  INV_X1    g484(.A(new_n551_), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n686_), .A2(new_n579_), .A3(new_n564_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n625_), .A2(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(G85gat), .B1(new_n688_), .B2(new_n568_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n656_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(new_n630_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n311_), .A2(new_n391_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n689_), .B1(new_n691_), .B2(new_n692_), .ZN(G1336gat));
  OAI21_X1  g492(.A(G92gat), .B1(new_n688_), .B2(new_n373_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n595_), .A2(new_n392_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n694_), .B1(new_n691_), .B2(new_n695_), .ZN(G1337gat));
  NOR2_X1   g495(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n387_), .A2(new_n389_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n690_), .A2(new_n698_), .A3(new_n359_), .A4(new_n630_), .ZN(new_n699_));
  OAI21_X1  g498(.A(G99gat), .B1(new_n688_), .B2(new_n378_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n697_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  AND2_X1   g500(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n701_), .B(new_n702_), .ZN(G1338gat));
  NAND3_X1  g502(.A1(new_n625_), .A2(new_n340_), .A3(new_n687_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(KEYINPUT109), .B(KEYINPUT52), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n704_), .A2(G106gat), .A3(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n704_), .B2(G106gat), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n340_), .A2(new_n388_), .ZN(new_n708_));
  OAI22_X1  g507(.A1(new_n706_), .A2(new_n707_), .B1(new_n691_), .B2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g509(.A(KEYINPUT115), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT54), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n547_), .A2(new_n578_), .A3(new_n664_), .A4(new_n713_), .ZN(new_n714_));
  AOI211_X1 g513(.A(new_n663_), .B(new_n620_), .C1(new_n545_), .C2(new_n546_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(KEYINPUT110), .B(KEYINPUT54), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n714_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n576_), .A2(KEYINPUT57), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n564_), .A2(new_n541_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n520_), .A2(new_n523_), .A3(KEYINPUT55), .A4(new_n524_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT111), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n427_), .B1(new_n449_), .B2(new_n452_), .ZN(new_n724_));
  OAI22_X1  g523(.A1(new_n724_), .A2(new_n432_), .B1(new_n430_), .B2(new_n433_), .ZN(new_n725_));
  AOI211_X1 g524(.A(new_n519_), .B(new_n495_), .C1(new_n725_), .C2(new_n407_), .ZN(new_n726_));
  AOI21_X1  g525(.A(KEYINPUT12), .B1(new_n455_), .B2(new_n496_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT111), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n728_), .A2(new_n729_), .A3(KEYINPUT55), .A4(new_n523_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n723_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT55), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n527_), .A2(new_n732_), .A3(new_n531_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n728_), .A2(new_n521_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(G230gat), .A3(G233gat), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n731_), .A2(new_n733_), .A3(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(new_n537_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT56), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n736_), .A2(KEYINPUT56), .A3(new_n537_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n721_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n554_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n552_), .A2(new_n553_), .A3(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n743_), .B1(new_n556_), .B2(new_n742_), .ZN(new_n744_));
  MUX2_X1   g543(.A(new_n744_), .B(new_n558_), .S(new_n561_), .Z(new_n745_));
  NAND3_X1  g544(.A1(new_n542_), .A2(new_n543_), .A3(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n720_), .B1(new_n741_), .B2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT112), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n564_), .A2(new_n541_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n736_), .A2(KEYINPUT56), .A3(new_n537_), .ZN(new_n751_));
  AOI21_X1  g550(.A(KEYINPUT56), .B1(new_n736_), .B2(new_n537_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n750_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(new_n746_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT112), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n754_), .A2(new_n755_), .A3(new_n720_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n749_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n745_), .A2(new_n541_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n620_), .B1(new_n759_), .B2(KEYINPUT58), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n745_), .A2(new_n541_), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n761_), .B(KEYINPUT58), .C1(new_n751_), .C2(new_n752_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n479_), .B1(new_n753_), .B2(new_n746_), .ZN(new_n764_));
  OAI22_X1  g563(.A1(new_n760_), .A2(new_n763_), .B1(new_n764_), .B2(KEYINPUT57), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n517_), .B1(new_n757_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT114), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n576_), .B1(new_n741_), .B2(new_n747_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT57), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n761_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT58), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n773_), .A2(new_n620_), .A3(new_n762_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n770_), .A2(new_n749_), .A3(new_n774_), .A4(new_n756_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT114), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n776_), .A3(new_n517_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n718_), .B1(new_n767_), .B2(new_n777_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n595_), .A2(new_n568_), .A3(new_n375_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT59), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n711_), .B1(new_n778_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT113), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n755_), .B1(new_n754_), .B2(new_n720_), .ZN(new_n784_));
  AOI211_X1 g583(.A(KEYINPUT112), .B(new_n719_), .C1(new_n753_), .C2(new_n746_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n578_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n787_));
  AOI22_X1  g586(.A1(new_n769_), .A2(new_n768_), .B1(new_n787_), .B2(new_n762_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n579_), .B1(new_n786_), .B2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n783_), .B1(new_n789_), .B2(new_n718_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n766_), .A2(KEYINPUT113), .A3(new_n717_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n790_), .A2(new_n791_), .A3(new_n779_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT59), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n775_), .A2(new_n776_), .A3(new_n517_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n776_), .B1(new_n775_), .B2(new_n517_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n717_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n781_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(KEYINPUT115), .A3(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(G113gat), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n565_), .A2(new_n799_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n782_), .A2(new_n793_), .A3(new_n798_), .A4(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n799_), .B1(new_n792_), .B2(new_n565_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT116), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n801_), .A2(KEYINPUT116), .A3(new_n802_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(G1340gat));
  AND2_X1   g606(.A1(new_n790_), .A2(new_n791_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n686_), .A2(KEYINPUT60), .ZN(new_n809_));
  MUX2_X1   g608(.A(new_n809_), .B(KEYINPUT60), .S(G120gat), .Z(new_n810_));
  NAND3_X1  g609(.A1(new_n808_), .A2(new_n779_), .A3(new_n810_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(KEYINPUT117), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n782_), .A2(new_n793_), .A3(new_n798_), .ZN(new_n813_));
  OAI21_X1  g612(.A(G120gat), .B1(new_n813_), .B2(new_n686_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(G1341gat));
  INV_X1    g614(.A(G127gat), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n517_), .A2(new_n816_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n782_), .A2(new_n793_), .A3(new_n798_), .A4(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n816_), .B1(new_n792_), .B2(new_n517_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT118), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT118), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n818_), .A2(new_n822_), .A3(new_n819_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(G1342gat));
  XNOR2_X1  g623(.A(KEYINPUT119), .B(G134gat), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n813_), .A2(new_n578_), .A3(new_n825_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n792_), .A2(new_n576_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n827_), .A2(G134gat), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n826_), .A2(new_n828_), .ZN(G1343gat));
  NOR3_X1   g628(.A1(new_n595_), .A2(new_n568_), .A3(new_n379_), .ZN(new_n830_));
  XOR2_X1   g629(.A(new_n830_), .B(KEYINPUT120), .Z(new_n831_));
  AND2_X1   g630(.A1(new_n808_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(new_n564_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n551_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(new_n835_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g635(.A1(new_n832_), .A2(new_n579_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(KEYINPUT61), .B(G155gat), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n837_), .B(new_n838_), .ZN(G1346gat));
  INV_X1    g638(.A(G162gat), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n832_), .A2(new_n840_), .A3(new_n479_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n832_), .A2(new_n620_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n842_), .B2(new_n840_), .ZN(G1347gat));
  NOR2_X1   g642(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n844_));
  AND2_X1   g643(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n595_), .A2(new_n568_), .A3(new_n359_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(KEYINPUT121), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n847_), .A2(new_n340_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n796_), .A2(KEYINPUT123), .A3(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT123), .B1(new_n796_), .B2(new_n848_), .ZN(new_n850_));
  OAI221_X1 g649(.A(new_n564_), .B1(new_n844_), .B2(new_n845_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n796_), .A2(new_n564_), .A3(new_n848_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(KEYINPUT122), .B(KEYINPUT62), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n852_), .A2(G169gat), .A3(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n853_), .B1(new_n852_), .B2(G169gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n851_), .B1(new_n854_), .B2(new_n855_), .ZN(G1348gat));
  OAI21_X1  g655(.A(new_n551_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n857_));
  INV_X1    g656(.A(G176gat), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n808_), .A2(new_n848_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n686_), .A2(new_n858_), .ZN(new_n860_));
  AOI22_X1  g659(.A1(new_n857_), .A2(new_n858_), .B1(new_n859_), .B2(new_n860_), .ZN(G1349gat));
  AOI21_X1  g660(.A(G183gat), .B1(new_n859_), .B2(new_n579_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n849_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n850_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n517_), .A2(new_n256_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n862_), .B1(new_n865_), .B2(new_n866_), .ZN(G1350gat));
  OAI211_X1 g666(.A(new_n479_), .B(new_n257_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n578_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n869_));
  INV_X1    g668(.A(G190gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n868_), .B1(new_n869_), .B2(new_n870_), .ZN(G1351gat));
  NOR3_X1   g670(.A1(new_n373_), .A2(new_n311_), .A3(new_n379_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n808_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n564_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n551_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(G204gat), .ZN(G1353gat));
  NOR3_X1   g677(.A1(KEYINPUT125), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n879_));
  OAI21_X1  g678(.A(KEYINPUT125), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n879_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n517_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n883_));
  XOR2_X1   g682(.A(new_n883_), .B(KEYINPUT124), .Z(new_n884_));
  NAND3_X1  g683(.A1(new_n808_), .A2(new_n872_), .A3(new_n884_), .ZN(new_n885_));
  MUX2_X1   g684(.A(new_n879_), .B(new_n882_), .S(new_n885_), .Z(G1354gat));
  XNOR2_X1  g685(.A(KEYINPUT127), .B(G218gat), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n873_), .A2(new_n578_), .A3(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n808_), .A2(new_n479_), .A3(new_n872_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT126), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n889_), .B(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n888_), .B1(new_n891_), .B2(new_n887_), .ZN(G1355gat));
endmodule


