//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1 0 0 1 0 0 0 1 0 1 1 0 1 0 1 1 1 1 0 0 0 1 1 1 1 0 0 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n607_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n720_, new_n721_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n840_, new_n842_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n875_, new_n876_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_;
  XOR2_X1   g000(.A(G78gat), .B(G106gat), .Z(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G141gat), .A2(G148gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT2), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n206_), .A2(new_n209_), .A3(new_n210_), .A4(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n212_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n204_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(new_n207_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n213_), .B1(KEYINPUT1), .B2(new_n215_), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n215_), .A2(KEYINPUT1), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n219_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT82), .B1(new_n217_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n222_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT82), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n212_), .A2(new_n216_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n223_), .A2(new_n227_), .A3(KEYINPUT29), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n228_), .B(KEYINPUT83), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G228gat), .A2(G233gat), .ZN(new_n230_));
  INV_X1    g029(.A(G197gat), .ZN(new_n231_));
  INV_X1    g030(.A(G204gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G197gat), .A2(G204gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(KEYINPUT21), .A3(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G211gat), .B(G218gat), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT21), .ZN(new_n238_));
  INV_X1    g037(.A(new_n234_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(G197gat), .A2(G204gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n238_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n241_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n237_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n229_), .A2(new_n230_), .A3(new_n243_), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n237_), .A2(new_n242_), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT29), .B1(new_n217_), .B2(new_n222_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n245_), .B1(new_n246_), .B2(KEYINPUT84), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n247_), .B1(KEYINPUT84), .B2(new_n246_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n248_), .A2(G228gat), .A3(G233gat), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n203_), .B1(new_n244_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G22gat), .B(G50gat), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n223_), .A2(new_n227_), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT28), .B1(new_n253_), .B2(KEYINPUT29), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NOR3_X1   g054(.A1(new_n253_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n252_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n256_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n252_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n258_), .A2(new_n254_), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n244_), .A2(new_n203_), .A3(new_n249_), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n251_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n262_), .B1(new_n251_), .B2(new_n263_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(G127gat), .B(G134gat), .Z(new_n267_));
  XOR2_X1   g066(.A(G113gat), .B(G120gat), .Z(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n223_), .A2(new_n227_), .A3(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n269_), .A2(new_n224_), .A3(new_n226_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(new_n272_), .A3(KEYINPUT4), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G225gat), .A2(G233gat), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n223_), .A2(new_n227_), .A3(new_n270_), .A4(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n273_), .A2(new_n275_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT90), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n271_), .A2(new_n272_), .A3(new_n274_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT93), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT93), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n271_), .A2(new_n272_), .A3(new_n283_), .A4(new_n274_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n273_), .A2(KEYINPUT90), .A3(new_n275_), .A4(new_n277_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n280_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G1gat), .B(G29gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT92), .ZN(new_n289_));
  XOR2_X1   g088(.A(G57gat), .B(G85gat), .Z(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT91), .B(KEYINPUT0), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n287_), .A2(new_n294_), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n280_), .A2(new_n285_), .A3(new_n293_), .A4(new_n286_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n297_), .A2(KEYINPUT96), .ZN(new_n298_));
  NAND2_X1  g097(.A1(KEYINPUT80), .A2(G169gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT22), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT22), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n301_), .A2(KEYINPUT80), .A3(G169gat), .ZN(new_n302_));
  INV_X1    g101(.A(G176gat), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n300_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G183gat), .A2(G190gat), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT23), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n308_));
  INV_X1    g107(.A(G183gat), .ZN(new_n309_));
  INV_X1    g108(.A(G190gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n307_), .A2(new_n308_), .A3(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n304_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(G169gat), .A2(G176gat), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n316_), .A2(KEYINPUT24), .A3(new_n313_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n305_), .A2(KEYINPUT23), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n306_), .A2(G183gat), .A3(G190gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT24), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n315_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n317_), .A2(new_n320_), .A3(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT25), .B(G183gat), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT26), .B1(new_n310_), .B2(KEYINPUT79), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT79), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT26), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n326_), .A2(new_n327_), .A3(G190gat), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n324_), .A2(new_n325_), .A3(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n314_), .B1(new_n323_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G227gat), .A2(G233gat), .ZN(new_n331_));
  INV_X1    g130(.A(G71gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(G99gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n330_), .B(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(new_n270_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G15gat), .B(G43gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT81), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT30), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT31), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n336_), .B(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n297_), .A2(KEYINPUT96), .ZN(new_n342_));
  AND3_X1   g141(.A1(new_n298_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT98), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G8gat), .B(G36gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT18), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G64gat), .B(G92gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT22), .B(G169gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n303_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(new_n313_), .A3(new_n312_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n321_), .A2(KEYINPUT85), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT85), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT24), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n320_), .B1(new_n357_), .B2(new_n316_), .ZN(new_n358_));
  AND2_X1   g157(.A1(G169gat), .A2(G176gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n359_), .A2(new_n315_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n327_), .A2(G190gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n309_), .A2(KEYINPUT25), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT25), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(G183gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n310_), .A2(KEYINPUT26), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n362_), .A2(new_n363_), .A3(new_n365_), .A4(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n361_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT86), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n358_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT26), .B(G190gat), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n360_), .A2(new_n357_), .B1(new_n324_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT86), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n353_), .B1(new_n370_), .B2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT87), .B1(new_n374_), .B2(new_n245_), .ZN(new_n375_));
  AND2_X1   g174(.A1(new_n354_), .A2(new_n356_), .ZN(new_n376_));
  AOI22_X1  g175(.A1(new_n376_), .A2(new_n315_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n377_), .B1(new_n372_), .B2(KEYINPUT86), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n368_), .A2(new_n369_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n352_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT87), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n380_), .A2(new_n381_), .A3(new_n243_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n330_), .A2(new_n243_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT20), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n375_), .A2(new_n382_), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT88), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT19), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n386_), .A2(new_n387_), .A3(new_n389_), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n245_), .B(new_n352_), .C1(new_n378_), .C2(new_n379_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n389_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n384_), .B1(new_n330_), .B2(new_n243_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n391_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT88), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n395_), .B1(new_n386_), .B2(new_n389_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n349_), .B1(new_n390_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT89), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT89), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n399_), .B(new_n349_), .C1(new_n390_), .C2(new_n396_), .ZN(new_n400_));
  OR3_X1    g199(.A1(new_n390_), .A2(new_n396_), .A3(new_n349_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n398_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  XOR2_X1   g201(.A(KEYINPUT97), .B(KEYINPUT27), .Z(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT27), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n391_), .A2(new_n393_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n389_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n408_), .B1(new_n386_), .B2(new_n389_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n406_), .B1(new_n409_), .B2(new_n348_), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n397_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n344_), .B1(new_n405_), .B2(new_n412_), .ZN(new_n413_));
  AOI211_X1 g212(.A(KEYINPUT98), .B(new_n411_), .C1(new_n402_), .C2(new_n404_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n266_), .B(new_n343_), .C1(new_n413_), .C2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT99), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NOR3_X1   g216(.A1(new_n390_), .A2(new_n396_), .A3(new_n349_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n418_), .B1(KEYINPUT89), .B2(new_n397_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n403_), .B1(new_n419_), .B2(new_n400_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT98), .B1(new_n420_), .B2(new_n411_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n411_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n344_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n421_), .A2(new_n423_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n424_), .A2(KEYINPUT99), .A3(new_n266_), .A4(new_n343_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n341_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n349_), .A2(KEYINPUT32), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n409_), .A2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n427_), .B(KEYINPUT94), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n429_), .B1(new_n390_), .B2(new_n396_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n297_), .A2(new_n428_), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT33), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n273_), .A2(new_n274_), .A3(new_n277_), .ZN(new_n433_));
  AND2_X1   g232(.A1(new_n271_), .A2(new_n272_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n293_), .B1(new_n434_), .B2(new_n275_), .ZN(new_n435_));
  AOI22_X1  g234(.A1(new_n296_), .A2(new_n432_), .B1(new_n433_), .B2(new_n435_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n280_), .A2(new_n286_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n437_), .A2(KEYINPUT33), .A3(new_n293_), .A4(new_n285_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n431_), .B1(new_n402_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(new_n266_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT95), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT95), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n440_), .A2(new_n266_), .A3(new_n443_), .ZN(new_n444_));
  OR2_X1    g243(.A1(new_n264_), .A2(new_n265_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n445_), .A2(new_n422_), .A3(new_n342_), .A4(new_n298_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n442_), .A2(new_n444_), .A3(new_n446_), .ZN(new_n447_));
  AOI22_X1  g246(.A1(new_n417_), .A2(new_n425_), .B1(new_n426_), .B2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G15gat), .B(G22gat), .ZN(new_n449_));
  INV_X1    g248(.A(G1gat), .ZN(new_n450_));
  INV_X1    g249(.A(G8gat), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT14), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n449_), .A2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G1gat), .B(G8gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G29gat), .B(G36gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G43gat), .B(G50gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  OR2_X1    g258(.A1(new_n455_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G229gat), .A2(G233gat), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n458_), .B(KEYINPUT15), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n455_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n455_), .B(new_n459_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n461_), .ZN(new_n466_));
  AOI22_X1  g265(.A1(new_n462_), .A2(new_n464_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G113gat), .B(G141gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G169gat), .B(G197gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n468_), .B(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT78), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n467_), .B(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(KEYINPUT10), .B(G99gat), .Z(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT64), .B(G106gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G99gat), .A2(G106gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT6), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT6), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(G99gat), .A3(G106gat), .ZN(new_n479_));
  AOI22_X1  g278(.A1(new_n474_), .A2(new_n475_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(KEYINPUT65), .B(KEYINPUT9), .Z(new_n481_));
  XNOR2_X1  g280(.A(KEYINPUT66), .B(G85gat), .ZN(new_n482_));
  XOR2_X1   g281(.A(KEYINPUT67), .B(G92gat), .Z(new_n483_));
  AOI21_X1  g282(.A(new_n481_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(G85gat), .ZN(new_n485_));
  INV_X1    g284(.A(G92gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT9), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G85gat), .A2(G92gat), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n487_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n480_), .B1(new_n484_), .B2(new_n490_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n487_), .A2(new_n489_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n477_), .A2(new_n479_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(G99gat), .A2(G106gat), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT7), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  OAI221_X1 g297(.A(new_n492_), .B1(KEYINPUT68), .B2(KEYINPUT8), .C1(new_n493_), .C2(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n492_), .B1(new_n493_), .B2(new_n498_), .ZN(new_n500_));
  AOI21_X1  g299(.A(KEYINPUT8), .B1(new_n492_), .B2(KEYINPUT68), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n491_), .A2(new_n499_), .A3(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G57gat), .B(G64gat), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n504_), .A2(KEYINPUT11), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(KEYINPUT11), .ZN(new_n506_));
  XOR2_X1   g305(.A(G71gat), .B(G78gat), .Z(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n506_), .A2(new_n507_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n503_), .A2(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(KEYINPUT69), .B1(new_n503_), .B2(new_n511_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT12), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n512_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G230gat), .A2(G233gat), .ZN(new_n517_));
  AOI211_X1 g316(.A(KEYINPUT69), .B(KEYINPUT12), .C1(new_n503_), .C2(new_n511_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n516_), .A2(new_n517_), .A3(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n503_), .A2(new_n511_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n512_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n517_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n520_), .A2(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G120gat), .B(G148gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G176gat), .B(G204gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n530_), .B(KEYINPUT71), .Z(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n525_), .A2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n520_), .A2(new_n524_), .A3(new_n530_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT13), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n533_), .B(new_n534_), .C1(KEYINPUT72), .C2(new_n538_), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT73), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G232gat), .A2(G233gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT34), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n543_), .A2(KEYINPUT35), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n544_), .B1(new_n463_), .B2(new_n503_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n545_), .B1(new_n459_), .B2(new_n503_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n543_), .A2(KEYINPUT35), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G190gat), .B(G218gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT74), .ZN(new_n550_));
  XOR2_X1   g349(.A(G134gat), .B(G162gat), .Z(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT36), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n548_), .A2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n548_), .A2(new_n553_), .A3(new_n552_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT37), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G231gat), .A2(G233gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n455_), .B(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(new_n510_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT75), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n563_), .ZN(new_n565_));
  XOR2_X1   g364(.A(G127gat), .B(G155gat), .Z(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT16), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G183gat), .B(G211gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT17), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n564_), .A2(new_n565_), .A3(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n569_), .B(new_n570_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT76), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(new_n574_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(new_n562_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n572_), .B1(new_n575_), .B2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT77), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n559_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NOR4_X1   g380(.A1(new_n448_), .A2(new_n473_), .A3(new_n541_), .A4(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n298_), .A2(new_n342_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(new_n450_), .A3(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n584_), .B(KEYINPUT100), .Z(new_n585_));
  OR2_X1    g384(.A1(new_n585_), .A2(KEYINPUT38), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(KEYINPUT38), .ZN(new_n587_));
  INV_X1    g386(.A(new_n557_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n448_), .A2(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n540_), .A2(new_n473_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n579_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT101), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n589_), .A2(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n450_), .B1(new_n594_), .B2(new_n583_), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n595_), .B(KEYINPUT102), .Z(new_n596_));
  NAND3_X1  g395(.A1(new_n586_), .A2(new_n587_), .A3(new_n596_), .ZN(G1324gat));
  INV_X1    g396(.A(new_n424_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n451_), .B1(new_n594_), .B2(new_n598_), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n599_), .A2(KEYINPUT39), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n582_), .A2(new_n451_), .A3(new_n598_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT103), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n599_), .A2(KEYINPUT39), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n600_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT40), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(G1325gat));
  INV_X1    g405(.A(G15gat), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n607_), .B1(new_n594_), .B2(new_n341_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT104), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n609_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n610_), .A2(KEYINPUT41), .A3(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n582_), .A2(new_n607_), .A3(new_n341_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(KEYINPUT41), .B1(new_n610_), .B2(new_n611_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n614_), .A2(new_n615_), .ZN(G1326gat));
  INV_X1    g415(.A(G22gat), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n617_), .B1(new_n594_), .B2(new_n445_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT42), .Z(new_n619_));
  NAND3_X1  g418(.A1(new_n582_), .A2(new_n617_), .A3(new_n445_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(G1327gat));
  INV_X1    g420(.A(KEYINPUT43), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n417_), .A2(new_n425_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n447_), .A2(new_n426_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n622_), .B1(new_n625_), .B2(new_n559_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n559_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n448_), .A2(KEYINPUT43), .A3(new_n627_), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n579_), .B(new_n590_), .C1(new_n626_), .C2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT44), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n625_), .A2(new_n622_), .A3(new_n559_), .ZN(new_n632_));
  OAI21_X1  g431(.A(KEYINPUT43), .B1(new_n448_), .B2(new_n627_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n634_), .A2(KEYINPUT44), .A3(new_n579_), .A4(new_n590_), .ZN(new_n635_));
  AND4_X1   g434(.A1(G29gat), .A2(new_n631_), .A3(new_n583_), .A4(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n579_), .A2(new_n588_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n637_), .A2(new_n540_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n625_), .A2(new_n472_), .A3(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT105), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT105), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n625_), .A2(new_n641_), .A3(new_n472_), .A4(new_n638_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(G29gat), .B1(new_n643_), .B2(new_n583_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n636_), .A2(new_n644_), .ZN(G1328gat));
  NAND3_X1  g444(.A1(new_n631_), .A2(new_n598_), .A3(new_n635_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(G36gat), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n424_), .A2(G36gat), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n640_), .A2(new_n642_), .A3(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT45), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n647_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT46), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n647_), .A2(KEYINPUT46), .A3(new_n650_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1329gat));
  INV_X1    g454(.A(G43gat), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n426_), .A2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n631_), .A2(new_n635_), .A3(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(KEYINPUT106), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT106), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n631_), .A2(new_n660_), .A3(new_n635_), .A4(new_n657_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n643_), .A2(new_n341_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(new_n656_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n659_), .A2(new_n661_), .A3(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT47), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT47), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n659_), .A2(new_n663_), .A3(new_n666_), .A4(new_n661_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(G1330gat));
  AND4_X1   g467(.A1(G50gat), .A2(new_n631_), .A3(new_n445_), .A4(new_n635_), .ZN(new_n669_));
  AOI21_X1  g468(.A(G50gat), .B1(new_n643_), .B2(new_n445_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1331gat));
  AND4_X1   g470(.A1(new_n473_), .A2(new_n589_), .A3(new_n541_), .A4(new_n591_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n672_), .A2(G57gat), .A3(new_n583_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT108), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n673_), .A2(new_n674_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n448_), .A2(new_n472_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n580_), .A2(new_n540_), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n678_), .B(KEYINPUT107), .Z(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(G57gat), .B1(new_n681_), .B2(new_n583_), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n675_), .A2(new_n676_), .A3(new_n682_), .ZN(G1332gat));
  NAND2_X1  g482(.A1(new_n672_), .A2(new_n598_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(G64gat), .ZN(new_n685_));
  XNOR2_X1  g484(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n685_), .B(new_n686_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n424_), .A2(G64gat), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT110), .Z(new_n689_));
  OAI21_X1  g488(.A(new_n687_), .B1(new_n680_), .B2(new_n689_), .ZN(G1333gat));
  AOI21_X1  g489(.A(new_n332_), .B1(new_n672_), .B2(new_n341_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT49), .Z(new_n692_));
  NAND3_X1  g491(.A1(new_n681_), .A2(new_n332_), .A3(new_n341_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1334gat));
  INV_X1    g493(.A(G78gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n681_), .A2(new_n695_), .A3(new_n445_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT50), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n672_), .A2(new_n445_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n698_), .B2(G78gat), .ZN(new_n699_));
  AOI211_X1 g498(.A(KEYINPUT50), .B(new_n695_), .C1(new_n672_), .C2(new_n445_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n696_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT111), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n701_), .B(new_n702_), .ZN(G1335gat));
  OAI21_X1  g502(.A(KEYINPUT112), .B1(new_n626_), .B2(new_n628_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT112), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n632_), .A2(new_n633_), .A3(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n540_), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n707_), .A2(new_n591_), .A3(new_n472_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n704_), .A2(new_n706_), .A3(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT113), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n710_), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n711_), .A2(new_n583_), .A3(new_n482_), .A4(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n541_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n714_), .A2(new_n637_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n677_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n583_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n485_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n713_), .A2(new_n718_), .ZN(G1336gat));
  NAND4_X1  g518(.A1(new_n711_), .A2(new_n598_), .A3(new_n483_), .A4(new_n712_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n486_), .B1(new_n716_), .B2(new_n424_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1337gat));
  INV_X1    g521(.A(new_n716_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n723_), .A2(new_n341_), .A3(new_n474_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT115), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n704_), .A2(new_n341_), .A3(new_n706_), .A4(new_n708_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT114), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n726_), .A2(new_n727_), .A3(G99gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n726_), .B2(G99gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT51), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT51), .ZN(new_n732_));
  OAI211_X1 g531(.A(new_n725_), .B(new_n732_), .C1(new_n728_), .C2(new_n729_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1338gat));
  NAND3_X1  g533(.A1(new_n723_), .A2(new_n445_), .A3(new_n475_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n707_), .A2(new_n472_), .A3(new_n266_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n634_), .A2(new_n579_), .A3(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT52), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n737_), .A2(new_n738_), .A3(G106gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n737_), .B2(G106gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n735_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g541(.A1(new_n424_), .A2(new_n341_), .A3(new_n266_), .A4(new_n583_), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n515_), .A2(new_n523_), .A3(new_n518_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n523_), .B1(new_n515_), .B2(new_n518_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(KEYINPUT55), .B2(new_n745_), .ZN(new_n746_));
  AND4_X1   g545(.A1(KEYINPUT55), .A2(new_n516_), .A3(new_n517_), .A4(new_n519_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n532_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT56), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  OAI211_X1 g549(.A(KEYINPUT56), .B(new_n532_), .C1(new_n746_), .C2(new_n747_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n464_), .A2(new_n460_), .A3(new_n466_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n465_), .A2(new_n461_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n470_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n755_), .B1(new_n470_), .B2(new_n467_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n534_), .A2(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT118), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n752_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT58), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n752_), .A2(new_n758_), .A3(KEYINPUT58), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n761_), .A2(new_n559_), .A3(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n534_), .A2(new_n472_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n745_), .A2(KEYINPUT55), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n520_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n744_), .A2(new_n745_), .A3(KEYINPUT55), .ZN(new_n767_));
  AOI211_X1 g566(.A(new_n749_), .B(new_n531_), .C1(new_n766_), .C2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT116), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n764_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n750_), .A2(KEYINPUT116), .A3(new_n751_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n535_), .A2(new_n756_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n588_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT119), .B1(new_n774_), .B2(KEYINPUT57), .ZN(new_n775_));
  AOI22_X1  g574(.A1(new_n770_), .A2(new_n771_), .B1(new_n535_), .B2(new_n756_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT119), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT57), .ZN(new_n778_));
  NOR4_X1   g577(.A1(new_n776_), .A2(new_n777_), .A3(new_n778_), .A4(new_n588_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n763_), .B1(new_n775_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT117), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n781_), .B1(new_n774_), .B2(KEYINPUT57), .ZN(new_n782_));
  OAI211_X1 g581(.A(KEYINPUT117), .B(new_n778_), .C1(new_n776_), .C2(new_n588_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n579_), .B1(new_n780_), .B2(new_n784_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n581_), .A2(new_n472_), .A3(new_n540_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n786_), .B(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n743_), .B1(new_n785_), .B2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(G113gat), .B1(new_n789_), .B2(new_n472_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT120), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT121), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT59), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n785_), .A2(new_n788_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n743_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n793_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n743_), .A2(KEYINPUT59), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n774_), .A2(KEYINPUT57), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n579_), .B1(new_n780_), .B2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n798_), .B1(new_n800_), .B2(new_n788_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n792_), .B1(new_n796_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n763_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n779_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n774_), .A2(KEYINPUT57), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n777_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n803_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n799_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n591_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n786_), .B(KEYINPUT54), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n797_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n811_), .B(KEYINPUT121), .C1(new_n793_), .C2(new_n789_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n802_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n472_), .A2(G113gat), .ZN(new_n814_));
  XOR2_X1   g613(.A(new_n814_), .B(KEYINPUT122), .Z(new_n815_));
  AOI21_X1  g614(.A(new_n791_), .B1(new_n813_), .B2(new_n815_), .ZN(G1340gat));
  INV_X1    g615(.A(G120gat), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n707_), .B2(KEYINPUT60), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n789_), .B(new_n818_), .C1(KEYINPUT60), .C2(new_n817_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n811_), .B(new_n541_), .C1(new_n793_), .C2(new_n789_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n819_), .B1(new_n821_), .B2(new_n817_), .ZN(G1341gat));
  NAND3_X1  g621(.A1(new_n802_), .A2(new_n591_), .A3(new_n812_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(G127gat), .ZN(new_n824_));
  INV_X1    g623(.A(new_n789_), .ZN(new_n825_));
  OR3_X1    g624(.A1(new_n825_), .A2(G127gat), .A3(new_n579_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(G1342gat));
  XNOR2_X1  g626(.A(KEYINPUT123), .B(G134gat), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n627_), .A2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n802_), .A2(new_n812_), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(G134gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(new_n825_), .B2(new_n557_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT124), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n830_), .A2(KEYINPUT124), .A3(new_n832_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(G1343gat));
  NOR2_X1   g636(.A1(new_n266_), .A2(new_n341_), .ZN(new_n838_));
  AND4_X1   g637(.A1(new_n583_), .A2(new_n794_), .A3(new_n424_), .A4(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n472_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g640(.A1(new_n839_), .A2(new_n541_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g642(.A1(new_n839_), .A2(new_n591_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(KEYINPUT61), .B(G155gat), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n844_), .B(new_n845_), .ZN(G1346gat));
  AOI21_X1  g645(.A(G162gat), .B1(new_n839_), .B2(new_n588_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n559_), .A2(G162gat), .ZN(new_n848_));
  XOR2_X1   g647(.A(new_n848_), .B(KEYINPUT125), .Z(new_n849_));
  AOI21_X1  g648(.A(new_n847_), .B1(new_n839_), .B2(new_n849_), .ZN(G1347gat));
  NOR2_X1   g649(.A1(new_n809_), .A2(new_n810_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n598_), .A2(new_n343_), .ZN(new_n852_));
  XOR2_X1   g651(.A(new_n852_), .B(KEYINPUT126), .Z(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n266_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n851_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n472_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n857_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n856_), .A2(new_n472_), .A3(new_n350_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(KEYINPUT62), .B1(new_n857_), .B2(G169gat), .ZN(new_n861_));
  OR2_X1    g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1348gat));
  AOI21_X1  g661(.A(G176gat), .B1(new_n856_), .B2(new_n540_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n445_), .B1(new_n785_), .B2(new_n788_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n853_), .A2(new_n303_), .A3(new_n714_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n863_), .B1(new_n864_), .B2(new_n865_), .ZN(G1349gat));
  NOR2_X1   g665(.A1(new_n579_), .A2(new_n324_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n864_), .A2(new_n591_), .A3(new_n854_), .ZN(new_n868_));
  AOI22_X1  g667(.A1(new_n856_), .A2(new_n867_), .B1(new_n868_), .B2(new_n309_), .ZN(G1350gat));
  NAND2_X1  g668(.A1(new_n588_), .A2(new_n371_), .ZN(new_n870_));
  XOR2_X1   g669(.A(new_n870_), .B(KEYINPUT127), .Z(new_n871_));
  NAND2_X1  g670(.A1(new_n856_), .A2(new_n871_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n851_), .A2(new_n855_), .A3(new_n627_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(new_n310_), .ZN(G1351gat));
  AND4_X1   g673(.A1(new_n717_), .A2(new_n794_), .A3(new_n598_), .A4(new_n838_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n472_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g676(.A1(new_n875_), .A2(new_n541_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g678(.A1(new_n875_), .A2(new_n591_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n881_));
  AND2_X1   g680(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n880_), .A2(new_n881_), .A3(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n883_), .B1(new_n880_), .B2(new_n881_), .ZN(G1354gat));
  INV_X1    g683(.A(G218gat), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n875_), .A2(new_n885_), .A3(new_n588_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n875_), .A2(new_n559_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(new_n885_), .ZN(G1355gat));
endmodule


