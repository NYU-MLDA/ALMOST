//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 1 0 0 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 0 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n787_, new_n788_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n891_, new_n892_, new_n894_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n933_, new_n934_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n941_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XOR2_X1   g002(.A(G85gat), .B(G92gat), .Z(new_n204_));
  NOR2_X1   g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT7), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT6), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n204_), .B1(new_n207_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT8), .ZN(new_n212_));
  OR3_X1    g011(.A1(new_n211_), .A2(KEYINPUT64), .A3(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(KEYINPUT8), .ZN(new_n214_));
  XOR2_X1   g013(.A(KEYINPUT10), .B(G99gat), .Z(new_n215_));
  INV_X1    g014(.A(G106gat), .ZN(new_n216_));
  AOI22_X1  g015(.A1(KEYINPUT9), .A2(new_n204_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G85gat), .ZN(new_n218_));
  INV_X1    g017(.A(G92gat), .ZN(new_n219_));
  NOR3_X1   g018(.A1(new_n218_), .A2(new_n219_), .A3(KEYINPUT9), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n210_), .A2(new_n220_), .ZN(new_n221_));
  AOI22_X1  g020(.A1(new_n211_), .A2(new_n214_), .B1(new_n217_), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n213_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G57gat), .B(G64gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT65), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT11), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n227_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G71gat), .B(G78gat), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n228_), .A2(new_n229_), .A3(new_n231_), .ZN(new_n232_));
  OR3_X1    g031(.A1(new_n226_), .A2(new_n227_), .A3(new_n231_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n224_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n223_), .A2(new_n233_), .A3(new_n232_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(KEYINPUT12), .A3(new_n236_), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n236_), .A2(KEYINPUT12), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n203_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n202_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G120gat), .B(G148gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G176gat), .B(G204gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  XOR2_X1   g044(.A(KEYINPUT67), .B(KEYINPUT5), .Z(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n241_), .B1(new_n242_), .B2(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n242_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n249_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n251_), .A2(KEYINPUT13), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n248_), .A2(KEYINPUT13), .A3(new_n250_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT37), .ZN(new_n256_));
  XOR2_X1   g055(.A(G29gat), .B(G36gat), .Z(new_n257_));
  XOR2_X1   g056(.A(G43gat), .B(G50gat), .Z(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT15), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n223_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G232gat), .A2(G233gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT35), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n259_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n261_), .B(new_n266_), .C1(new_n267_), .C2(new_n223_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n264_), .A2(new_n265_), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n269_), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT69), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(G190gat), .B(G218gat), .Z(new_n273_));
  XNOR2_X1  g072(.A(G134gat), .B(G162gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT36), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n277_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n276_), .A2(KEYINPUT36), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n272_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NOR3_X1   g080(.A1(new_n272_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n256_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n278_), .A2(new_n279_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n272_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n286_), .A2(KEYINPUT37), .A3(new_n280_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n283_), .A2(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(G127gat), .B(G155gat), .Z(new_n289_));
  XNOR2_X1  g088(.A(G183gat), .B(G211gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(KEYINPUT71), .B(KEYINPUT16), .Z(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n293_), .A2(KEYINPUT17), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G15gat), .B(G22gat), .ZN(new_n295_));
  INV_X1    g094(.A(G1gat), .ZN(new_n296_));
  INV_X1    g095(.A(G8gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT14), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n295_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G1gat), .B(G8gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G231gat), .A2(G233gat), .ZN(new_n302_));
  XOR2_X1   g101(.A(new_n301_), .B(new_n302_), .Z(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(new_n234_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT17), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n305_), .A2(KEYINPUT70), .ZN(new_n306_));
  AOI211_X1 g105(.A(new_n294_), .B(new_n304_), .C1(new_n293_), .C2(new_n306_), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n304_), .A2(new_n293_), .A3(new_n306_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n288_), .A2(new_n309_), .ZN(new_n310_));
  XOR2_X1   g109(.A(KEYINPUT98), .B(KEYINPUT27), .Z(new_n311_));
  NAND2_X1  g110(.A1(G226gat), .A2(G233gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n312_), .B(KEYINPUT90), .ZN(new_n313_));
  XOR2_X1   g112(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n314_));
  XOR2_X1   g113(.A(new_n313_), .B(new_n314_), .Z(new_n315_));
  INV_X1    g114(.A(G183gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT25), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT25), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(G183gat), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(G190gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT26), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT26), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(G190gat), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT91), .B(KEYINPUT24), .ZN(new_n326_));
  NOR2_X1   g125(.A1(G169gat), .A2(G176gat), .ZN(new_n327_));
  AOI22_X1  g126(.A1(new_n320_), .A2(new_n325_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G183gat), .A2(G190gat), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT23), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n326_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G169gat), .A2(G176gat), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n336_), .A2(new_n327_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n333_), .B1(new_n334_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(G176gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT73), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT73), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(G176gat), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT22), .B(G169gat), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n336_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n316_), .A2(new_n321_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n331_), .A2(new_n346_), .A3(new_n332_), .ZN(new_n347_));
  AOI22_X1  g146(.A1(new_n328_), .A2(new_n338_), .B1(new_n345_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT86), .ZN(new_n350_));
  INV_X1    g149(.A(G218gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(G211gat), .ZN(new_n352_));
  INV_X1    g151(.A(G211gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(G218gat), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT85), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n352_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n355_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n350_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n353_), .A2(G218gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n351_), .A2(G211gat), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT85), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n352_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n361_), .A2(KEYINPUT86), .A3(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n358_), .A2(new_n363_), .A3(KEYINPUT21), .ZN(new_n364_));
  INV_X1    g163(.A(G204gat), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n365_), .A2(G197gat), .ZN(new_n366_));
  INV_X1    g165(.A(G197gat), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT83), .B1(new_n367_), .B2(G204gat), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT83), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n369_), .A2(new_n365_), .A3(G197gat), .ZN(new_n370_));
  AOI211_X1 g169(.A(KEYINPUT87), .B(new_n366_), .C1(new_n368_), .C2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT87), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n368_), .A2(new_n370_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n366_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n372_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n371_), .A2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n364_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n361_), .A2(new_n362_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT82), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n379_), .B1(new_n365_), .B2(G197gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n365_), .A2(G197gat), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n367_), .A2(KEYINPUT82), .A3(G204gat), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n380_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT21), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n378_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT21), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n373_), .A2(new_n386_), .A3(new_n374_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT84), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n366_), .B1(new_n368_), .B2(new_n370_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT84), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n389_), .A2(new_n390_), .A3(new_n386_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n385_), .B1(new_n388_), .B2(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n349_), .B1(new_n377_), .B2(new_n392_), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n393_), .A2(KEYINPUT20), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n389_), .B(new_n372_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n386_), .B1(new_n378_), .B2(new_n350_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n395_), .A2(new_n396_), .A3(new_n363_), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n362_), .A2(new_n361_), .B1(new_n383_), .B2(KEYINPUT21), .ZN(new_n398_));
  AND4_X1   g197(.A1(new_n390_), .A2(new_n373_), .A3(new_n386_), .A4(new_n374_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n390_), .B1(new_n389_), .B2(new_n386_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n398_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n317_), .A2(new_n319_), .A3(new_n322_), .A4(new_n324_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n332_), .ZN(new_n403_));
  AOI21_X1  g202(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT24), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n327_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(G169gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n339_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n409_), .A2(KEYINPUT24), .A3(new_n335_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n402_), .A2(new_n405_), .A3(new_n407_), .A4(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n408_), .A2(KEYINPUT22), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT22), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(G169gat), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n340_), .A2(new_n342_), .A3(new_n412_), .A4(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(new_n347_), .A3(new_n335_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n411_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT74), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n411_), .A2(KEYINPUT74), .A3(new_n416_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n397_), .A2(new_n401_), .A3(new_n419_), .A4(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n315_), .B1(new_n394_), .B2(new_n421_), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n401_), .B(new_n348_), .C1(new_n376_), .C2(new_n364_), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n358_), .A2(KEYINPUT21), .A3(new_n363_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n388_), .A2(new_n391_), .ZN(new_n425_));
  AOI22_X1  g224(.A1(new_n424_), .A2(new_n395_), .B1(new_n425_), .B2(new_n398_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n420_), .ZN(new_n427_));
  AOI21_X1  g226(.A(KEYINPUT74), .B1(new_n411_), .B2(new_n416_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n423_), .B(KEYINPUT20), .C1(new_n426_), .C2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n315_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G8gat), .B(G36gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT18), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G64gat), .B(G92gat), .ZN(new_n435_));
  XOR2_X1   g234(.A(new_n434_), .B(new_n435_), .Z(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  OR3_X1    g236(.A1(new_n422_), .A2(new_n432_), .A3(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n437_), .B1(new_n422_), .B2(new_n432_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n311_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT97), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT95), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n430_), .A2(new_n442_), .A3(new_n431_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n442_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n444_));
  AND4_X1   g243(.A1(KEYINPUT20), .A2(new_n393_), .A3(new_n421_), .A4(new_n315_), .ZN(new_n445_));
  NOR3_X1   g244(.A1(new_n443_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n441_), .B1(new_n446_), .B2(new_n436_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n444_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n430_), .A2(new_n442_), .A3(new_n431_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n445_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n451_), .A2(KEYINPUT97), .A3(new_n437_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n447_), .A2(new_n452_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n438_), .A2(KEYINPUT27), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n440_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  XOR2_X1   g254(.A(G1gat), .B(G29gat), .Z(new_n456_));
  XNOR2_X1  g255(.A(G57gat), .B(G85gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(G155gat), .A2(G162gat), .ZN(new_n461_));
  AND2_X1   g260(.A1(G155gat), .A2(G162gat), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT1), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n461_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G155gat), .A2(G162gat), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n465_), .A2(KEYINPUT78), .A3(KEYINPUT1), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(KEYINPUT78), .B1(new_n465_), .B2(KEYINPUT1), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n464_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G141gat), .A2(G148gat), .ZN(new_n470_));
  INV_X1    g269(.A(G141gat), .ZN(new_n471_));
  INV_X1    g270(.A(G148gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n469_), .A2(new_n470_), .A3(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT79), .B1(new_n462_), .B2(new_n461_), .ZN(new_n475_));
  INV_X1    g274(.A(G155gat), .ZN(new_n476_));
  INV_X1    g275(.A(G162gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT79), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n478_), .A2(new_n479_), .A3(new_n465_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n475_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT3), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n482_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT2), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n470_), .A2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n483_), .A2(new_n485_), .A3(new_n486_), .A4(new_n487_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n481_), .A2(KEYINPUT80), .A3(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(KEYINPUT80), .B1(new_n481_), .B2(new_n488_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n474_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT76), .ZN(new_n492_));
  INV_X1    g291(.A(G127gat), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n493_), .A2(G134gat), .ZN(new_n494_));
  INV_X1    g293(.A(G134gat), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n495_), .A2(G127gat), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n492_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(G127gat), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n493_), .A2(G134gat), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n498_), .A2(new_n499_), .A3(KEYINPUT76), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G113gat), .B(G120gat), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n497_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n501_), .B1(new_n497_), .B2(new_n500_), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n491_), .A2(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n502_), .A2(new_n503_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n506_), .B(new_n474_), .C1(new_n490_), .C2(new_n489_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n507_), .A3(KEYINPUT4), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT92), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n505_), .A2(new_n507_), .A3(KEYINPUT92), .A4(KEYINPUT4), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G225gat), .A2(G233gat), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n514_), .B1(new_n505_), .B2(KEYINPUT4), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n512_), .A2(KEYINPUT93), .A3(new_n516_), .ZN(new_n517_));
  AND2_X1   g316(.A1(new_n505_), .A2(new_n507_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(new_n513_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n515_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n521_), .A2(KEYINPUT93), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n460_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT96), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n521_), .A2(KEYINPUT93), .B1(new_n518_), .B2(new_n513_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n512_), .A2(new_n516_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT93), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n460_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n525_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n523_), .A2(new_n524_), .A3(new_n530_), .ZN(new_n531_));
  OAI211_X1 g330(.A(KEYINPUT96), .B(new_n460_), .C1(new_n520_), .C2(new_n522_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n455_), .A2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n506_), .B(KEYINPUT31), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G71gat), .B(G99gat), .ZN(new_n537_));
  INV_X1    g336(.A(G43gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G227gat), .A2(G233gat), .ZN(new_n540_));
  INV_X1    g339(.A(G15gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n539_), .B(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT30), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n427_), .A2(new_n428_), .A3(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(KEYINPUT30), .B1(new_n419_), .B2(new_n420_), .ZN(new_n546_));
  OAI21_X1  g345(.A(KEYINPUT75), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n544_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n419_), .A2(KEYINPUT30), .A3(new_n420_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT75), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n548_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n543_), .B1(new_n547_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n543_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n536_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n543_), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n548_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n550_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n556_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n559_), .A2(new_n553_), .A3(new_n535_), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n555_), .A2(KEYINPUT77), .A3(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(KEYINPUT77), .B1(new_n555_), .B2(new_n560_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n473_), .A2(new_n470_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n468_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(new_n466_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n564_), .B1(new_n566_), .B2(new_n464_), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n462_), .A2(new_n461_), .A3(KEYINPUT79), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n479_), .B1(new_n478_), .B2(new_n465_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n488_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT80), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n481_), .A2(KEYINPUT80), .A3(new_n488_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n567_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT29), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n576_), .B(KEYINPUT28), .Z(new_n577_));
  OAI22_X1  g376(.A1(new_n392_), .A2(new_n377_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT88), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n579_), .B1(new_n377_), .B2(new_n392_), .ZN(new_n580_));
  INV_X1    g379(.A(G228gat), .ZN(new_n581_));
  INV_X1    g380(.A(G233gat), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n578_), .A2(new_n580_), .A3(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G78gat), .B(G106gat), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n397_), .A2(new_n401_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n491_), .A2(KEYINPUT29), .ZN(new_n587_));
  INV_X1    g386(.A(new_n583_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n586_), .B(new_n587_), .C1(new_n579_), .C2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n584_), .A2(new_n585_), .A3(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(KEYINPUT81), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n585_), .B1(new_n584_), .B2(new_n589_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n577_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G22gat), .B(G50gat), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n584_), .A2(new_n589_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n585_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n577_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n597_), .A2(new_n598_), .A3(KEYINPUT81), .A4(new_n590_), .ZN(new_n599_));
  AND3_X1   g398(.A1(new_n593_), .A2(new_n594_), .A3(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n594_), .B1(new_n593_), .B2(new_n599_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n563_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n593_), .A2(new_n599_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n594_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n555_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n560_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n593_), .A2(new_n594_), .A3(new_n599_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n605_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n602_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n436_), .A2(KEYINPUT32), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n612_), .B1(new_n422_), .B2(new_n432_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n613_), .B1(new_n451_), .B2(new_n612_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n531_), .A2(new_n532_), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT33), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n530_), .A2(new_n616_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n438_), .A2(new_n439_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n525_), .A2(new_n528_), .A3(KEYINPUT33), .A4(new_n529_), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n512_), .B(new_n513_), .C1(KEYINPUT4), .C2(new_n505_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n518_), .A2(new_n514_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n620_), .A2(new_n460_), .A3(new_n621_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n617_), .A2(new_n618_), .A3(new_n619_), .A4(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n615_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n562_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n555_), .A2(new_n560_), .A3(KEYINPUT77), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NOR3_X1   g426(.A1(new_n627_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n628_));
  AOI22_X1  g427(.A1(new_n534_), .A2(new_n611_), .B1(new_n624_), .B2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n260_), .A2(new_n301_), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n267_), .A2(new_n301_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(G229gat), .A2(G233gat), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n630_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n267_), .B(new_n301_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n632_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n633_), .A2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(G113gat), .B(G141gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G169gat), .B(G197gat), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n638_), .B(new_n639_), .Z(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n637_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n633_), .A2(new_n636_), .A3(new_n640_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT72), .Z(new_n645_));
  OAI21_X1  g444(.A(KEYINPUT99), .B1(new_n629_), .B2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n611_), .A2(new_n533_), .A3(new_n455_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n624_), .A2(new_n628_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT99), .ZN(new_n650_));
  INV_X1    g449(.A(new_n645_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n649_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n652_));
  AOI211_X1 g451(.A(new_n255_), .B(new_n310_), .C1(new_n646_), .C2(new_n652_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n653_), .A2(new_n296_), .A3(new_n532_), .A4(new_n531_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n655_));
  OR3_X1    g454(.A1(new_n654_), .A2(KEYINPUT101), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n286_), .A2(new_n280_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n629_), .A2(new_n657_), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n658_), .A2(new_n644_), .A3(new_n254_), .A4(new_n309_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n659_), .A2(new_n533_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n660_), .A2(new_n296_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n654_), .B1(new_n661_), .B2(new_n655_), .ZN(new_n662_));
  OAI21_X1  g461(.A(KEYINPUT101), .B1(new_n654_), .B2(new_n655_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n656_), .A2(new_n662_), .A3(new_n663_), .ZN(G1324gat));
  OAI21_X1  g463(.A(G8gat), .B1(new_n659_), .B2(new_n455_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT39), .ZN(new_n666_));
  INV_X1    g465(.A(new_n455_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n653_), .A2(new_n297_), .A3(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT40), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(G1325gat));
  OAI21_X1  g470(.A(G15gat), .B1(new_n659_), .B2(new_n563_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n672_), .B(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n653_), .A2(new_n541_), .A3(new_n627_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n676_), .B(new_n677_), .ZN(G1326gat));
  NOR2_X1   g477(.A1(new_n600_), .A2(new_n601_), .ZN(new_n679_));
  OAI21_X1  g478(.A(G22gat), .B1(new_n659_), .B2(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT42), .ZN(new_n681_));
  INV_X1    g480(.A(G22gat), .ZN(new_n682_));
  INV_X1    g481(.A(new_n679_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n653_), .A2(new_n682_), .A3(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n681_), .A2(new_n684_), .ZN(G1327gat));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n686_));
  INV_X1    g485(.A(new_n657_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n686_), .B1(new_n687_), .B2(new_n309_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n309_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n657_), .A2(KEYINPUT104), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(new_n254_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n646_), .B2(new_n652_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n694_), .A2(new_n533_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n695_), .A2(G29gat), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n254_), .A2(new_n644_), .A3(new_n689_), .ZN(new_n698_));
  OAI21_X1  g497(.A(KEYINPUT43), .B1(new_n629_), .B2(new_n288_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n700_));
  INV_X1    g499(.A(new_n288_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n602_), .A2(new_n610_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n455_), .A2(new_n533_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n679_), .A2(new_n563_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(new_n615_), .B2(new_n623_), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n700_), .B(new_n701_), .C1(new_n704_), .C2(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n698_), .B1(new_n699_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT103), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n697_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  AOI211_X1 g509(.A(KEYINPUT103), .B(new_n698_), .C1(new_n699_), .C2(new_n707_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n712_), .B1(KEYINPUT44), .B2(new_n708_), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n531_), .A2(G29gat), .A3(new_n532_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n696_), .B1(new_n713_), .B2(new_n714_), .ZN(G1328gat));
  INV_X1    g514(.A(KEYINPUT106), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n716_), .A2(KEYINPUT46), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n455_), .B1(new_n708_), .B2(KEYINPUT44), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n718_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n717_), .B1(new_n719_), .B2(G36gat), .ZN(new_n720_));
  INV_X1    g519(.A(new_n692_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n455_), .A2(G36gat), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n629_), .A2(KEYINPUT99), .A3(new_n645_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n650_), .B1(new_n649_), .B2(new_n651_), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n721_), .B(new_n722_), .C1(new_n723_), .C2(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n725_), .A2(KEYINPUT105), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n727_), .B1(new_n693_), .B2(new_n722_), .ZN(new_n728_));
  OAI21_X1  g527(.A(KEYINPUT45), .B1(new_n726_), .B2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n725_), .A2(KEYINPUT105), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT45), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n693_), .A2(new_n727_), .A3(new_n722_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n730_), .A2(new_n731_), .A3(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n729_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n716_), .A2(KEYINPUT46), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n720_), .A2(new_n734_), .A3(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n720_), .B2(new_n734_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n736_), .A2(new_n737_), .ZN(G1329gat));
  XOR2_X1   g537(.A(KEYINPUT107), .B(G43gat), .Z(new_n739_));
  OAI21_X1  g538(.A(new_n739_), .B1(new_n694_), .B2(new_n563_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n708_), .A2(KEYINPUT44), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n741_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n608_), .A2(G43gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n740_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g544(.A(G50gat), .B1(new_n693_), .B2(new_n683_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n683_), .A2(G50gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n713_), .B2(new_n747_), .ZN(G1331gat));
  NAND4_X1  g547(.A1(new_n658_), .A2(new_n645_), .A3(new_n255_), .A4(new_n309_), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT108), .Z(new_n750_));
  NAND3_X1  g549(.A1(new_n750_), .A2(new_n532_), .A3(new_n531_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(G57gat), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n629_), .A2(new_n644_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n310_), .A2(new_n254_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n533_), .A2(G57gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n752_), .B1(new_n755_), .B2(new_n756_), .ZN(G1332gat));
  INV_X1    g556(.A(KEYINPUT48), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n750_), .A2(new_n667_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n759_), .B2(G64gat), .ZN(new_n760_));
  INV_X1    g559(.A(G64gat), .ZN(new_n761_));
  AOI211_X1 g560(.A(KEYINPUT48), .B(new_n761_), .C1(new_n750_), .C2(new_n667_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n667_), .A2(new_n761_), .ZN(new_n763_));
  OAI22_X1  g562(.A1(new_n760_), .A2(new_n762_), .B1(new_n755_), .B2(new_n763_), .ZN(G1333gat));
  INV_X1    g563(.A(KEYINPUT49), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n750_), .A2(new_n627_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(G71gat), .ZN(new_n767_));
  INV_X1    g566(.A(G71gat), .ZN(new_n768_));
  AOI211_X1 g567(.A(KEYINPUT49), .B(new_n768_), .C1(new_n750_), .C2(new_n627_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n627_), .A2(new_n768_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT109), .ZN(new_n771_));
  OAI22_X1  g570(.A1(new_n767_), .A2(new_n769_), .B1(new_n755_), .B2(new_n771_), .ZN(G1334gat));
  OR3_X1    g571(.A1(new_n755_), .A2(G78gat), .A3(new_n679_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n750_), .A2(new_n683_), .ZN(new_n774_));
  XOR2_X1   g573(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n775_));
  AND3_X1   g574(.A1(new_n774_), .A2(G78gat), .A3(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n774_), .B2(G78gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n776_), .B2(new_n777_), .ZN(G1335gat));
  AND3_X1   g577(.A1(new_n753_), .A2(new_n255_), .A3(new_n691_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n779_), .A2(new_n218_), .A3(new_n532_), .A4(new_n531_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n644_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n255_), .A2(new_n781_), .A3(new_n689_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n782_), .B1(new_n699_), .B2(new_n707_), .ZN(new_n783_));
  XOR2_X1   g582(.A(new_n783_), .B(KEYINPUT111), .Z(new_n784_));
  AND3_X1   g583(.A1(new_n784_), .A2(new_n532_), .A3(new_n531_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n780_), .B1(new_n785_), .B2(new_n218_), .ZN(G1336gat));
  NAND3_X1  g585(.A1(new_n779_), .A2(new_n219_), .A3(new_n667_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n784_), .A2(new_n667_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n787_), .B1(new_n788_), .B2(new_n219_), .ZN(G1337gat));
  NAND2_X1  g588(.A1(new_n783_), .A2(new_n627_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(G99gat), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n779_), .A2(new_n608_), .A3(new_n215_), .ZN(new_n792_));
  XOR2_X1   g591(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n793_));
  NAND3_X1  g592(.A1(new_n791_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT114), .ZN(new_n795_));
  INV_X1    g594(.A(new_n791_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n792_), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT51), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT112), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n798_), .A2(new_n799_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n795_), .B1(new_n800_), .B2(new_n801_), .ZN(G1338gat));
  NAND3_X1  g601(.A1(new_n779_), .A2(new_n216_), .A3(new_n683_), .ZN(new_n803_));
  AOI211_X1 g602(.A(KEYINPUT115), .B(new_n216_), .C1(new_n783_), .C2(new_n683_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT115), .ZN(new_n805_));
  INV_X1    g604(.A(new_n782_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n700_), .B1(new_n649_), .B2(new_n701_), .ZN(new_n807_));
  AOI211_X1 g606(.A(KEYINPUT43), .B(new_n288_), .C1(new_n647_), .C2(new_n648_), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n683_), .B(new_n806_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n805_), .B1(new_n809_), .B2(G106gat), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n804_), .A2(new_n810_), .A3(KEYINPUT52), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n812_));
  AOI211_X1 g611(.A(new_n679_), .B(new_n782_), .C1(new_n699_), .C2(new_n707_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT115), .B1(new_n813_), .B2(new_n216_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n809_), .A2(new_n805_), .A3(G106gat), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n812_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n803_), .B1(new_n811_), .B2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT53), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n819_), .B(new_n803_), .C1(new_n811_), .C2(new_n816_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(G1339gat));
  NAND4_X1  g620(.A1(new_n254_), .A2(new_n288_), .A3(new_n645_), .A4(new_n309_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n822_), .B(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n239_), .A2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n237_), .A2(new_n238_), .A3(new_n203_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n247_), .B1(new_n239_), .B2(new_n825_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n828_), .A2(new_n829_), .A3(KEYINPUT116), .A4(KEYINPUT56), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n781_), .B1(new_n241_), .B2(new_n247_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT56), .B1(new_n828_), .B2(new_n829_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n833_), .A2(KEYINPUT116), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n828_), .A2(KEYINPUT56), .A3(new_n829_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n832_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n640_), .B1(new_n634_), .B2(new_n632_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT117), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n630_), .A2(new_n631_), .A3(new_n635_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n643_), .B1(new_n839_), .B2(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n251_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n687_), .B1(new_n836_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845_));
  OAI21_X1  g644(.A(KEYINPUT118), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT58), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n842_), .B1(new_n241_), .B2(new_n247_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n835_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(new_n833_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n288_), .B1(new_n847_), .B2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n847_), .B2(new_n850_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n849_), .A2(KEYINPUT116), .A3(new_n833_), .ZN(new_n853_));
  OAI22_X1  g652(.A1(new_n853_), .A2(new_n832_), .B1(new_n251_), .B2(new_n842_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT118), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n854_), .A2(new_n855_), .A3(KEYINPUT57), .A4(new_n687_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n844_), .A2(new_n845_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n846_), .A2(new_n852_), .A3(new_n856_), .A4(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n824_), .B1(new_n858_), .B2(new_n689_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n667_), .A2(new_n533_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n860_), .A2(new_n608_), .A3(new_n679_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(KEYINPUT119), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  OAI22_X1  g662(.A1(new_n859_), .A2(new_n863_), .B1(KEYINPUT120), .B2(KEYINPUT59), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n858_), .A2(new_n689_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n824_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n862_), .ZN(new_n868_));
  XOR2_X1   g667(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n869_));
  OAI21_X1  g668(.A(new_n864_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  XOR2_X1   g669(.A(KEYINPUT121), .B(G113gat), .Z(new_n871_));
  NOR3_X1   g670(.A1(new_n870_), .A2(new_n645_), .A3(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n868_), .A2(new_n781_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(G113gat), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n872_), .A2(new_n874_), .ZN(G1340gat));
  OAI21_X1  g674(.A(G120gat), .B1(new_n870_), .B2(new_n254_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT60), .ZN(new_n877_));
  AOI21_X1  g676(.A(G120gat), .B1(new_n255_), .B2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n878_), .B1(new_n877_), .B2(G120gat), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n867_), .A2(new_n862_), .A3(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n876_), .A2(new_n880_), .ZN(G1341gat));
  NOR3_X1   g680(.A1(new_n859_), .A2(new_n689_), .A3(new_n863_), .ZN(new_n882_));
  OR3_X1    g681(.A1(new_n882_), .A2(KEYINPUT122), .A3(G127gat), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n689_), .A2(new_n493_), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n864_), .B(new_n884_), .C1(new_n868_), .C2(new_n869_), .ZN(new_n885_));
  OAI21_X1  g684(.A(KEYINPUT122), .B1(new_n882_), .B2(G127gat), .ZN(new_n886_));
  AND3_X1   g685(.A1(new_n883_), .A2(new_n885_), .A3(new_n886_), .ZN(G1342gat));
  OAI21_X1  g686(.A(G134gat), .B1(new_n870_), .B2(new_n288_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n657_), .A2(new_n495_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n868_), .B2(new_n889_), .ZN(G1343gat));
  NOR2_X1   g689(.A1(new_n859_), .A2(new_n602_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n891_), .A2(new_n644_), .A3(new_n860_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g692(.A1(new_n891_), .A2(new_n255_), .A3(new_n860_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g694(.A1(new_n891_), .A2(new_n309_), .A3(new_n860_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(KEYINPUT61), .B(G155gat), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n896_), .B(new_n897_), .ZN(G1346gat));
  NAND4_X1  g697(.A1(new_n891_), .A2(new_n477_), .A3(new_n657_), .A4(new_n860_), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n891_), .A2(new_n701_), .A3(new_n860_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(new_n477_), .ZN(G1347gat));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT62), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n455_), .B1(new_n532_), .B2(new_n531_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n627_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n644_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT123), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n907_), .B(new_n908_), .ZN(new_n909_));
  NOR3_X1   g708(.A1(new_n859_), .A2(new_n683_), .A3(new_n909_), .ZN(new_n910_));
  OAI211_X1 g709(.A(new_n902_), .B(new_n903_), .C1(new_n910_), .C2(new_n408_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n859_), .A2(new_n683_), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n912_), .A2(new_n344_), .A3(new_n644_), .A4(new_n906_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n902_), .B1(new_n910_), .B2(new_n408_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(KEYINPUT62), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n910_), .A2(new_n902_), .A3(new_n408_), .ZN(new_n916_));
  OAI211_X1 g715(.A(new_n911_), .B(new_n913_), .C1(new_n915_), .C2(new_n916_), .ZN(G1348gat));
  NAND2_X1  g716(.A1(new_n912_), .A2(KEYINPUT125), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT125), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n919_), .B1(new_n859_), .B2(new_n683_), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n918_), .A2(new_n920_), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n905_), .A2(new_n339_), .A3(new_n254_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n912_), .A2(new_n255_), .A3(new_n906_), .ZN(new_n923_));
  AOI22_X1  g722(.A1(new_n921_), .A2(new_n922_), .B1(new_n343_), .B2(new_n923_), .ZN(G1349gat));
  NOR2_X1   g723(.A1(new_n689_), .A2(new_n320_), .ZN(new_n925_));
  NAND4_X1  g724(.A1(new_n867_), .A2(new_n679_), .A3(new_n906_), .A4(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(KEYINPUT126), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT126), .ZN(new_n928_));
  NAND4_X1  g727(.A1(new_n912_), .A2(new_n928_), .A3(new_n906_), .A4(new_n925_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n929_), .ZN(new_n930_));
  NAND4_X1  g729(.A1(new_n918_), .A2(new_n309_), .A3(new_n906_), .A4(new_n920_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n316_), .B2(new_n931_), .ZN(G1350gat));
  AND2_X1   g731(.A1(new_n657_), .A2(new_n325_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n912_), .A2(new_n906_), .A3(new_n933_), .ZN(new_n934_));
  NOR4_X1   g733(.A1(new_n859_), .A2(new_n683_), .A3(new_n288_), .A4(new_n905_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n935_), .B2(new_n321_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(KEYINPUT127), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT127), .ZN(new_n938_));
  OAI211_X1 g737(.A(new_n934_), .B(new_n938_), .C1(new_n321_), .C2(new_n935_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n937_), .A2(new_n939_), .ZN(G1351gat));
  NAND3_X1  g739(.A1(new_n891_), .A2(new_n644_), .A3(new_n904_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g741(.A1(new_n891_), .A2(new_n255_), .A3(new_n904_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(G204gat), .ZN(G1353gat));
  AND3_X1   g743(.A1(new_n891_), .A2(new_n309_), .A3(new_n904_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n946_));
  AND2_X1   g745(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n945_), .B1(new_n946_), .B2(new_n947_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n948_), .B1(new_n945_), .B2(new_n946_), .ZN(G1354gat));
  NAND4_X1  g748(.A1(new_n891_), .A2(new_n351_), .A3(new_n657_), .A4(new_n904_), .ZN(new_n950_));
  AND3_X1   g749(.A1(new_n891_), .A2(new_n701_), .A3(new_n904_), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n950_), .B1(new_n951_), .B2(new_n351_), .ZN(G1355gat));
endmodule


