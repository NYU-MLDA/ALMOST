//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 0 0 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n860_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT20), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(G197gat), .B(G204gat), .Z(new_n206_));
  XNOR2_X1  g005(.A(G211gat), .B(G218gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n206_), .B1(KEYINPUT21), .B2(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT21), .B1(new_n207_), .B2(KEYINPUT86), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  AND3_X1   g009(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n211_));
  AOI21_X1  g010(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT24), .ZN(new_n214_));
  INV_X1    g013(.A(G169gat), .ZN(new_n215_));
  INV_X1    g014(.A(G176gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n213_), .A2(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n215_), .A2(new_n216_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220_));
  NOR3_X1   g019(.A1(new_n219_), .A2(new_n214_), .A3(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n218_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT25), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(G183gat), .ZN(new_n224_));
  INV_X1    g023(.A(G183gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT25), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT88), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(KEYINPUT25), .B(G183gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT88), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT26), .B(G190gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n229_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  OR2_X1    g032(.A1(G183gat), .A2(G190gat), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n219_), .B1(new_n213_), .B2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT22), .B(G169gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(new_n216_), .ZN(new_n237_));
  AOI22_X1  g036(.A1(new_n222_), .A2(new_n233_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT90), .ZN(new_n239_));
  AND3_X1   g038(.A1(new_n210_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n239_), .B1(new_n210_), .B2(new_n238_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n205_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n210_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT77), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n224_), .A2(new_n244_), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n232_), .B(new_n245_), .C1(new_n230_), .C2(new_n244_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n221_), .ZN(new_n247_));
  AOI21_X1  g046(.A(KEYINPUT78), .B1(new_n213_), .B2(new_n217_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G183gat), .A2(G190gat), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT23), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n252_));
  AND4_X1   g051(.A1(KEYINPUT78), .A2(new_n217_), .A3(new_n251_), .A4(new_n252_), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n246_), .B(new_n247_), .C1(new_n248_), .C2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT80), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n237_), .A2(KEYINPUT79), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT79), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n236_), .A2(new_n257_), .A3(new_n216_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(new_n235_), .A3(new_n258_), .ZN(new_n259_));
  AND3_X1   g058(.A1(new_n254_), .A2(new_n255_), .A3(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n255_), .B1(new_n254_), .B2(new_n259_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n243_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(KEYINPUT89), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n254_), .A2(new_n259_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT80), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n254_), .A2(new_n255_), .A3(new_n259_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT89), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(new_n268_), .A3(new_n243_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n242_), .B1(new_n263_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n203_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n210_), .A2(new_n238_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n272_), .A2(new_n204_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n265_), .A2(new_n266_), .A3(new_n210_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n271_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G8gat), .B(G36gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT18), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(G64gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(G92gat), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT32), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NOR3_X1   g080(.A1(new_n270_), .A2(new_n275_), .A3(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n273_), .A2(new_n274_), .A3(new_n271_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n210_), .A2(new_n238_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(KEYINPUT20), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n285_), .B1(new_n263_), .B2(new_n269_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n283_), .B1(new_n286_), .B2(new_n271_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n282_), .B1(new_n287_), .B2(new_n281_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G155gat), .B(G162gat), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n289_), .A2(KEYINPUT1), .ZN(new_n290_));
  INV_X1    g089(.A(G141gat), .ZN(new_n291_));
  INV_X1    g090(.A(G148gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G141gat), .A2(G148gat), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n290_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT3), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n298_), .A2(new_n291_), .A3(new_n292_), .A4(KEYINPUT83), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT83), .ZN(new_n300_));
  OAI22_X1  g099(.A1(new_n300_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT2), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n295_), .A2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n299_), .A2(new_n301_), .A3(new_n303_), .A4(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT84), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n289_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n303_), .A2(new_n304_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n308_), .A2(KEYINPUT84), .A3(new_n301_), .A4(new_n299_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n297_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G127gat), .B(G134gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G113gat), .B(G120gat), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n312_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT91), .B1(new_n310_), .B2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n307_), .A2(new_n309_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n297_), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n317_), .A2(new_n315_), .A3(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n316_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n310_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n315_), .ZN(new_n322_));
  NOR3_X1   g121(.A1(new_n321_), .A2(KEYINPUT91), .A3(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT4), .B1(new_n320_), .B2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G225gat), .A2(G233gat), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  OR3_X1    g125(.A1(new_n310_), .A2(KEYINPUT4), .A3(new_n315_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n324_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n325_), .B1(new_n320_), .B2(new_n323_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G1gat), .B(G29gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(KEYINPUT0), .ZN(new_n331_));
  INV_X1    g130(.A(G57gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(G85gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n333_), .B(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n328_), .A2(new_n329_), .A3(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n336_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT95), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n337_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  AOI211_X1 g139(.A(KEYINPUT95), .B(new_n336_), .C1(new_n328_), .C2(new_n329_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n288_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT96), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT96), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n288_), .B(new_n344_), .C1(new_n340_), .C2(new_n341_), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n316_), .A2(new_n319_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n323_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT93), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT93), .B1(new_n320_), .B2(new_n323_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(new_n350_), .A3(new_n326_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(new_n335_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT94), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n351_), .A2(KEYINPUT94), .A3(new_n335_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n324_), .A2(new_n325_), .A3(new_n327_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n270_), .A2(new_n275_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(new_n279_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT33), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n337_), .B1(KEYINPUT92), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(KEYINPUT92), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n337_), .A2(KEYINPUT92), .A3(new_n360_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n357_), .A2(new_n359_), .A3(new_n363_), .A4(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n343_), .A2(new_n345_), .A3(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n210_), .B1(new_n321_), .B2(KEYINPUT29), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G228gat), .A2(G233gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G78gat), .B(G106gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n369_), .A2(new_n370_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n321_), .A2(KEYINPUT29), .ZN(new_n375_));
  XOR2_X1   g174(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n376_));
  XNOR2_X1  g175(.A(G22gat), .B(G50gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n375_), .B(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n379_), .B1(new_n371_), .B2(KEYINPUT87), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n374_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n374_), .A2(new_n380_), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n366_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT97), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT97), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n366_), .A2(new_n387_), .A3(new_n384_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n340_), .A2(new_n341_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n383_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  OR2_X1    g190(.A1(new_n359_), .A2(KEYINPUT27), .ZN(new_n392_));
  INV_X1    g191(.A(new_n279_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n358_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n287_), .ZN(new_n395_));
  XOR2_X1   g194(.A(new_n279_), .B(KEYINPUT98), .Z(new_n396_));
  OAI211_X1 g195(.A(new_n394_), .B(KEYINPUT27), .C1(new_n395_), .C2(new_n396_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n392_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n391_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n386_), .A2(new_n388_), .A3(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G15gat), .B(G43gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G71gat), .B(G99gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G227gat), .A2(G233gat), .ZN(new_n404_));
  XOR2_X1   g203(.A(new_n403_), .B(new_n404_), .Z(new_n405_));
  XOR2_X1   g204(.A(new_n267_), .B(KEYINPUT30), .Z(new_n406_));
  OR2_X1    g205(.A1(new_n406_), .A2(KEYINPUT81), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(KEYINPUT81), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n405_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n408_), .A2(new_n405_), .ZN(new_n410_));
  OR2_X1    g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(KEYINPUT82), .B(KEYINPUT31), .Z(new_n412_));
  XNOR2_X1  g211(.A(new_n315_), .B(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n411_), .B(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n400_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n398_), .A2(new_n384_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n389_), .ZN(new_n418_));
  NOR3_X1   g217(.A1(new_n417_), .A2(new_n415_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n416_), .A2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G15gat), .B(G22gat), .ZN(new_n422_));
  INV_X1    g221(.A(G1gat), .ZN(new_n423_));
  INV_X1    g222(.A(G8gat), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT14), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n422_), .A2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G1gat), .B(G8gat), .ZN(new_n427_));
  XOR2_X1   g226(.A(new_n426_), .B(new_n427_), .Z(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(G50gat), .ZN(new_n430_));
  INV_X1    g229(.A(G36gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(G29gat), .ZN(new_n432_));
  INV_X1    g231(.A(G29gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(G36gat), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT68), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n432_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n435_), .B1(new_n432_), .B2(new_n434_), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n437_), .A2(new_n438_), .A3(G43gat), .ZN(new_n439_));
  INV_X1    g238(.A(G43gat), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n433_), .A2(G36gat), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n431_), .A2(G29gat), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT68), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n440_), .B1(new_n443_), .B2(new_n436_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n430_), .B1(new_n439_), .B2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(G43gat), .B1(new_n437_), .B2(new_n438_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n443_), .A2(new_n440_), .A3(new_n436_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n446_), .A2(new_n447_), .A3(G50gat), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n445_), .A2(KEYINPUT15), .A3(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(KEYINPUT15), .B1(new_n445_), .B2(new_n448_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n429_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G229gat), .A2(G233gat), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n445_), .A2(new_n428_), .A3(new_n448_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n451_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n428_), .B1(new_n445_), .B2(new_n448_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n453_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n452_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G113gat), .B(G141gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(new_n215_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(G197gat), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n454_), .A2(new_n459_), .A3(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT75), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT76), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT76), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n463_), .A2(new_n464_), .A3(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n466_), .A2(new_n468_), .ZN(new_n469_));
  AND2_X1   g268(.A1(new_n454_), .A2(new_n459_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n470_), .A2(new_n462_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n469_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n466_), .A2(new_n471_), .A3(new_n468_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n421_), .A2(KEYINPUT99), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT99), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n419_), .B1(new_n400_), .B2(new_n415_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n478_), .B1(new_n479_), .B2(new_n475_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT7), .ZN(new_n482_));
  INV_X1    g281(.A(G99gat), .ZN(new_n483_));
  INV_X1    g282(.A(G106gat), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G99gat), .A2(G106gat), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT6), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n490_));
  NAND4_X1  g289(.A1(new_n485_), .A2(new_n488_), .A3(new_n489_), .A4(new_n490_), .ZN(new_n491_));
  OR2_X1    g290(.A1(G85gat), .A2(G92gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G85gat), .A2(G92gat), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n491_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(KEYINPUT64), .A2(KEYINPUT8), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n491_), .A2(new_n496_), .A3(new_n494_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(KEYINPUT10), .B(G99gat), .Z(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n484_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n488_), .A2(new_n489_), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n493_), .A2(KEYINPUT9), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n492_), .A2(KEYINPUT9), .A3(new_n493_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .A4(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n500_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G71gat), .B(G78gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G57gat), .B(G64gat), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT11), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n508_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n509_), .A2(KEYINPUT11), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n509_), .A2(new_n508_), .A3(KEYINPUT11), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT12), .B1(new_n507_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n507_), .A2(new_n516_), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n516_), .A2(KEYINPUT12), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT66), .ZN(new_n522_));
  INV_X1    g321(.A(new_n506_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n523_), .B1(new_n500_), .B2(KEYINPUT65), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT65), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n498_), .A2(new_n525_), .A3(new_n499_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n522_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n491_), .A2(new_n496_), .A3(new_n494_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n496_), .B1(new_n491_), .B2(new_n494_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT65), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n530_), .A2(new_n526_), .A3(new_n522_), .A4(new_n506_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n521_), .B1(new_n527_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT67), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n519_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n530_), .A2(new_n526_), .A3(new_n506_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT66), .ZN(new_n537_));
  AOI211_X1 g336(.A(new_n534_), .B(new_n520_), .C1(new_n537_), .C2(new_n531_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G230gat), .A2(G233gat), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n535_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n540_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n518_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n507_), .A2(new_n516_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n542_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n541_), .A2(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(G120gat), .B(G148gat), .Z(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(G204gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT5), .B(G176gat), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n548_), .B(new_n549_), .Z(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n546_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n546_), .A2(new_n551_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT13), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n553_), .A2(KEYINPUT13), .A3(new_n554_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G127gat), .B(G155gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT16), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(new_n225_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(G211gat), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT17), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  AND2_X1   g364(.A1(new_n563_), .A2(new_n564_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n429_), .B(new_n516_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G231gat), .A2(G233gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT74), .ZN(new_n570_));
  AOI211_X1 g369(.A(new_n565_), .B(new_n566_), .C1(new_n569_), .C2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n571_), .B1(new_n570_), .B2(new_n569_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n565_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT73), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n572_), .A2(new_n575_), .ZN(new_n576_));
  OAI22_X1  g375(.A1(new_n527_), .A2(new_n532_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n577_));
  AND4_X1   g376(.A1(new_n448_), .A2(new_n445_), .A3(new_n500_), .A4(new_n506_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G232gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT34), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT35), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT70), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n580_), .A2(KEYINPUT35), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n578_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n577_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n586_), .A2(new_n582_), .A3(new_n581_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n581_), .A2(new_n582_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n577_), .A2(new_n588_), .A3(new_n585_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G134gat), .B(G162gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT69), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(G190gat), .ZN(new_n593_));
  INV_X1    g392(.A(G218gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n595_), .A2(KEYINPUT36), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(KEYINPUT36), .ZN(new_n597_));
  OAI21_X1  g396(.A(KEYINPUT72), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n597_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n595_), .A2(KEYINPUT36), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT72), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n599_), .A2(new_n600_), .A3(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n590_), .B1(new_n598_), .B2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(KEYINPUT37), .B1(new_n603_), .B2(KEYINPUT71), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n599_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n604_), .B(new_n606_), .ZN(new_n607_));
  AND4_X1   g406(.A1(new_n481_), .A2(new_n559_), .A3(new_n576_), .A4(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n608_), .A2(new_n423_), .A3(new_n418_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT38), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n479_), .A2(new_n606_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n559_), .A2(new_n476_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n576_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(G1gat), .B1(new_n616_), .B2(new_n389_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n609_), .A2(new_n610_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n618_), .A2(KEYINPUT100), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(KEYINPUT100), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n611_), .B(new_n617_), .C1(new_n619_), .C2(new_n620_), .ZN(G1324gat));
  OAI21_X1  g420(.A(G8gat), .B1(new_n616_), .B2(new_n398_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n623_), .A2(KEYINPUT101), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(KEYINPUT101), .ZN(new_n625_));
  OR3_X1    g424(.A1(new_n622_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n398_), .A2(G8gat), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n608_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n622_), .A2(new_n624_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n626_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n630_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g430(.A(G15gat), .B1(new_n616_), .B2(new_n415_), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n632_), .B(KEYINPUT41), .Z(new_n633_));
  INV_X1    g432(.A(G15gat), .ZN(new_n634_));
  INV_X1    g433(.A(new_n415_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n608_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n633_), .A2(new_n636_), .ZN(G1326gat));
  OAI21_X1  g436(.A(G22gat), .B1(new_n616_), .B2(new_n384_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT42), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n384_), .A2(G22gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT102), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n608_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n639_), .A2(new_n642_), .ZN(G1327gat));
  INV_X1    g442(.A(new_n606_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n644_), .A2(new_n576_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n559_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n481_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(G29gat), .B1(new_n649_), .B2(new_n418_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n613_), .A2(new_n576_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(KEYINPUT43), .B1(new_n479_), .B2(new_n607_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT43), .ZN(new_n654_));
  INV_X1    g453(.A(new_n607_), .ZN(new_n655_));
  AOI22_X1  g454(.A1(new_n385_), .A2(KEYINPUT97), .B1(new_n391_), .B2(new_n398_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n635_), .B1(new_n656_), .B2(new_n388_), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n654_), .B(new_n655_), .C1(new_n657_), .C2(new_n419_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n652_), .B1(new_n653_), .B2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(KEYINPUT44), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n661_), .A2(new_n433_), .A3(new_n389_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n653_), .A2(new_n658_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(new_n651_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT103), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n659_), .A2(KEYINPUT103), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n666_), .A2(new_n667_), .A3(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n650_), .B1(new_n662_), .B2(new_n669_), .ZN(G1328gat));
  XNOR2_X1  g469(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n398_), .A2(KEYINPUT104), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n398_), .A2(KEYINPUT104), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n675_), .A2(G36gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(KEYINPUT99), .B1(new_n421_), .B2(new_n476_), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n479_), .A2(new_n478_), .A3(new_n475_), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n647_), .B(new_n676_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n680_), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n481_), .A2(new_n647_), .A3(new_n682_), .A4(new_n676_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n398_), .B1(new_n659_), .B2(KEYINPUT44), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n667_), .B1(new_n659_), .B2(KEYINPUT103), .ZN(new_n686_));
  AOI211_X1 g485(.A(new_n665_), .B(new_n652_), .C1(new_n653_), .C2(new_n658_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n685_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n684_), .B1(new_n688_), .B2(G36gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n672_), .B1(new_n689_), .B2(KEYINPUT106), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT106), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n431_), .B1(new_n669_), .B2(new_n685_), .ZN(new_n692_));
  OAI211_X1 g491(.A(new_n691_), .B(new_n671_), .C1(new_n692_), .C2(new_n684_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n690_), .A2(new_n693_), .ZN(G1329gat));
  XNOR2_X1  g493(.A(KEYINPUT109), .B(G43gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n695_), .B1(new_n648_), .B2(new_n415_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT108), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n635_), .A2(G43gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(new_n659_), .B2(KEYINPUT44), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n697_), .B1(new_n669_), .B2(new_n699_), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n697_), .B(new_n699_), .C1(new_n686_), .C2(new_n687_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n696_), .B1(new_n700_), .B2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT47), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT47), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n705_), .B(new_n696_), .C1(new_n700_), .C2(new_n702_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1330gat));
  AOI21_X1  g506(.A(G50gat), .B1(new_n649_), .B2(new_n383_), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n661_), .A2(new_n430_), .A3(new_n384_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n709_), .B2(new_n669_), .ZN(G1331gat));
  NOR3_X1   g509(.A1(new_n559_), .A2(new_n476_), .A3(new_n614_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n612_), .A2(new_n711_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n712_), .A2(new_n332_), .A3(new_n389_), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n421_), .A2(new_n607_), .A3(new_n711_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n715_), .A2(KEYINPUT110), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n389_), .B1(new_n715_), .B2(KEYINPUT110), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n713_), .B1(new_n718_), .B2(new_n332_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT111), .Z(G1332gat));
  OAI21_X1  g519(.A(G64gat), .B1(new_n712_), .B2(new_n675_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT48), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n675_), .A2(G64gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(new_n715_), .B2(new_n723_), .ZN(G1333gat));
  OAI21_X1  g523(.A(G71gat), .B1(new_n712_), .B2(new_n415_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT49), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n415_), .A2(G71gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n715_), .B2(new_n727_), .ZN(G1334gat));
  OAI21_X1  g527(.A(G78gat), .B1(new_n712_), .B2(new_n384_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT50), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n384_), .A2(G78gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n715_), .B2(new_n731_), .ZN(G1335gat));
  NOR2_X1   g531(.A1(new_n559_), .A2(new_n476_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(new_n614_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n734_), .B1(new_n653_), .B2(new_n658_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(G85gat), .B1(new_n736_), .B2(new_n389_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n733_), .A2(new_n645_), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n479_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n740_), .A2(new_n334_), .A3(new_n418_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n737_), .A2(new_n741_), .ZN(G1336gat));
  OAI21_X1  g541(.A(G92gat), .B1(new_n736_), .B2(new_n675_), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n398_), .A2(G92gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(new_n739_), .B2(new_n744_), .ZN(G1337gat));
  NAND2_X1  g544(.A1(new_n735_), .A2(new_n635_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n635_), .A2(new_n501_), .ZN(new_n747_));
  AOI22_X1  g546(.A1(new_n746_), .A2(G99gat), .B1(new_n740_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT51), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT112), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n748_), .A2(new_n749_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT113), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(G1338gat));
  NAND3_X1  g553(.A1(new_n740_), .A2(new_n484_), .A3(new_n383_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT52), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n735_), .A2(new_n383_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n757_), .B2(G106gat), .ZN(new_n758_));
  AOI211_X1 g557(.A(KEYINPUT52), .B(new_n484_), .C1(new_n735_), .C2(new_n383_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n755_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  XOR2_X1   g559(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n761_));
  XNOR2_X1  g560(.A(new_n760_), .B(new_n761_), .ZN(G1339gat));
  NAND2_X1  g561(.A1(new_n517_), .A2(new_n518_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n520_), .B1(new_n537_), .B2(new_n531_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n764_), .B2(KEYINPUT67), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n765_), .A2(new_n542_), .A3(new_n538_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n542_), .B1(new_n765_), .B2(new_n538_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(KEYINPUT55), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769_));
  NOR4_X1   g568(.A1(new_n765_), .A2(new_n538_), .A3(new_n769_), .A4(new_n542_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n551_), .B1(new_n768_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT56), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n540_), .B1(new_n535_), .B2(new_n539_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n541_), .B1(new_n774_), .B2(new_n769_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n770_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n550_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT56), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n773_), .A2(new_n778_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n451_), .A2(new_n453_), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n780_), .A2(KEYINPUT116), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(KEYINPUT116), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(new_n458_), .A3(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n462_), .B1(new_n457_), .B2(new_n452_), .ZN(new_n784_));
  AOI22_X1  g583(.A1(new_n783_), .A2(new_n784_), .B1(new_n470_), .B2(new_n462_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n553_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n779_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT58), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n779_), .A2(KEYINPUT58), .A3(new_n786_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n655_), .A3(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n772_), .B1(new_n777_), .B2(KEYINPUT115), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n771_), .A2(new_n794_), .A3(KEYINPUT56), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n552_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n793_), .A2(new_n795_), .A3(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n555_), .A2(new_n785_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n792_), .B1(new_n799_), .B2(new_n644_), .ZN(new_n800_));
  AOI211_X1 g599(.A(KEYINPUT57), .B(new_n606_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n791_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT117), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  OAI211_X1 g603(.A(KEYINPUT117), .B(new_n791_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(new_n614_), .A3(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT118), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n559_), .A2(new_n607_), .A3(new_n475_), .A4(new_n576_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n808_), .B(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n806_), .A2(new_n807_), .A3(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n807_), .B1(new_n806_), .B2(new_n811_), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n417_), .A2(new_n415_), .A3(new_n389_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n812_), .A2(new_n813_), .A3(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(G113gat), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(new_n817_), .A3(new_n476_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT119), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n810_), .B1(new_n614_), .B2(new_n802_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT59), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n814_), .A2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n819_), .B1(new_n820_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n822_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n802_), .A2(new_n614_), .ZN(new_n825_));
  OAI211_X1 g624(.A(KEYINPUT119), .B(new_n824_), .C1(new_n825_), .C2(new_n810_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n823_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n806_), .A2(new_n811_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT118), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n806_), .A2(new_n807_), .A3(new_n811_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n830_), .A3(new_n814_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n827_), .B1(new_n831_), .B2(KEYINPUT59), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n832_), .A2(new_n476_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n818_), .B1(new_n833_), .B2(new_n817_), .ZN(G1340gat));
  INV_X1    g633(.A(new_n559_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n827_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n835_), .B(new_n836_), .C1(new_n816_), .C2(new_n821_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT121), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(KEYINPUT120), .B(G120gat), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n832_), .A2(KEYINPUT121), .A3(new_n835_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n839_), .A2(new_n841_), .A3(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n840_), .B1(new_n559_), .B2(KEYINPUT60), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n816_), .B(new_n844_), .C1(KEYINPUT60), .C2(new_n840_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(G1341gat));
  INV_X1    g645(.A(G127gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n816_), .A2(new_n847_), .A3(new_n576_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n832_), .A2(new_n576_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(new_n847_), .ZN(G1342gat));
  INV_X1    g649(.A(G134gat), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n816_), .A2(new_n851_), .A3(new_n606_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n832_), .A2(new_n655_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n851_), .ZN(G1343gat));
  NOR2_X1   g653(.A1(new_n812_), .A2(new_n813_), .ZN(new_n855_));
  AND4_X1   g654(.A1(new_n415_), .A2(new_n675_), .A3(new_n383_), .A4(new_n418_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n475_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(new_n291_), .ZN(G1344gat));
  NOR2_X1   g658(.A1(new_n857_), .A2(new_n559_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(new_n292_), .ZN(G1345gat));
  INV_X1    g660(.A(new_n857_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n576_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(KEYINPUT61), .B(G155gat), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n863_), .B(new_n864_), .ZN(G1346gat));
  AOI21_X1  g664(.A(G162gat), .B1(new_n862_), .B2(new_n606_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n655_), .A2(G162gat), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(KEYINPUT122), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n866_), .B1(new_n862_), .B2(new_n868_), .ZN(G1347gat));
  NOR3_X1   g668(.A1(new_n675_), .A2(new_n415_), .A3(new_n418_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n384_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n820_), .A2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(G169gat), .B1(new_n873_), .B2(new_n475_), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n874_), .A2(KEYINPUT123), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(KEYINPUT123), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n875_), .A2(KEYINPUT62), .A3(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n872_), .A2(new_n236_), .A3(new_n476_), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n877_), .B(new_n878_), .C1(KEYINPUT62), .C2(new_n876_), .ZN(G1348gat));
  AOI21_X1  g678(.A(G176gat), .B1(new_n872_), .B2(new_n835_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n812_), .A2(new_n813_), .A3(new_n383_), .ZN(new_n881_));
  AND3_X1   g680(.A1(new_n870_), .A2(G176gat), .A3(new_n835_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n880_), .B1(new_n881_), .B2(new_n882_), .ZN(G1349gat));
  AOI211_X1 g682(.A(new_n614_), .B(new_n873_), .C1(new_n229_), .C2(new_n231_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n881_), .A2(new_n576_), .A3(new_n870_), .ZN(new_n885_));
  OR2_X1    g684(.A1(new_n885_), .A2(KEYINPUT124), .ZN(new_n886_));
  AOI21_X1  g685(.A(G183gat), .B1(new_n885_), .B2(KEYINPUT124), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n884_), .B1(new_n886_), .B2(new_n887_), .ZN(G1350gat));
  OAI21_X1  g687(.A(G190gat), .B1(new_n873_), .B2(new_n607_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n872_), .A2(new_n232_), .A3(new_n606_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1351gat));
  NOR3_X1   g690(.A1(new_n675_), .A2(new_n635_), .A3(new_n390_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n855_), .A2(new_n892_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n476_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g695(.A1(new_n893_), .A2(new_n559_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT125), .ZN(new_n898_));
  AND2_X1   g697(.A1(new_n898_), .A2(G204gat), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n898_), .A2(G204gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n897_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n901_), .B1(new_n897_), .B2(new_n900_), .ZN(G1353gat));
  INV_X1    g701(.A(KEYINPUT126), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n855_), .A2(new_n576_), .A3(new_n892_), .ZN(new_n904_));
  XOR2_X1   g703(.A(KEYINPUT63), .B(G211gat), .Z(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n903_), .B1(new_n904_), .B2(new_n906_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n904_), .A2(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n907_), .A2(new_n909_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n904_), .A2(new_n903_), .A3(new_n906_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1354gat));
  NAND4_X1  g711(.A1(new_n829_), .A2(new_n655_), .A3(new_n830_), .A4(new_n892_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(G218gat), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n606_), .A2(new_n594_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n914_), .B1(new_n893_), .B2(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT127), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n916_), .B(new_n917_), .ZN(G1355gat));
endmodule


