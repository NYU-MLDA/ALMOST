//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 0 0 1 0 0 0 1 1 1 0 0 0 0 1 1 0 0 1 1 0 0 0 0 0 1 0 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n878_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n916_, new_n917_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_;
  NAND2_X1  g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT87), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT90), .B(KEYINPUT2), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT91), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT91), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n203_), .A2(new_n207_), .A3(new_n204_), .ZN(new_n208_));
  INV_X1    g007(.A(G141gat), .ZN(new_n209_));
  INV_X1    g008(.A(G148gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(new_n210_), .A3(KEYINPUT3), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT3), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n212_), .B1(G141gat), .B2(G148gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n202_), .ZN(new_n214_));
  AOI22_X1  g013(.A1(new_n211_), .A2(new_n213_), .B1(new_n214_), .B2(KEYINPUT2), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n206_), .A2(new_n208_), .A3(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n217_), .B1(new_n219_), .B2(KEYINPUT1), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT88), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n222_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT89), .ZN(new_n225_));
  OR3_X1    g024(.A1(new_n217_), .A2(new_n225_), .A3(KEYINPUT1), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n225_), .B1(new_n217_), .B2(KEYINPUT1), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n223_), .A2(new_n224_), .A3(new_n226_), .A4(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n203_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n229_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n230_));
  AOI22_X1  g029(.A1(new_n216_), .A2(new_n220_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G113gat), .B(G120gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT84), .ZN(new_n233_));
  XOR2_X1   g032(.A(G127gat), .B(G134gat), .Z(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n231_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT85), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n233_), .A2(new_n234_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n233_), .A2(new_n234_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n237_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n237_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n236_), .B1(new_n243_), .B2(new_n231_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT4), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G225gat), .A2(G233gat), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n241_), .B1(new_n235_), .B2(new_n237_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n216_), .A2(new_n220_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n230_), .A2(new_n228_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(KEYINPUT4), .B1(new_n248_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n245_), .A2(new_n247_), .A3(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n248_), .A2(new_n251_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n247_), .B1(new_n255_), .B2(new_n236_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n254_), .A2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G1gat), .B(G29gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(G85gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT0), .B(G57gat), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n260_), .B(new_n261_), .Z(new_n262_));
  NAND2_X1  g061(.A1(new_n258_), .A2(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n252_), .B1(KEYINPUT4), .B2(new_n244_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n256_), .B1(new_n264_), .B2(new_n247_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n262_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n263_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n248_), .B(KEYINPUT86), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT31), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n243_), .B(KEYINPUT86), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT31), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n272_), .A2(new_n274_), .A3(KEYINPUT83), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G15gat), .B(G43gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT82), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT30), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n275_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n278_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n272_), .A2(new_n274_), .A3(KEYINPUT83), .A4(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G183gat), .A2(G190gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT23), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT80), .B(G183gat), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n284_), .B1(G190gat), .B2(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(G169gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT81), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT24), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n292_), .B1(G169gat), .B2(G176gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT81), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n290_), .B(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(new_n292_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n294_), .A2(new_n297_), .A3(new_n284_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT26), .B(G190gat), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n285_), .A2(KEYINPUT25), .ZN(new_n301_));
  OR2_X1    g100(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n300_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n289_), .B1(new_n298_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G227gat), .A2(G233gat), .ZN(new_n305_));
  INV_X1    g104(.A(G71gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(G99gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n304_), .B(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n282_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n279_), .A2(new_n309_), .A3(new_n281_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT20), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n294_), .A2(new_n297_), .A3(new_n284_), .ZN(new_n315_));
  XOR2_X1   g114(.A(KEYINPUT25), .B(G183gat), .Z(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT96), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n299_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n315_), .A2(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n284_), .B1(G183gat), .B2(G190gat), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(new_n288_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G197gat), .B(G204gat), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT21), .ZN(new_n324_));
  OR2_X1    g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n324_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G211gat), .B(G218gat), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n325_), .A2(new_n326_), .A3(new_n327_), .ZN(new_n328_));
  OR3_X1    g127(.A1(new_n323_), .A2(new_n327_), .A3(new_n324_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n314_), .B1(new_n322_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G226gat), .A2(G233gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT19), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n304_), .A2(new_n330_), .ZN(new_n335_));
  AND3_X1   g134(.A1(new_n331_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  AOI22_X1  g135(.A1(new_n315_), .A2(new_n318_), .B1(new_n288_), .B2(new_n320_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n330_), .B1(new_n337_), .B2(KEYINPUT101), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT101), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n322_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n304_), .A2(new_n330_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT97), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT97), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n304_), .A2(new_n344_), .A3(new_n330_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n341_), .A2(KEYINPUT20), .A3(new_n343_), .A4(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n336_), .B1(new_n346_), .B2(new_n333_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT102), .ZN(new_n348_));
  XOR2_X1   g147(.A(G8gat), .B(G36gat), .Z(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G64gat), .B(G92gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  OR3_X1    g152(.A1(new_n347_), .A2(new_n348_), .A3(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n348_), .B1(new_n347_), .B2(new_n353_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n331_), .A2(new_n335_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(new_n333_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n330_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n333_), .B1(new_n337_), .B2(new_n359_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n360_), .A2(new_n343_), .A3(KEYINPUT20), .A4(new_n345_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n358_), .A2(new_n353_), .A3(new_n361_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n362_), .A2(KEYINPUT27), .ZN(new_n363_));
  INV_X1    g162(.A(new_n353_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n361_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n334_), .B1(new_n331_), .B2(new_n335_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n364_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(new_n362_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT103), .B(KEYINPUT27), .ZN(new_n369_));
  AOI22_X1  g168(.A1(new_n356_), .A2(new_n363_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT29), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n231_), .A2(new_n371_), .ZN(new_n372_));
  XOR2_X1   g171(.A(G22gat), .B(G50gat), .Z(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT28), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n372_), .B(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(G78gat), .B(G106gat), .Z(new_n376_));
  OAI21_X1  g175(.A(new_n330_), .B1(new_n231_), .B2(new_n371_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n330_), .A2(KEYINPUT93), .ZN(new_n378_));
  OAI21_X1  g177(.A(G233gat), .B1(KEYINPUT92), .B2(G228gat), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n379_), .B1(KEYINPUT92), .B2(G228gat), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n377_), .A2(new_n378_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n378_), .A2(new_n380_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n382_), .B(new_n330_), .C1(new_n231_), .C2(new_n371_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n376_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n375_), .B1(new_n384_), .B2(KEYINPUT94), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT95), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT95), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n387_), .B(new_n375_), .C1(new_n384_), .C2(KEYINPUT94), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n381_), .A2(new_n383_), .A3(new_n376_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n390_), .A2(new_n384_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n389_), .B(new_n392_), .ZN(new_n393_));
  AND4_X1   g192(.A1(new_n269_), .A2(new_n313_), .A3(new_n370_), .A4(new_n393_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n353_), .A2(KEYINPUT32), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n358_), .A2(KEYINPUT100), .A3(new_n361_), .ZN(new_n396_));
  AND3_X1   g195(.A1(new_n347_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  NOR3_X1   g196(.A1(new_n365_), .A2(new_n366_), .A3(KEYINPUT100), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n398_), .A2(new_n395_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n268_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n264_), .A2(new_n247_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n266_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n367_), .B(new_n362_), .C1(new_n401_), .C2(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT33), .B1(new_n265_), .B2(new_n266_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n266_), .B1(new_n254_), .B2(new_n257_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT33), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n403_), .B1(new_n404_), .B2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n400_), .B1(new_n408_), .B2(KEYINPUT99), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n245_), .A2(new_n253_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n402_), .B1(new_n410_), .B2(new_n246_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n368_), .A2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n405_), .A2(new_n406_), .ZN(new_n413_));
  NOR3_X1   g212(.A1(new_n265_), .A2(KEYINPUT33), .A3(new_n266_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n412_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT99), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n393_), .B1(new_n409_), .B2(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n389_), .A2(new_n392_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n391_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n420_));
  NOR3_X1   g219(.A1(new_n419_), .A2(new_n268_), .A3(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n370_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n418_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n313_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n394_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(G29gat), .B(G36gat), .Z(new_n426_));
  INV_X1    g225(.A(KEYINPUT70), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G29gat), .B(G36gat), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT70), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G43gat), .B(G50gat), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n428_), .A2(new_n430_), .A3(new_n432_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(G1gat), .ZN(new_n438_));
  INV_X1    g237(.A(G8gat), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT14), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n440_), .A2(KEYINPUT74), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(KEYINPUT74), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G15gat), .B(G22gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n441_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  XOR2_X1   g243(.A(G1gat), .B(G8gat), .Z(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n437_), .B(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n447_), .A2(G229gat), .A3(G233gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n437_), .A2(KEYINPUT15), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT15), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n436_), .A2(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n446_), .B1(new_n449_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n446_), .A2(new_n437_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G229gat), .A2(G233gat), .ZN(new_n454_));
  XOR2_X1   g253(.A(new_n454_), .B(KEYINPUT78), .Z(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n448_), .B1(new_n452_), .B2(new_n456_), .ZN(new_n457_));
  XOR2_X1   g256(.A(G113gat), .B(G141gat), .Z(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT79), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G169gat), .B(G197gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n457_), .B(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G57gat), .B(G64gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(KEYINPUT11), .ZN(new_n466_));
  XOR2_X1   g265(.A(G71gat), .B(G78gat), .Z(new_n467_));
  OR2_X1    g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n465_), .A2(KEYINPUT11), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n466_), .A2(new_n467_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n468_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT12), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G99gat), .A2(G106gat), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT65), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n476_), .A2(KEYINPUT6), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT6), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n478_), .A2(KEYINPUT65), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n475_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(KEYINPUT65), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n476_), .A2(KEYINPUT6), .ZN(new_n482_));
  AND2_X1   g281(.A1(G99gat), .A2(G106gat), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT7), .ZN(new_n486_));
  INV_X1    g285(.A(G99gat), .ZN(new_n487_));
  INV_X1    g286(.A(G106gat), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n480_), .A2(new_n484_), .A3(new_n485_), .A4(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT8), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G85gat), .A2(G92gat), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(G85gat), .A2(G92gat), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  AND3_X1   g294(.A1(new_n490_), .A2(new_n491_), .A3(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n491_), .B1(new_n490_), .B2(new_n495_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT66), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT9), .ZN(new_n500_));
  OR2_X1    g299(.A1(G85gat), .A2(G92gat), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n500_), .B1(new_n501_), .B2(new_n492_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n505_));
  OAI21_X1  g304(.A(G92gat), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n502_), .B1(new_n500_), .B2(new_n506_), .ZN(new_n507_));
  OR2_X1    g306(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(new_n488_), .A3(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n480_), .A2(new_n484_), .A3(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n499_), .B1(new_n507_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n484_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n483_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT9), .B1(new_n493_), .B2(new_n494_), .ZN(new_n516_));
  INV_X1    g315(.A(G92gat), .ZN(new_n517_));
  OR2_X1    g316(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n517_), .B1(new_n518_), .B2(new_n503_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n516_), .B1(new_n519_), .B2(KEYINPUT9), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n515_), .A2(new_n520_), .A3(KEYINPUT66), .A4(new_n510_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n512_), .A2(new_n521_), .ZN(new_n522_));
  NOR3_X1   g321(.A1(new_n498_), .A2(new_n522_), .A3(KEYINPUT67), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT67), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n512_), .A2(new_n521_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n489_), .A2(new_n485_), .ZN(new_n526_));
  NOR3_X1   g325(.A1(new_n513_), .A2(new_n514_), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n495_), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT8), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n490_), .A2(new_n491_), .A3(new_n495_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n524_), .B1(new_n525_), .B2(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n474_), .B1(new_n523_), .B2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n515_), .A2(new_n520_), .A3(new_n510_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n534_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n535_));
  AOI21_X1  g334(.A(KEYINPUT12), .B1(new_n535_), .B2(new_n472_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n471_), .B(new_n534_), .C1(new_n496_), .C2(new_n497_), .ZN(new_n538_));
  INV_X1    g337(.A(G230gat), .ZN(new_n539_));
  INV_X1    g338(.A(G233gat), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n538_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n533_), .A2(new_n537_), .A3(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT68), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n539_), .A2(new_n540_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n535_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n546_), .A2(new_n471_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n538_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n545_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(KEYINPUT67), .B1(new_n498_), .B2(new_n522_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n525_), .A2(new_n531_), .A3(new_n524_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n536_), .B1(new_n552_), .B2(new_n474_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT68), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n553_), .A2(new_n554_), .A3(new_n542_), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n544_), .A2(new_n549_), .A3(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(G120gat), .B(G148gat), .Z(new_n557_));
  XNOR2_X1  g356(.A(G176gat), .B(G204gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n556_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n556_), .A2(new_n562_), .ZN(new_n564_));
  AND3_X1   g363(.A1(new_n563_), .A2(KEYINPUT13), .A3(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(KEYINPUT13), .B1(new_n563_), .B2(new_n564_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G232gat), .A2(G233gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT34), .ZN(new_n569_));
  OAI22_X1  g368(.A1(new_n535_), .A2(new_n436_), .B1(KEYINPUT35), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT71), .ZN(new_n571_));
  OAI211_X1 g370(.A(KEYINPUT35), .B(new_n569_), .C1(new_n570_), .C2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n449_), .A2(new_n451_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n552_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n570_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n572_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT35), .ZN(new_n577_));
  INV_X1    g376(.A(new_n569_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n531_), .A2(new_n437_), .A3(new_n534_), .ZN(new_n579_));
  AOI211_X1 g378(.A(new_n577_), .B(new_n578_), .C1(new_n579_), .C2(KEYINPUT71), .ZN(new_n580_));
  AOI22_X1  g379(.A1(new_n550_), .A2(new_n551_), .B1(new_n449_), .B2(new_n451_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n580_), .B1(new_n581_), .B2(new_n570_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n576_), .A2(new_n582_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n583_), .A2(KEYINPUT73), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G190gat), .B(G218gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT72), .ZN(new_n586_));
  XOR2_X1   g385(.A(G134gat), .B(G162gat), .Z(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n588_), .B1(new_n583_), .B2(KEYINPUT36), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(KEYINPUT36), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n584_), .B1(new_n589_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n583_), .A2(KEYINPUT73), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT36), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n594_), .B1(new_n576_), .B2(new_n582_), .ZN(new_n595_));
  OAI211_X1 g394(.A(new_n593_), .B(new_n590_), .C1(new_n595_), .C2(new_n588_), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n592_), .A2(KEYINPUT37), .A3(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(KEYINPUT37), .B1(new_n592_), .B2(new_n596_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n471_), .B(new_n600_), .Z(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT75), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(new_n446_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT77), .ZN(new_n604_));
  XOR2_X1   g403(.A(G127gat), .B(G155gat), .Z(new_n605_));
  XNOR2_X1  g404(.A(G183gat), .B(G211gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(KEYINPUT17), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n604_), .B(new_n610_), .ZN(new_n611_));
  OR3_X1    g410(.A1(new_n603_), .A2(KEYINPUT17), .A3(new_n609_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n567_), .A2(new_n599_), .A3(new_n613_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n425_), .A2(new_n464_), .A3(new_n614_), .ZN(new_n615_));
  XOR2_X1   g414(.A(new_n615_), .B(KEYINPUT104), .Z(new_n616_));
  NAND3_X1  g415(.A1(new_n616_), .A2(new_n438_), .A3(new_n268_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT38), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n592_), .A2(new_n596_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n425_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n567_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n613_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n623_), .A2(new_n464_), .A3(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n622_), .A2(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G1gat), .B1(new_n626_), .B2(new_n269_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n617_), .A2(new_n618_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n619_), .A2(new_n627_), .A3(new_n628_), .ZN(G1324gat));
  NOR2_X1   g428(.A1(new_n370_), .A2(G8gat), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n616_), .A2(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G8gat), .B1(new_n626_), .B2(new_n370_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n632_), .A2(KEYINPUT39), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(KEYINPUT39), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n631_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT40), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n631_), .B(KEYINPUT40), .C1(new_n633_), .C2(new_n634_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(G1325gat));
  OAI21_X1  g438(.A(G15gat), .B1(new_n626_), .B2(new_n424_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT41), .Z(new_n641_));
  INV_X1    g440(.A(G15gat), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n616_), .A2(new_n642_), .A3(new_n313_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(G1326gat));
  OAI21_X1  g443(.A(G22gat), .B1(new_n626_), .B2(new_n393_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT42), .ZN(new_n646_));
  INV_X1    g445(.A(G22gat), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n419_), .A2(new_n420_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n616_), .A2(new_n647_), .A3(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n649_), .ZN(G1327gat));
  INV_X1    g449(.A(KEYINPUT106), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n624_), .A2(new_n567_), .A3(new_n463_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT43), .ZN(new_n654_));
  INV_X1    g453(.A(new_n599_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n313_), .B1(new_n418_), .B2(new_n422_), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n654_), .B(new_n655_), .C1(new_n656_), .C2(new_n394_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n355_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n347_), .A2(new_n348_), .A3(new_n353_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n363_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n368_), .A2(new_n369_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n663_), .A2(new_n648_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n664_), .A2(new_n313_), .A3(new_n269_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n415_), .A2(new_n416_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n408_), .A2(KEYINPUT99), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n666_), .A2(new_n667_), .A3(new_n400_), .ZN(new_n668_));
  AOI22_X1  g467(.A1(new_n668_), .A2(new_n393_), .B1(new_n421_), .B2(new_n370_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n665_), .B1(new_n669_), .B2(new_n313_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n654_), .B1(new_n670_), .B2(new_n655_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n653_), .B1(new_n658_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT44), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(KEYINPUT43), .B1(new_n425_), .B2(new_n599_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(new_n657_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n676_), .A2(KEYINPUT44), .A3(new_n653_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n674_), .A2(new_n268_), .A3(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(G29gat), .ZN(new_n679_));
  INV_X1    g478(.A(G29gat), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n623_), .A2(new_n613_), .A3(new_n620_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n670_), .A2(new_n681_), .A3(new_n463_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT105), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT105), .ZN(new_n684_));
  NAND4_X1  g483(.A1(new_n670_), .A2(new_n681_), .A3(new_n684_), .A4(new_n463_), .ZN(new_n685_));
  AND4_X1   g484(.A1(new_n680_), .A2(new_n683_), .A3(new_n268_), .A4(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n651_), .B1(new_n679_), .B2(new_n687_), .ZN(new_n688_));
  AOI211_X1 g487(.A(KEYINPUT106), .B(new_n686_), .C1(new_n678_), .C2(G29gat), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1328gat));
  INV_X1    g489(.A(KEYINPUT46), .ZN(new_n691_));
  INV_X1    g490(.A(G36gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(KEYINPUT44), .B1(new_n676_), .B2(new_n653_), .ZN(new_n693_));
  AOI211_X1 g492(.A(new_n673_), .B(new_n652_), .C1(new_n675_), .C2(new_n657_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n692_), .B1(new_n695_), .B2(new_n663_), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n683_), .A2(new_n692_), .A3(new_n663_), .A4(new_n685_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT45), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n691_), .B1(new_n696_), .B2(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n697_), .B(KEYINPUT45), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n693_), .A2(new_n694_), .A3(new_n370_), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n701_), .B(KEYINPUT46), .C1(new_n702_), .C2(new_n692_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n700_), .A2(new_n703_), .ZN(G1329gat));
  AND2_X1   g503(.A1(new_n313_), .A2(G43gat), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n674_), .A2(new_n677_), .A3(new_n705_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n683_), .A2(new_n685_), .ZN(new_n707_));
  AOI21_X1  g506(.A(G43gat), .B1(new_n707_), .B2(new_n313_), .ZN(new_n708_));
  OR3_X1    g507(.A1(new_n706_), .A2(KEYINPUT47), .A3(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(KEYINPUT47), .B1(new_n706_), .B2(new_n708_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1330gat));
  INV_X1    g510(.A(G50gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n707_), .A2(new_n712_), .A3(new_n648_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n695_), .A2(new_n714_), .A3(new_n648_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(G50gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n714_), .B1(new_n695_), .B2(new_n648_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n713_), .B1(new_n716_), .B2(new_n717_), .ZN(G1331gat));
  NOR2_X1   g517(.A1(new_n425_), .A2(new_n463_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n655_), .A2(new_n624_), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n719_), .A2(new_n623_), .A3(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(G57gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(new_n722_), .A3(new_n268_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n624_), .A2(new_n567_), .A3(new_n463_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n622_), .A2(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(G57gat), .B1(new_n725_), .B2(new_n269_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n723_), .A2(new_n726_), .ZN(G1332gat));
  OAI21_X1  g526(.A(G64gat), .B1(new_n725_), .B2(new_n370_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT48), .ZN(new_n729_));
  INV_X1    g528(.A(G64gat), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n721_), .A2(new_n730_), .A3(new_n663_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(G1333gat));
  NAND3_X1  g531(.A1(new_n721_), .A2(new_n306_), .A3(new_n313_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n622_), .A2(new_n313_), .A3(new_n724_), .ZN(new_n734_));
  XOR2_X1   g533(.A(KEYINPUT108), .B(KEYINPUT49), .Z(new_n735_));
  AND3_X1   g534(.A1(new_n734_), .A2(G71gat), .A3(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n734_), .B2(G71gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n733_), .B1(new_n736_), .B2(new_n737_), .ZN(G1334gat));
  OAI21_X1  g537(.A(G78gat), .B1(new_n725_), .B2(new_n393_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT50), .ZN(new_n740_));
  INV_X1    g539(.A(G78gat), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n721_), .A2(new_n741_), .A3(new_n648_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(G1335gat));
  NOR3_X1   g542(.A1(new_n567_), .A2(new_n613_), .A3(new_n620_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n719_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(G85gat), .B1(new_n746_), .B2(new_n268_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n567_), .A2(new_n463_), .A3(new_n613_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n676_), .A2(new_n748_), .ZN(new_n749_));
  XOR2_X1   g548(.A(new_n749_), .B(KEYINPUT109), .Z(new_n750_));
  AOI21_X1  g549(.A(new_n269_), .B1(new_n518_), .B2(new_n503_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n747_), .B1(new_n750_), .B2(new_n751_), .ZN(G1336gat));
  OAI21_X1  g551(.A(new_n517_), .B1(new_n745_), .B2(new_n370_), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT110), .Z(new_n754_));
  NOR2_X1   g553(.A1(new_n370_), .A2(new_n517_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n750_), .B2(new_n755_), .ZN(G1337gat));
  NAND4_X1  g555(.A1(new_n746_), .A2(new_n313_), .A3(new_n508_), .A4(new_n509_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n749_), .A2(new_n313_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(new_n758_), .B2(new_n487_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n760_), .B(new_n757_), .C1(new_n758_), .C2(new_n487_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1338gat));
  NAND3_X1  g563(.A1(new_n746_), .A2(new_n488_), .A3(new_n648_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n676_), .A2(new_n648_), .A3(new_n748_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n766_), .A2(new_n767_), .A3(G106gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n766_), .B2(G106gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n765_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n770_), .A2(new_n772_), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n765_), .B(new_n771_), .C1(new_n768_), .C2(new_n769_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(G1339gat));
  OR3_X1    g574(.A1(new_n614_), .A2(KEYINPUT54), .A3(new_n463_), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT54), .B1(new_n614_), .B2(new_n463_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n564_), .A2(new_n463_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n554_), .B1(new_n553_), .B2(new_n542_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n473_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n781_));
  NOR4_X1   g580(.A1(new_n781_), .A2(KEYINPUT68), .A3(new_n536_), .A4(new_n541_), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n780_), .A2(new_n782_), .A3(KEYINPUT55), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n533_), .A2(new_n538_), .A3(new_n537_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n545_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n785_), .B1(new_n786_), .B2(new_n543_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n561_), .B1(new_n783_), .B2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT56), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n544_), .A2(new_n786_), .A3(new_n555_), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n781_), .A2(new_n536_), .A3(new_n541_), .ZN(new_n792_));
  AOI22_X1  g591(.A1(KEYINPUT55), .A2(new_n792_), .B1(new_n784_), .B2(new_n545_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(KEYINPUT56), .A3(new_n561_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n779_), .B1(new_n790_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n453_), .ZN(new_n797_));
  OR3_X1    g596(.A1(new_n452_), .A2(new_n797_), .A3(new_n455_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n461_), .B1(new_n447_), .B2(new_n455_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n800_), .B1(new_n457_), .B2(new_n462_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n620_), .B1(new_n796_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  OAI211_X1 g604(.A(KEYINPUT57), .B(new_n620_), .C1(new_n796_), .C2(new_n802_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n801_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n564_), .A2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n809_), .B1(new_n790_), .B2(new_n795_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT58), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n801_), .B1(new_n556_), .B2(new_n562_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT56), .B1(new_n794_), .B2(new_n561_), .ZN(new_n814_));
  AOI211_X1 g613(.A(new_n789_), .B(new_n562_), .C1(new_n791_), .C2(new_n793_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n813_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n817_));
  AOI21_X1  g616(.A(KEYINPUT58), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n813_), .B(KEYINPUT113), .C1(new_n814_), .C2(new_n815_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n599_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT114), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n812_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT58), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n810_), .B2(KEYINPUT113), .ZN(new_n824_));
  INV_X1    g623(.A(new_n819_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n655_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT114), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n807_), .B1(new_n822_), .B2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n778_), .B1(new_n828_), .B2(new_n613_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n664_), .A2(new_n313_), .A3(new_n268_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n831_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(KEYINPUT115), .ZN(new_n833_));
  INV_X1    g632(.A(G113gat), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n463_), .A2(new_n834_), .ZN(new_n835_));
  OR2_X1    g634(.A1(new_n831_), .A2(KEYINPUT116), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT59), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n831_), .A2(KEYINPUT116), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n836_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n829_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n837_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n842_), .A2(new_n843_), .A3(new_n464_), .ZN(new_n844_));
  OAI22_X1  g643(.A1(new_n833_), .A2(new_n835_), .B1(new_n844_), .B2(new_n834_), .ZN(G1340gat));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n846_));
  INV_X1    g645(.A(new_n807_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n655_), .B(new_n821_), .C1(new_n824_), .C2(new_n825_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n811_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n820_), .A2(new_n821_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n847_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  AOI22_X1  g650(.A1(new_n851_), .A2(new_n624_), .B1(new_n777_), .B2(new_n776_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n623_), .B1(new_n852_), .B2(new_n839_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n846_), .B1(new_n853_), .B2(new_n843_), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT59), .B1(new_n852_), .B2(new_n830_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n855_), .A2(new_n841_), .A3(KEYINPUT117), .A4(new_n623_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n854_), .A2(new_n856_), .A3(G120gat), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT115), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n832_), .B(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT60), .ZN(new_n860_));
  AOI21_X1  g659(.A(G120gat), .B1(new_n623_), .B2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n861_), .B1(new_n860_), .B2(G120gat), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n859_), .A2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n857_), .A2(new_n863_), .ZN(G1341gat));
  INV_X1    g663(.A(G127gat), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n613_), .A2(new_n865_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n842_), .A2(new_n843_), .A3(new_n624_), .ZN(new_n867_));
  OAI22_X1  g666(.A1(new_n833_), .A2(new_n866_), .B1(new_n867_), .B2(new_n865_), .ZN(G1342gat));
  INV_X1    g667(.A(G134gat), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n621_), .A2(new_n869_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n842_), .A2(new_n843_), .A3(new_n599_), .ZN(new_n871_));
  OAI22_X1  g670(.A1(new_n833_), .A2(new_n870_), .B1(new_n871_), .B2(new_n869_), .ZN(G1343gat));
  NOR4_X1   g671(.A1(new_n393_), .A2(new_n313_), .A3(new_n663_), .A4(new_n269_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n829_), .A2(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n874_), .A2(new_n464_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT118), .B(G141gat), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n875_), .B(new_n876_), .ZN(G1344gat));
  NOR2_X1   g676(.A1(new_n874_), .A2(new_n567_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(new_n210_), .ZN(G1345gat));
  NOR2_X1   g678(.A1(new_n874_), .A2(new_n624_), .ZN(new_n880_));
  XOR2_X1   g679(.A(KEYINPUT61), .B(G155gat), .Z(new_n881_));
  XNOR2_X1  g680(.A(new_n880_), .B(new_n881_), .ZN(G1346gat));
  INV_X1    g681(.A(new_n874_), .ZN(new_n883_));
  AOI21_X1  g682(.A(G162gat), .B1(new_n883_), .B2(new_n621_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n655_), .A2(G162gat), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(KEYINPUT119), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n884_), .B1(new_n883_), .B2(new_n886_), .ZN(G1347gat));
  INV_X1    g686(.A(G169gat), .ZN(new_n888_));
  XOR2_X1   g687(.A(KEYINPUT120), .B(KEYINPUT62), .Z(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n424_), .A2(new_n268_), .A3(new_n648_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n829_), .A2(new_n663_), .A3(new_n463_), .A4(new_n891_), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n888_), .B(new_n890_), .C1(new_n892_), .C2(KEYINPUT22), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n890_), .B1(new_n892_), .B2(KEYINPUT22), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n892_), .A2(new_n890_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n896_), .A2(new_n888_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n894_), .B1(new_n895_), .B2(new_n897_), .ZN(G1348gat));
  NAND2_X1  g697(.A1(new_n851_), .A2(new_n624_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n370_), .B1(new_n899_), .B2(new_n778_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n900_), .A2(new_n623_), .A3(new_n891_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G176gat), .ZN(G1349gat));
  NAND4_X1  g701(.A1(new_n900_), .A2(new_n317_), .A3(new_n613_), .A4(new_n891_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n829_), .A2(new_n663_), .A3(new_n613_), .A4(new_n891_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n285_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n906_));
  AND3_X1   g705(.A1(new_n903_), .A2(new_n905_), .A3(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n903_), .B2(new_n905_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n907_), .A2(new_n908_), .ZN(G1350gat));
  NAND4_X1  g708(.A1(new_n900_), .A2(new_n299_), .A3(new_n621_), .A4(new_n891_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n900_), .A2(new_n655_), .A3(new_n891_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT122), .ZN(new_n912_));
  AND3_X1   g711(.A1(new_n911_), .A2(new_n912_), .A3(G190gat), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n912_), .B1(new_n911_), .B2(G190gat), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n910_), .B1(new_n913_), .B2(new_n914_), .ZN(G1351gat));
  NOR3_X1   g714(.A1(new_n313_), .A2(new_n393_), .A3(new_n268_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n900_), .A2(new_n463_), .A3(new_n916_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(G197gat), .ZN(G1352gat));
  AND2_X1   g717(.A1(new_n900_), .A2(new_n916_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(new_n623_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(KEYINPUT123), .B(G204gat), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n920_), .A2(new_n922_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n919_), .A2(new_n623_), .A3(new_n921_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1353gat));
  INV_X1    g724(.A(KEYINPUT124), .ZN(new_n926_));
  NOR3_X1   g725(.A1(new_n926_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n927_));
  AOI211_X1 g726(.A(new_n927_), .B(new_n624_), .C1(KEYINPUT63), .C2(G211gat), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n919_), .A2(new_n928_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n926_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n930_));
  INV_X1    g729(.A(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n929_), .A2(new_n931_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n919_), .A2(new_n930_), .A3(new_n928_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1354gat));
  NAND4_X1  g733(.A1(new_n829_), .A2(new_n663_), .A3(new_n621_), .A4(new_n916_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT125), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n935_), .B(new_n936_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(KEYINPUT126), .B(G218gat), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n599_), .A2(new_n938_), .ZN(new_n939_));
  XOR2_X1   g738(.A(new_n939_), .B(KEYINPUT127), .Z(new_n940_));
  AOI22_X1  g739(.A1(new_n937_), .A2(new_n938_), .B1(new_n919_), .B2(new_n940_), .ZN(G1355gat));
endmodule


