//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 1 1 0 1 0 0 1 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 0 1 0 1 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n630_,
    new_n631_, new_n632_, new_n633_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n806_, new_n807_,
    new_n808_, new_n810_, new_n811_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n819_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT15), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G15gat), .B(G22gat), .ZN(new_n209_));
  INV_X1    g008(.A(G1gat), .ZN(new_n210_));
  INV_X1    g009(.A(G8gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT14), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G1gat), .B(G8gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n208_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G229gat), .A2(G233gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n206_), .A2(new_n215_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n216_), .A2(new_n217_), .A3(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n206_), .B(new_n215_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(G229gat), .A3(G233gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G169gat), .B(G197gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n224_), .B(G141gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n225_), .B(KEYINPUT79), .ZN(new_n226_));
  INV_X1    g025(.A(G113gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n226_), .B(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n223_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n220_), .A2(new_n222_), .A3(new_n228_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G230gat), .A2(G233gat), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  XOR2_X1   g033(.A(G85gat), .B(G92gat), .Z(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G99gat), .A2(G106gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n239_));
  NOR2_X1   g038(.A1(G99gat), .A2(G106gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n239_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n242_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n235_), .B1(new_n238_), .B2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT8), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT9), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n235_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G85gat), .A2(G92gat), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT64), .B1(new_n248_), .B2(new_n246_), .ZN(new_n249_));
  XOR2_X1   g048(.A(KEYINPUT10), .B(G99gat), .Z(new_n250_));
  INV_X1    g049(.A(G106gat), .ZN(new_n251_));
  AOI22_X1  g050(.A1(new_n247_), .A2(new_n249_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n238_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(KEYINPUT64), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n245_), .A2(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(G57gat), .B(G64gat), .Z(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n258_), .A2(KEYINPUT11), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n258_), .A2(KEYINPUT11), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G71gat), .B(G78gat), .ZN(new_n261_));
  OR3_X1    g060(.A1(new_n259_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n258_), .A2(new_n261_), .A3(KEYINPUT11), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n256_), .A2(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n245_), .A2(new_n255_), .A3(new_n264_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n266_), .A2(KEYINPUT12), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT12), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n256_), .A2(new_n269_), .A3(new_n265_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n234_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n233_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT67), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  OR2_X1    g072(.A1(new_n272_), .A2(KEYINPUT67), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G120gat), .B(G148gat), .ZN(new_n276_));
  INV_X1    g075(.A(G204gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT5), .ZN(new_n279_));
  INV_X1    g078(.A(G176gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n275_), .A2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n273_), .A2(new_n274_), .A3(new_n281_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT13), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n283_), .A2(KEYINPUT13), .A3(new_n284_), .ZN(new_n288_));
  AND2_X1   g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT68), .ZN(new_n290_));
  NOR2_X1   g089(.A1(G141gat), .A2(G148gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT3), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT88), .ZN(new_n296_));
  NAND2_X1  g095(.A1(KEYINPUT87), .A2(KEYINPUT2), .ZN(new_n297_));
  NOR2_X1   g096(.A1(KEYINPUT87), .A2(KEYINPUT2), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G141gat), .A2(G148gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n297_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(KEYINPUT87), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n295_), .A2(new_n296_), .A3(new_n300_), .A4(new_n301_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n300_), .A2(new_n294_), .A3(new_n293_), .A4(new_n301_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT88), .ZN(new_n304_));
  OR2_X1    g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n302_), .A2(new_n304_), .A3(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT1), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n305_), .A2(new_n309_), .A3(new_n306_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n311_), .A2(new_n299_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n291_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n310_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT86), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n310_), .A2(new_n312_), .A3(KEYINPUT86), .A4(new_n313_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n308_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G127gat), .B(G134gat), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n320_), .A2(G113gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(G113gat), .ZN(new_n322_));
  AND3_X1   g121(.A1(new_n321_), .A2(G120gat), .A3(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(G120gat), .B1(new_n321_), .B2(new_n322_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n319_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n323_), .A2(new_n324_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n326_), .A2(new_n318_), .A3(new_n308_), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G225gat), .A2(G233gat), .ZN(new_n329_));
  XOR2_X1   g128(.A(new_n329_), .B(KEYINPUT96), .Z(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  AND3_X1   g130(.A1(new_n328_), .A2(KEYINPUT98), .A3(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(KEYINPUT98), .B1(new_n328_), .B2(new_n331_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n325_), .A2(KEYINPUT4), .A3(new_n327_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT95), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT95), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n325_), .A2(new_n337_), .A3(new_n327_), .A4(KEYINPUT4), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n325_), .A2(KEYINPUT4), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n336_), .A2(new_n330_), .A3(new_n338_), .A4(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n334_), .A2(new_n340_), .ZN(new_n341_));
  XOR2_X1   g140(.A(G1gat), .B(G29gat), .Z(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G57gat), .B(G85gat), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n344_), .B(new_n345_), .Z(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n341_), .A2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n346_), .B1(new_n334_), .B2(new_n340_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n319_), .A2(KEYINPUT29), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G22gat), .B(G50gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT28), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n351_), .B(new_n353_), .Z(new_n354_));
  XOR2_X1   g153(.A(G211gat), .B(G218gat), .Z(new_n355_));
  INV_X1    g154(.A(KEYINPUT89), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n356_), .B1(new_n277_), .B2(G197gat), .ZN(new_n357_));
  INV_X1    g156(.A(G197gat), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n358_), .A2(KEYINPUT89), .A3(G204gat), .ZN(new_n359_));
  AOI22_X1  g158(.A1(new_n357_), .A2(new_n359_), .B1(G197gat), .B2(new_n277_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT21), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  XOR2_X1   g161(.A(G197gat), .B(G204gat), .Z(new_n363_));
  AOI21_X1  g162(.A(new_n355_), .B1(KEYINPUT21), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n360_), .A2(new_n361_), .ZN(new_n365_));
  AOI22_X1  g164(.A1(new_n355_), .A2(new_n362_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n366_), .B1(new_n319_), .B2(KEYINPUT29), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G228gat), .A2(G233gat), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n368_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G78gat), .B(G106gat), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n372_), .B(KEYINPUT90), .Z(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n371_), .A2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n369_), .A2(new_n373_), .A3(new_n370_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n354_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT92), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n369_), .A2(KEYINPUT92), .A3(new_n373_), .A4(new_n370_), .ZN(new_n380_));
  AND3_X1   g179(.A1(new_n379_), .A2(new_n354_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT91), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n382_), .B1(new_n371_), .B2(new_n374_), .ZN(new_n383_));
  AOI211_X1 g182(.A(KEYINPUT91), .B(new_n373_), .C1(new_n369_), .C2(new_n370_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n377_), .B1(new_n381_), .B2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n326_), .B(KEYINPUT31), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G15gat), .B(G43gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(G183gat), .ZN(new_n391_));
  INV_X1    g190(.A(G190gat), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT23), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT23), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n394_), .A2(G183gat), .A3(G190gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n391_), .A2(new_n392_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  AND2_X1   g197(.A1(G169gat), .A2(G176gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT22), .B(G169gat), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n399_), .B1(new_n400_), .B2(new_n280_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n398_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n399_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT81), .ZN(new_n404_));
  NOR3_X1   g203(.A1(new_n404_), .A2(G169gat), .A3(G176gat), .ZN(new_n405_));
  INV_X1    g204(.A(G169gat), .ZN(new_n406_));
  AOI21_X1  g205(.A(KEYINPUT81), .B1(new_n406_), .B2(new_n280_), .ZN(new_n407_));
  OAI211_X1 g206(.A(KEYINPUT24), .B(new_n403_), .C1(new_n405_), .C2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT82), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT24), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n406_), .A2(new_n280_), .A3(KEYINPUT81), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n404_), .B1(G169gat), .B2(G176gat), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n410_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT82), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(new_n414_), .A3(new_n403_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n409_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT83), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n395_), .A2(new_n417_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n394_), .A2(KEYINPUT83), .A3(G183gat), .A4(G190gat), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n393_), .A3(new_n419_), .ZN(new_n420_));
  OR3_X1    g219(.A1(new_n392_), .A2(KEYINPUT80), .A3(KEYINPUT26), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT25), .B(G183gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT26), .B1(new_n392_), .B2(KEYINPUT80), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n411_), .A2(new_n412_), .A3(new_n410_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n420_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n402_), .B1(new_n416_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT84), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT84), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n429_), .B(new_n402_), .C1(new_n416_), .C2(new_n426_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G227gat), .A2(G233gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(G71gat), .ZN(new_n433_));
  XOR2_X1   g232(.A(KEYINPUT30), .B(G99gat), .Z(new_n434_));
  XOR2_X1   g233(.A(new_n433_), .B(new_n434_), .Z(new_n435_));
  NAND2_X1  g234(.A1(new_n431_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n431_), .A2(new_n435_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n390_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n438_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n440_), .A2(new_n436_), .A3(new_n389_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT85), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT85), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n439_), .A2(new_n441_), .A3(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n388_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n387_), .B1(new_n442_), .B2(KEYINPUT85), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n386_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n428_), .A2(new_n366_), .A3(new_n430_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT20), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n420_), .A2(new_n397_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT94), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT94), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n420_), .A2(new_n453_), .A3(new_n397_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n452_), .A2(new_n401_), .A3(new_n454_), .ZN(new_n455_));
  AOI211_X1 g254(.A(new_n410_), .B(new_n399_), .C1(new_n411_), .C2(new_n412_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT26), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(G190gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n392_), .A2(KEYINPUT26), .ZN(new_n459_));
  AND2_X1   g258(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n460_));
  NOR2_X1   g259(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n458_), .B(new_n459_), .C1(new_n460_), .C2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT93), .B1(new_n456_), .B2(new_n463_), .ZN(new_n464_));
  NOR3_X1   g263(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n465_), .B1(new_n393_), .B2(new_n395_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT93), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n408_), .A2(new_n467_), .A3(new_n462_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n464_), .A2(new_n466_), .A3(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n455_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n366_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n450_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n449_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G226gat), .A2(G233gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT19), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT18), .B(G64gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(G92gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G8gat), .B(G36gat), .ZN(new_n479_));
  XOR2_X1   g278(.A(new_n478_), .B(new_n479_), .Z(new_n480_));
  INV_X1    g279(.A(new_n430_), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n420_), .A2(new_n425_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n482_), .A2(new_n424_), .A3(new_n409_), .A4(new_n415_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n429_), .B1(new_n483_), .B2(new_n402_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n471_), .B1(new_n481_), .B2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n455_), .A2(new_n469_), .A3(new_n366_), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n486_), .A2(KEYINPUT20), .ZN(new_n487_));
  INV_X1    g286(.A(new_n475_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n485_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n476_), .A2(new_n480_), .A3(new_n489_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n473_), .A2(new_n475_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n487_), .A2(KEYINPUT100), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n486_), .A2(KEYINPUT20), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT100), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n492_), .A2(new_n485_), .A3(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n491_), .B1(new_n496_), .B2(new_n475_), .ZN(new_n497_));
  OAI211_X1 g296(.A(KEYINPUT27), .B(new_n490_), .C1(new_n497_), .C2(new_n480_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n480_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n366_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n500_));
  NOR3_X1   g299(.A1(new_n500_), .A2(new_n475_), .A3(new_n493_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n488_), .B1(new_n449_), .B2(new_n472_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n499_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(new_n490_), .ZN(new_n504_));
  XOR2_X1   g303(.A(KEYINPUT101), .B(KEYINPUT27), .Z(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(KEYINPUT102), .B1(new_n504_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT102), .ZN(new_n508_));
  AOI211_X1 g307(.A(new_n508_), .B(new_n505_), .C1(new_n503_), .C2(new_n490_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n498_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT103), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT103), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n498_), .B(new_n512_), .C1(new_n507_), .C2(new_n509_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n448_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n443_), .A2(new_n445_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(new_n387_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n447_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n518_), .A2(new_n510_), .A3(new_n386_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n350_), .B1(new_n514_), .B2(new_n519_), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n328_), .A2(new_n331_), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n336_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n522_));
  OAI211_X1 g321(.A(KEYINPUT33), .B(new_n521_), .C1(new_n522_), .C2(new_n330_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n347_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT33), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n341_), .A2(new_n525_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n503_), .A2(new_n490_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n334_), .A2(KEYINPUT33), .A3(new_n346_), .A4(new_n340_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n524_), .A2(new_n526_), .A3(new_n527_), .A4(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT99), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n480_), .A2(KEYINPUT32), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n476_), .A2(new_n489_), .A3(new_n531_), .ZN(new_n532_));
  OAI221_X1 g331(.A(new_n532_), .B1(new_n497_), .B2(new_n531_), .C1(new_n348_), .C2(new_n349_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n504_), .B1(new_n523_), .B2(new_n347_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT99), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n534_), .A2(new_n535_), .A3(new_n526_), .A4(new_n528_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n530_), .A2(new_n533_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n386_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n518_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n520_), .A2(new_n540_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n245_), .A2(new_n255_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n206_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n544_), .B1(new_n542_), .B2(new_n207_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G232gat), .A2(G233gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT34), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n547_), .A2(KEYINPUT35), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n545_), .A2(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n547_), .A2(KEYINPUT35), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n544_), .B(new_n551_), .C1(new_n542_), .C2(new_n207_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n549_), .A2(KEYINPUT73), .A3(new_n552_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n552_), .A2(KEYINPUT73), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(KEYINPUT72), .A2(KEYINPUT36), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT71), .B(G134gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(G162gat), .ZN(new_n558_));
  XOR2_X1   g357(.A(G190gat), .B(G218gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT72), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT36), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n560_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n555_), .A2(new_n556_), .A3(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n560_), .B(new_n562_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n553_), .A2(new_n554_), .A3(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n564_), .A2(KEYINPUT74), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(new_n568_), .A3(KEYINPUT37), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT37), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n564_), .B(new_n566_), .C1(KEYINPUT74), .C2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT16), .B(G183gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(G211gat), .ZN(new_n575_));
  XOR2_X1   g374(.A(G127gat), .B(G155gat), .Z(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT17), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT76), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G231gat), .A2(G233gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n215_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(new_n264_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n580_), .A2(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n584_), .B(KEYINPUT77), .Z(new_n585_));
  NOR3_X1   g384(.A1(new_n583_), .A2(new_n578_), .A3(new_n577_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT75), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT78), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n573_), .A2(new_n590_), .ZN(new_n591_));
  AND4_X1   g390(.A1(new_n232_), .A2(new_n290_), .A3(new_n541_), .A4(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n350_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n592_), .A2(new_n210_), .A3(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT38), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n287_), .A2(new_n288_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n596_), .A2(new_n588_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n541_), .A2(new_n567_), .A3(new_n597_), .A4(new_n232_), .ZN(new_n598_));
  OAI21_X1  g397(.A(G1gat), .B1(new_n598_), .B2(new_n350_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT104), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n595_), .A2(new_n600_), .ZN(G1324gat));
  NAND2_X1  g400(.A1(KEYINPUT105), .A2(KEYINPUT39), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n508_), .B1(new_n527_), .B2(new_n505_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n504_), .A2(KEYINPUT102), .A3(new_n506_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n512_), .B1(new_n605_), .B2(new_n498_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n513_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  OAI211_X1 g408(.A(G8gat), .B(new_n602_), .C1(new_n598_), .C2(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(KEYINPUT105), .A2(KEYINPUT39), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n592_), .A2(new_n211_), .A3(new_n608_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n610_), .A2(new_n611_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n612_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT106), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT106), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n612_), .A2(new_n613_), .A3(new_n617_), .A4(new_n614_), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n616_), .A2(KEYINPUT40), .A3(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(KEYINPUT40), .B1(new_n616_), .B2(new_n618_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(new_n620_), .ZN(G1325gat));
  INV_X1    g420(.A(G15gat), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n592_), .A2(new_n622_), .A3(new_n518_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT108), .Z(new_n624_));
  INV_X1    g423(.A(new_n518_), .ZN(new_n625_));
  OAI21_X1  g424(.A(G15gat), .B1(new_n598_), .B2(new_n625_), .ZN(new_n626_));
  XOR2_X1   g425(.A(KEYINPUT107), .B(KEYINPUT41), .Z(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n624_), .A2(new_n628_), .ZN(G1326gat));
  OAI21_X1  g428(.A(G22gat), .B1(new_n598_), .B2(new_n386_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT42), .ZN(new_n631_));
  INV_X1    g430(.A(G22gat), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n592_), .A2(new_n632_), .A3(new_n538_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(G1327gat));
  INV_X1    g433(.A(new_n232_), .ZN(new_n635_));
  NOR3_X1   g434(.A1(new_n589_), .A2(new_n596_), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n567_), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n541_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(G29gat), .B1(new_n638_), .B2(new_n593_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT110), .ZN(new_n640_));
  XNOR2_X1  g439(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n537_), .A2(new_n539_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n448_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n644_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n518_), .A2(new_n386_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n510_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n645_), .A2(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n643_), .B1(new_n649_), .B2(new_n350_), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n640_), .B(new_n642_), .C1(new_n650_), .C2(new_n572_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n572_), .B1(new_n520_), .B2(new_n540_), .ZN(new_n652_));
  OAI21_X1  g451(.A(KEYINPUT110), .B1(new_n652_), .B2(new_n641_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT43), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n651_), .A2(new_n653_), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(new_n636_), .ZN(new_n657_));
  XOR2_X1   g456(.A(KEYINPUT111), .B(KEYINPUT44), .Z(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n656_), .A2(new_n660_), .A3(new_n636_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n350_), .B1(new_n659_), .B2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n639_), .B1(new_n662_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g462(.A(G36gat), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n638_), .A2(new_n664_), .A3(new_n608_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT45), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n609_), .B1(new_n659_), .B2(new_n661_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n666_), .B1(new_n667_), .B2(new_n664_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT46), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  OAI211_X1 g469(.A(new_n666_), .B(KEYINPUT46), .C1(new_n667_), .C2(new_n664_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1329gat));
  XNOR2_X1  g471(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n656_), .A2(new_n660_), .A3(new_n636_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n658_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n676_), .B1(new_n656_), .B2(new_n636_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n518_), .B1(new_n675_), .B2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(G43gat), .ZN(new_n679_));
  INV_X1    g478(.A(G43gat), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n638_), .A2(new_n680_), .A3(new_n518_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n674_), .B1(new_n679_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n681_), .ZN(new_n683_));
  AOI211_X1 g482(.A(new_n673_), .B(new_n683_), .C1(new_n678_), .C2(G43gat), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n682_), .A2(new_n684_), .ZN(G1330gat));
  AOI21_X1  g484(.A(G50gat), .B1(new_n638_), .B2(new_n538_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n386_), .B1(new_n659_), .B2(new_n661_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n687_), .B2(G50gat), .ZN(G1331gat));
  NOR2_X1   g487(.A1(new_n289_), .A2(new_n232_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n591_), .A2(new_n541_), .A3(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n690_), .A2(new_n350_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n290_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n692_), .A2(new_n567_), .A3(new_n541_), .ZN(new_n693_));
  NOR3_X1   g492(.A1(new_n693_), .A2(new_n232_), .A3(new_n590_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(new_n593_), .ZN(new_n695_));
  MUX2_X1   g494(.A(new_n691_), .B(new_n695_), .S(G57gat), .Z(G1332gat));
  OR3_X1    g495(.A1(new_n690_), .A2(G64gat), .A3(new_n609_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n694_), .A2(new_n608_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(G64gat), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n699_), .A2(KEYINPUT48), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n699_), .A2(KEYINPUT48), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n697_), .B1(new_n700_), .B2(new_n701_), .ZN(G1333gat));
  OR3_X1    g501(.A1(new_n690_), .A2(G71gat), .A3(new_n625_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n694_), .A2(new_n518_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(G71gat), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n705_), .A2(KEYINPUT49), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n705_), .A2(KEYINPUT49), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n703_), .B1(new_n706_), .B2(new_n707_), .ZN(G1334gat));
  NAND2_X1  g507(.A1(new_n694_), .A2(new_n538_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(G78gat), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n710_), .A2(KEYINPUT50), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n710_), .A2(KEYINPUT50), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n386_), .A2(G78gat), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT113), .Z(new_n714_));
  OAI22_X1  g513(.A1(new_n711_), .A2(new_n712_), .B1(new_n690_), .B2(new_n714_), .ZN(G1335gat));
  NOR2_X1   g514(.A1(new_n290_), .A2(new_n589_), .ZN(new_n716_));
  NOR3_X1   g515(.A1(new_n650_), .A2(new_n567_), .A3(new_n232_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(G85gat), .B1(new_n718_), .B2(new_n593_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n289_), .A2(new_n589_), .A3(new_n232_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n656_), .A2(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n593_), .A2(G85gat), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT114), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n719_), .B1(new_n721_), .B2(new_n723_), .ZN(G1336gat));
  AOI21_X1  g523(.A(G92gat), .B1(new_n718_), .B2(new_n608_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n721_), .A2(G92gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n726_), .B2(new_n608_), .ZN(G1337gat));
  NAND2_X1  g526(.A1(new_n721_), .A2(new_n518_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(G99gat), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n718_), .A2(new_n250_), .A3(new_n518_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(KEYINPUT51), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT51), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n729_), .A2(new_n733_), .A3(new_n730_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(G1338gat));
  NAND3_X1  g534(.A1(new_n656_), .A2(new_n538_), .A3(new_n720_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(G106gat), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT52), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n716_), .A2(new_n717_), .A3(new_n251_), .A4(new_n538_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT115), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n736_), .A2(KEYINPUT52), .A3(G106gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n739_), .A2(new_n741_), .A3(new_n742_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g543(.A1(new_n572_), .A2(new_n289_), .A3(new_n635_), .A4(new_n589_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT54), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n284_), .A2(new_n232_), .ZN(new_n747_));
  OR2_X1    g546(.A1(KEYINPUT116), .A2(KEYINPUT55), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n271_), .A2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n268_), .A2(new_n234_), .A3(new_n270_), .ZN(new_n750_));
  XOR2_X1   g549(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n271_), .B2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n282_), .B1(new_n749_), .B2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT56), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  OAI211_X1 g554(.A(KEYINPUT56), .B(new_n282_), .C1(new_n749_), .C2(new_n752_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n747_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n221_), .A2(new_n217_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n216_), .A2(new_n219_), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n229_), .B(new_n758_), .C1(new_n759_), .C2(new_n217_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n231_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n761_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n567_), .B1(new_n757_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT57), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT57), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n765_), .B(new_n567_), .C1(new_n757_), .C2(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT58), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n755_), .A2(KEYINPUT117), .A3(new_n756_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n761_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n771_), .B(new_n284_), .C1(new_n756_), .C2(KEYINPUT117), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n770_), .B2(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n756_), .A2(KEYINPUT117), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n774_), .A2(new_n761_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n775_), .A2(new_n769_), .A3(KEYINPUT58), .A4(new_n284_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n573_), .A2(new_n773_), .A3(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n767_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n588_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n746_), .A2(new_n779_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n645_), .A2(new_n350_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n227_), .B1(new_n782_), .B2(new_n635_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT118), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  OR2_X1    g584(.A1(new_n783_), .A2(new_n784_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n778_), .A2(new_n590_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT119), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n778_), .A2(KEYINPUT119), .A3(new_n590_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n789_), .A2(new_n746_), .A3(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT59), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n792_), .A3(new_n781_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n782_), .A2(KEYINPUT59), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n232_), .A2(G113gat), .ZN(new_n797_));
  XOR2_X1   g596(.A(new_n797_), .B(KEYINPUT120), .Z(new_n798_));
  AOI22_X1  g597(.A1(new_n785_), .A2(new_n786_), .B1(new_n796_), .B2(new_n798_), .ZN(G1340gat));
  OAI21_X1  g598(.A(G120gat), .B1(new_n795_), .B2(new_n290_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n782_), .ZN(new_n801_));
  INV_X1    g600(.A(G120gat), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n802_), .B1(new_n289_), .B2(KEYINPUT60), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n801_), .B(new_n803_), .C1(KEYINPUT60), .C2(new_n802_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n800_), .A2(new_n804_), .ZN(G1341gat));
  AOI21_X1  g604(.A(G127gat), .B1(new_n801_), .B2(new_n589_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n793_), .A2(new_n794_), .A3(G127gat), .ZN(new_n807_));
  INV_X1    g606(.A(new_n588_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n806_), .B1(new_n807_), .B2(new_n808_), .ZN(G1342gat));
  AOI21_X1  g608(.A(G134gat), .B1(new_n801_), .B2(new_n637_), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n793_), .A2(new_n794_), .A3(G134gat), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n810_), .B1(new_n811_), .B2(new_n573_), .ZN(G1343gat));
  NAND3_X1  g611(.A1(new_n609_), .A2(new_n593_), .A3(new_n646_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT121), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n814_), .B1(new_n746_), .B2(new_n779_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n232_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n692_), .ZN(new_n818_));
  XOR2_X1   g617(.A(KEYINPUT122), .B(G148gat), .Z(new_n819_));
  XNOR2_X1  g618(.A(new_n818_), .B(new_n819_), .ZN(G1345gat));
  NAND2_X1  g619(.A1(new_n815_), .A2(new_n589_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(KEYINPUT61), .B(G155gat), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n821_), .B(new_n822_), .ZN(G1346gat));
  AOI21_X1  g622(.A(G162gat), .B1(new_n815_), .B2(new_n637_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n815_), .A2(G162gat), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n824_), .B1(new_n826_), .B2(new_n573_), .ZN(G1347gat));
  NOR2_X1   g626(.A1(new_n609_), .A2(new_n593_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n518_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n829_), .A2(new_n635_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n791_), .A2(new_n386_), .A3(new_n400_), .A4(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n830_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT123), .ZN(new_n833_));
  OR2_X1    g632(.A1(new_n832_), .A2(KEYINPUT123), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n791_), .A2(new_n386_), .A3(new_n833_), .A4(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT62), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n835_), .A2(new_n836_), .A3(G169gat), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n836_), .B1(new_n835_), .B2(G169gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n831_), .B1(new_n837_), .B2(new_n838_), .ZN(G1348gat));
  INV_X1    g638(.A(new_n829_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n791_), .A2(new_n596_), .A3(new_n386_), .A4(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n280_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n538_), .B1(new_n746_), .B2(new_n779_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n843_), .A2(G176gat), .A3(new_n692_), .A4(new_n840_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT124), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT124), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n842_), .A2(new_n844_), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n848_), .ZN(G1349gat));
  NOR2_X1   g648(.A1(new_n829_), .A2(new_n590_), .ZN(new_n850_));
  AOI21_X1  g649(.A(G183gat), .B1(new_n843_), .B2(new_n850_), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n791_), .A2(new_n386_), .A3(new_n840_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n588_), .A2(new_n422_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n851_), .B1(new_n852_), .B2(new_n853_), .ZN(G1350gat));
  NAND4_X1  g653(.A1(new_n791_), .A2(new_n386_), .A3(new_n573_), .A4(new_n840_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(G190gat), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n637_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n791_), .A2(new_n386_), .A3(new_n840_), .A4(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT125), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n856_), .A2(KEYINPUT125), .A3(new_n858_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1351gat));
  NAND3_X1  g662(.A1(new_n780_), .A2(new_n646_), .A3(new_n828_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT126), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n780_), .A2(KEYINPUT126), .A3(new_n646_), .A4(new_n828_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n635_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(new_n358_), .ZN(G1352gat));
  AOI21_X1  g668(.A(new_n290_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(new_n277_), .ZN(G1353gat));
  XNOR2_X1  g670(.A(KEYINPUT63), .B(G211gat), .ZN(new_n872_));
  AOI211_X1 g671(.A(new_n588_), .B(new_n872_), .C1(new_n866_), .C2(new_n867_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n866_), .A2(new_n867_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n808_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n873_), .B1(new_n875_), .B2(new_n876_), .ZN(G1354gat));
  AOI21_X1  g676(.A(G218gat), .B1(new_n874_), .B2(new_n637_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n573_), .A2(G218gat), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(KEYINPUT127), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n878_), .B1(new_n874_), .B2(new_n880_), .ZN(G1355gat));
endmodule


