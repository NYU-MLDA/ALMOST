//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 0 1 1 0 1 0 1 0 1 1 1 1 1 1 1 1 1 1 0 0 0 1 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n750_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n792_, new_n793_, new_n794_, new_n796_, new_n797_,
    new_n798_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n904_, new_n906_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_, new_n935_,
    new_n936_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n944_, new_n946_, new_n947_, new_n948_, new_n950_,
    new_n951_, new_n952_, new_n954_, new_n955_, new_n956_, new_n958_,
    new_n959_;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G64gat), .B(G92gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G226gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT19), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT20), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n215_));
  INV_X1    g014(.A(G183gat), .ZN(new_n216_));
  INV_X1    g015(.A(G190gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n214_), .A2(new_n215_), .A3(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT93), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n214_), .A2(new_n218_), .A3(KEYINPUT93), .A4(new_n215_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224_));
  INV_X1    g023(.A(G169gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT22), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT22), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(G169gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT92), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G176gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n226_), .A2(new_n228_), .A3(KEYINPUT92), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n223_), .A2(new_n224_), .A3(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n216_), .A2(KEYINPUT25), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT25), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(G183gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n217_), .A2(KEYINPUT26), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT26), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(G190gat), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n236_), .A2(new_n238_), .A3(new_n239_), .A4(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(G169gat), .A2(G176gat), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT24), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  AND3_X1   g044(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n246_));
  AOI21_X1  g045(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n225_), .A2(new_n232_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(KEYINPUT24), .A3(new_n224_), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n242_), .A2(new_n245_), .A3(new_n248_), .A4(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT91), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT25), .B(G183gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT26), .B(G190gat), .ZN(new_n254_));
  AOI22_X1  g053(.A1(new_n253_), .A2(new_n254_), .B1(new_n244_), .B2(new_n243_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n214_), .A2(new_n215_), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n257_));
  AND2_X1   g056(.A1(G169gat), .A2(G176gat), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n256_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT91), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n255_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n235_), .A2(new_n252_), .A3(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT86), .ZN(new_n264_));
  INV_X1    g063(.A(G204gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n264_), .B1(new_n265_), .B2(G197gat), .ZN(new_n266_));
  INV_X1    g065(.A(G197gat), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n267_), .A2(KEYINPUT86), .A3(G204gat), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT21), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n265_), .A2(G197gat), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n266_), .A2(new_n268_), .A3(new_n269_), .A4(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n265_), .A2(G197gat), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n267_), .A2(G204gat), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT21), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(G218gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(G211gat), .ZN(new_n276_));
  INV_X1    g075(.A(G211gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(G218gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n271_), .A2(new_n274_), .A3(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n266_), .A2(new_n270_), .A3(new_n268_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n269_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n281_), .A2(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n211_), .B1(new_n263_), .B2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT22), .B(G169gat), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n258_), .B1(new_n287_), .B2(new_n232_), .ZN(new_n288_));
  AOI22_X1  g087(.A1(new_n255_), .A2(new_n260_), .B1(new_n288_), .B2(new_n219_), .ZN(new_n289_));
  AND3_X1   g088(.A1(new_n281_), .A2(KEYINPUT87), .A3(new_n284_), .ZN(new_n290_));
  AOI21_X1  g089(.A(KEYINPUT87), .B1(new_n281_), .B2(new_n284_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n289_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n210_), .B1(new_n286_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n290_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n291_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n289_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n294_), .A2(new_n295_), .A3(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n267_), .A2(G204gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(new_n270_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n279_), .B1(KEYINPUT21), .B2(new_n299_), .ZN(new_n300_));
  AOI22_X1  g099(.A1(new_n300_), .A2(new_n271_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n235_), .A2(new_n301_), .A3(new_n252_), .A4(new_n262_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n209_), .A2(new_n211_), .ZN(new_n303_));
  AND3_X1   g102(.A1(new_n297_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n207_), .B1(new_n293_), .B2(new_n304_), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n223_), .A2(new_n224_), .A3(new_n234_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n252_), .A2(new_n262_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n285_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n308_), .A2(KEYINPUT20), .A3(new_n292_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(new_n209_), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n302_), .A2(new_n303_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n297_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n310_), .A2(new_n206_), .A3(new_n312_), .ZN(new_n313_));
  OR3_X1    g112(.A1(KEYINPUT81), .A2(G141gat), .A3(G148gat), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT81), .B1(G141gat), .B2(G148gat), .ZN(new_n315_));
  AOI22_X1  g114(.A1(new_n314_), .A2(new_n315_), .B1(G141gat), .B2(G148gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G155gat), .A2(G162gat), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT82), .B1(new_n317_), .B2(KEYINPUT1), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT82), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT1), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n319_), .A2(new_n320_), .A3(G155gat), .A4(G162gat), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n318_), .A2(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n320_), .B1(G155gat), .B2(G162gat), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n323_), .A2(new_n317_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n316_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(G141gat), .ZN(new_n326_));
  INV_X1    g125(.A(G148gat), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n326_), .A2(new_n327_), .A3(KEYINPUT3), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT3), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n329_), .B1(G141gat), .B2(G148gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n328_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT83), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G141gat), .A2(G148gat), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT2), .ZN(new_n335_));
  AOI22_X1  g134(.A1(new_n332_), .A2(new_n333_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  AND3_X1   g135(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT83), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n331_), .A2(new_n336_), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n317_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(G155gat), .A2(G162gat), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n339_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(G127gat), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n344_), .A2(G134gat), .ZN(new_n345_));
  INV_X1    g144(.A(G134gat), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n346_), .A2(G127gat), .ZN(new_n347_));
  INV_X1    g146(.A(G113gat), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n348_), .A2(G120gat), .ZN(new_n349_));
  INV_X1    g148(.A(G120gat), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n350_), .A2(G113gat), .ZN(new_n351_));
  OAI22_X1  g150(.A1(new_n345_), .A2(new_n347_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G127gat), .B(G134gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G113gat), .B(G120gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n352_), .A2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n325_), .A2(new_n343_), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT95), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n325_), .A2(new_n343_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT80), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n361_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n362_), .B1(new_n356_), .B2(new_n361_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n360_), .A2(new_n363_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n325_), .A2(new_n343_), .A3(KEYINPUT95), .A4(new_n356_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n359_), .A2(new_n364_), .A3(KEYINPUT4), .A4(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT4), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n360_), .A2(new_n363_), .A3(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n366_), .A2(new_n367_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n367_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n359_), .A2(new_n364_), .A3(new_n371_), .A4(new_n365_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G1gat), .B(G29gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(G85gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT0), .B(G57gat), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n374_), .B(new_n375_), .Z(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n370_), .A2(new_n372_), .A3(new_n377_), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n305_), .A2(new_n313_), .A3(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n366_), .A2(new_n371_), .A3(new_n369_), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n359_), .A2(new_n364_), .A3(new_n367_), .A4(new_n365_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n380_), .A2(new_n381_), .A3(new_n376_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT97), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT33), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n380_), .A2(KEYINPUT97), .A3(new_n381_), .A4(new_n376_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n384_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n377_), .A2(new_n385_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n380_), .A2(new_n388_), .A3(new_n381_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT96), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT96), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n380_), .A2(new_n388_), .A3(new_n391_), .A4(new_n381_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n379_), .A2(new_n387_), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n380_), .A2(new_n381_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n377_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n382_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n235_), .A2(new_n251_), .A3(new_n301_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT98), .B(KEYINPUT20), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NOR3_X1   g199(.A1(new_n290_), .A2(new_n291_), .A3(new_n289_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n209_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n308_), .A2(KEYINPUT20), .A3(new_n210_), .A4(new_n292_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n206_), .A2(KEYINPUT32), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n309_), .A2(new_n209_), .B1(new_n311_), .B2(new_n297_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n397_), .B(new_n406_), .C1(new_n408_), .C2(new_n405_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n394_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G78gat), .B(G106gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G228gat), .A2(G233gat), .ZN(new_n412_));
  INV_X1    g211(.A(new_n342_), .ZN(new_n413_));
  AOI22_X1  g212(.A1(new_n330_), .A2(new_n328_), .B1(new_n337_), .B2(KEYINPUT83), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n413_), .B1(new_n414_), .B2(new_n336_), .ZN(new_n415_));
  AOI22_X1  g214(.A1(new_n318_), .A2(new_n321_), .B1(new_n323_), .B2(new_n317_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n315_), .ZN(new_n417_));
  NOR3_X1   g216(.A1(KEYINPUT81), .A2(G141gat), .A3(G148gat), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n334_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n416_), .A2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT29), .B1(new_n415_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT88), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n301_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT29), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n424_), .B1(new_n325_), .B2(new_n343_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT88), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n412_), .B1(new_n423_), .B2(new_n426_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n294_), .A2(new_n421_), .A3(new_n295_), .A4(new_n412_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  OAI211_X1 g228(.A(KEYINPUT90), .B(new_n411_), .C1(new_n427_), .C2(new_n429_), .ZN(new_n430_));
  XOR2_X1   g229(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n431_));
  NOR2_X1   g230(.A1(new_n415_), .A2(new_n420_), .ZN(new_n432_));
  AOI21_X1  g231(.A(KEYINPUT84), .B1(new_n432_), .B2(new_n424_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n325_), .A2(new_n343_), .A3(KEYINPUT84), .A4(new_n424_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n431_), .B1(new_n433_), .B2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G22gat), .B(G50gat), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n325_), .A2(new_n343_), .A3(new_n424_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT84), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n431_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(new_n434_), .A3(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n436_), .A2(new_n437_), .A3(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n437_), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n440_), .A2(new_n434_), .A3(new_n441_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n441_), .B1(new_n440_), .B2(new_n434_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n444_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n412_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n285_), .B1(new_n425_), .B2(KEYINPUT88), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n421_), .A2(new_n422_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n448_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n411_), .A2(KEYINPUT90), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n451_), .A2(new_n428_), .A3(new_n452_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n430_), .A2(new_n443_), .A3(new_n447_), .A4(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n411_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n411_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n451_), .A2(new_n456_), .A3(new_n428_), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n455_), .A2(KEYINPUT89), .A3(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n447_), .A2(new_n443_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT89), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n460_), .B(new_n411_), .C1(new_n427_), .C2(new_n429_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n454_), .B1(new_n458_), .B2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n410_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n305_), .A2(new_n313_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT27), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n404_), .A2(new_n207_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT99), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n467_), .B1(new_n407_), .B2(new_n206_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n404_), .A2(KEYINPUT99), .A3(new_n207_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n471_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n397_), .ZN(new_n475_));
  NAND4_X1  g274(.A1(new_n463_), .A2(new_n468_), .A3(new_n474_), .A4(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT100), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n455_), .A2(new_n457_), .A3(KEYINPUT89), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(new_n461_), .A3(new_n459_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n397_), .B1(new_n479_), .B2(new_n454_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT100), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n480_), .A2(new_n481_), .A3(new_n468_), .A4(new_n474_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n465_), .A2(new_n477_), .A3(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G227gat), .A2(G233gat), .ZN(new_n484_));
  INV_X1    g283(.A(G15gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(G71gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(G99gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT78), .B(G43gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n289_), .B(KEYINPUT30), .Z(new_n491_));
  INV_X1    g290(.A(KEYINPUT79), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n491_), .A2(new_n492_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n490_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n495_), .B1(new_n493_), .B2(new_n490_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n363_), .B(KEYINPUT31), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n496_), .A2(new_n498_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n483_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT101), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT101), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n483_), .A2(new_n505_), .A3(new_n502_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n501_), .A2(new_n475_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n474_), .A2(new_n468_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(new_n464_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n504_), .A2(new_n506_), .A3(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(G15gat), .B(G22gat), .Z(new_n513_));
  INV_X1    g312(.A(KEYINPUT74), .ZN(new_n514_));
  INV_X1    g313(.A(G1gat), .ZN(new_n515_));
  INV_X1    g314(.A(G8gat), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT14), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n513_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n518_), .B1(new_n514_), .B2(new_n517_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G1gat), .B(G8gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT75), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n519_), .B(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G29gat), .B(G36gat), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n523_), .A2(KEYINPUT70), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(KEYINPUT70), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G43gat), .B(G50gat), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n524_), .A2(new_n525_), .A3(new_n527_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n522_), .B(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT77), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G229gat), .A2(G233gat), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT15), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n531_), .B(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(new_n522_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n531_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n522_), .A2(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n542_), .A2(new_n536_), .ZN(new_n543_));
  AOI22_X1  g342(.A1(new_n534_), .A2(new_n536_), .B1(new_n540_), .B2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G113gat), .B(G141gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G169gat), .B(G197gat), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n545_), .B(new_n546_), .Z(new_n547_));
  XNOR2_X1  g346(.A(new_n544_), .B(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n512_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT102), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G230gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT10), .B(G99gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT64), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n553_), .A2(G106gat), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT9), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G85gat), .A2(G92gat), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n555_), .B1(new_n556_), .B2(KEYINPUT65), .ZN(new_n557_));
  AND3_X1   g356(.A1(new_n556_), .A2(KEYINPUT65), .A3(new_n555_), .ZN(new_n558_));
  INV_X1    g357(.A(G85gat), .ZN(new_n559_));
  INV_X1    g358(.A(G92gat), .ZN(new_n560_));
  AOI211_X1 g359(.A(new_n557_), .B(new_n558_), .C1(new_n559_), .C2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G99gat), .A2(G106gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT6), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NOR3_X1   g363(.A1(new_n554_), .A2(new_n561_), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT66), .ZN(new_n567_));
  INV_X1    g366(.A(G99gat), .ZN(new_n568_));
  INV_X1    g367(.A(G106gat), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n567_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT7), .ZN(new_n571_));
  OAI21_X1  g370(.A(KEYINPUT66), .B1(G99gat), .B2(G106gat), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n570_), .A2(new_n571_), .A3(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT67), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n575_), .A2(new_n563_), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT8), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G85gat), .B(G92gat), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n577_), .A2(new_n578_), .A3(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n578_), .B1(new_n577_), .B2(new_n580_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n566_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G57gat), .B(G64gat), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n585_), .A2(KEYINPUT11), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(KEYINPUT11), .ZN(new_n587_));
  XOR2_X1   g386(.A(G71gat), .B(G78gat), .Z(new_n588_));
  NAND3_X1  g387(.A1(new_n586_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n587_), .A2(new_n588_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n584_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n577_), .A2(new_n580_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT8), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n565_), .B1(new_n595_), .B2(new_n581_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n596_), .A2(new_n591_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n593_), .B1(KEYINPUT68), .B2(new_n597_), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n597_), .A2(KEYINPUT68), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n551_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n584_), .A2(new_n592_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n596_), .A2(new_n591_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n601_), .A2(KEYINPUT12), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT12), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n584_), .A2(new_n604_), .A3(new_n592_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n600_), .B1(new_n551_), .B2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G120gat), .B(G148gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT5), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G176gat), .B(G204gat), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n609_), .B(new_n610_), .Z(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n607_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n607_), .A2(new_n612_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT13), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT69), .ZN(new_n618_));
  XOR2_X1   g417(.A(G190gat), .B(G218gat), .Z(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT72), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G134gat), .B(G162gat), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n620_), .B(new_n621_), .Z(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(KEYINPUT71), .B1(new_n596_), .B2(new_n538_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G232gat), .A2(G233gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT34), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n626_), .A2(KEYINPUT35), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n624_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n596_), .A2(new_n531_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n629_), .B1(new_n538_), .B2(new_n596_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n626_), .A2(KEYINPUT35), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n632_), .B1(new_n624_), .B2(new_n627_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n631_), .B1(new_n630_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT73), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n623_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT36), .B1(new_n634_), .B2(new_n623_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  AOI211_X1 g437(.A(KEYINPUT36), .B(new_n623_), .C1(new_n634_), .C2(new_n635_), .ZN(new_n639_));
  OAI21_X1  g438(.A(KEYINPUT37), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT36), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n636_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT37), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n642_), .B(new_n643_), .C1(new_n636_), .C2(new_n637_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n640_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(G231gat), .A2(G233gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n591_), .B(new_n646_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(new_n522_), .Z(new_n648_));
  XOR2_X1   g447(.A(G127gat), .B(G155gat), .Z(new_n649_));
  XNOR2_X1  g448(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(G183gat), .B(G211gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT17), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n648_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n648_), .A2(KEYINPUT17), .A3(new_n653_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n645_), .A2(new_n657_), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n550_), .A2(new_n618_), .A3(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n659_), .A2(new_n515_), .A3(new_n397_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT38), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT103), .ZN(new_n663_));
  INV_X1    g462(.A(new_n548_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n663_), .B1(new_n617_), .B2(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n615_), .B(KEYINPUT13), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n666_), .A2(KEYINPUT103), .A3(new_n548_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n657_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n638_), .A2(new_n639_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n671_), .A2(KEYINPUT104), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(KEYINPUT104), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n674_), .A2(new_n512_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n668_), .A2(new_n669_), .A3(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G1gat), .B1(new_n676_), .B2(new_n475_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n660_), .A2(new_n661_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n662_), .A2(new_n677_), .A3(new_n678_), .ZN(G1324gat));
  INV_X1    g478(.A(new_n508_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n659_), .A2(new_n516_), .A3(new_n680_), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n668_), .A2(new_n680_), .A3(new_n669_), .A4(new_n675_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT39), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n682_), .A2(new_n683_), .A3(G8gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n682_), .B2(G8gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n681_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n686_), .B(new_n687_), .Z(G1325gat));
  NAND3_X1  g487(.A1(new_n659_), .A2(new_n485_), .A3(new_n501_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT107), .Z(new_n690_));
  NAND4_X1  g489(.A1(new_n668_), .A2(new_n501_), .A3(new_n669_), .A4(new_n675_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(G15gat), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n692_), .A2(KEYINPUT41), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(KEYINPUT41), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(KEYINPUT106), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT106), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n693_), .A2(new_n697_), .A3(new_n694_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n690_), .A2(new_n696_), .A3(new_n698_), .ZN(G1326gat));
  INV_X1    g498(.A(G22gat), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n463_), .B(KEYINPUT108), .Z(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n659_), .A2(new_n700_), .A3(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(G22gat), .B1(new_n676_), .B2(new_n701_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n704_), .A2(KEYINPUT42), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(KEYINPUT42), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n703_), .B1(new_n705_), .B2(new_n706_), .ZN(G1327gat));
  NAND2_X1  g506(.A1(new_n671_), .A2(new_n657_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n617_), .A2(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n550_), .A2(new_n709_), .ZN(new_n710_));
  OR3_X1    g509(.A1(new_n710_), .A2(G29gat), .A3(new_n475_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n640_), .A2(new_n644_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n510_), .B1(new_n503_), .B2(KEYINPUT101), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n506_), .B2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n512_), .B2(new_n645_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT109), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n512_), .A2(new_n716_), .A3(new_n645_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n717_), .A2(new_n719_), .A3(new_n720_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n665_), .A2(new_n657_), .A3(new_n667_), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT44), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n723_), .A2(new_n475_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n721_), .A2(KEYINPUT44), .A3(new_n722_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n726_), .A2(KEYINPUT110), .A3(G29gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(KEYINPUT110), .B1(new_n726_), .B2(G29gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n711_), .B1(new_n727_), .B2(new_n728_), .ZN(G1328gat));
  INV_X1    g528(.A(G36gat), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n550_), .A2(new_n730_), .A3(new_n680_), .A4(new_n709_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(KEYINPUT111), .B(KEYINPUT45), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n731_), .B(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n723_), .A2(new_n508_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n735_), .A2(new_n725_), .ZN(new_n736_));
  OAI211_X1 g535(.A(KEYINPUT46), .B(new_n734_), .C1(new_n736_), .C2(new_n730_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT46), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n730_), .B1(new_n735_), .B2(new_n725_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n739_), .B2(new_n733_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n737_), .A2(new_n740_), .ZN(G1329gat));
  INV_X1    g540(.A(new_n723_), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n742_), .A2(G43gat), .A3(new_n501_), .A4(new_n725_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(KEYINPUT112), .B(G43gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n744_), .B1(new_n710_), .B2(new_n502_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g546(.A(new_n710_), .ZN(new_n748_));
  AOI21_X1  g547(.A(G50gat), .B1(new_n748_), .B2(new_n702_), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n742_), .A2(G50gat), .A3(new_n463_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n750_), .B2(new_n725_), .ZN(G1331gat));
  XNOR2_X1  g550(.A(new_n666_), .B(KEYINPUT69), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n548_), .A2(new_n657_), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n752_), .A2(new_n675_), .A3(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(G57gat), .A3(new_n397_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT114), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n755_), .A2(new_n756_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n617_), .A2(new_n658_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT113), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n548_), .B1(new_n714_), .B2(new_n506_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(G57gat), .B1(new_n763_), .B2(new_n397_), .ZN(new_n764_));
  NOR3_X1   g563(.A1(new_n757_), .A2(new_n758_), .A3(new_n764_), .ZN(G1332gat));
  INV_X1    g564(.A(G64gat), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n754_), .B2(new_n680_), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n767_), .B(KEYINPUT48), .Z(new_n768_));
  NOR2_X1   g567(.A1(new_n508_), .A2(G64gat), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT115), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n768_), .B1(new_n762_), .B2(new_n770_), .ZN(G1333gat));
  INV_X1    g570(.A(G71gat), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n772_), .B1(new_n754_), .B2(new_n501_), .ZN(new_n773_));
  XOR2_X1   g572(.A(new_n773_), .B(KEYINPUT49), .Z(new_n774_));
  NAND3_X1  g573(.A1(new_n763_), .A2(new_n772_), .A3(new_n501_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1334gat));
  OR3_X1    g575(.A1(new_n762_), .A2(G78gat), .A3(new_n701_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n754_), .A2(new_n702_), .ZN(new_n778_));
  XOR2_X1   g577(.A(KEYINPUT116), .B(KEYINPUT50), .Z(new_n779_));
  AND3_X1   g578(.A1(new_n778_), .A2(G78gat), .A3(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n778_), .B2(G78gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n777_), .B1(new_n780_), .B2(new_n781_), .ZN(G1335gat));
  NOR2_X1   g581(.A1(new_n618_), .A2(new_n708_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n761_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(G85gat), .B1(new_n785_), .B2(new_n397_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n666_), .A2(new_n548_), .A3(new_n669_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n721_), .A2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n397_), .A2(G85gat), .ZN(new_n789_));
  XOR2_X1   g588(.A(new_n789_), .B(KEYINPUT117), .Z(new_n790_));
  AOI21_X1  g589(.A(new_n786_), .B1(new_n788_), .B2(new_n790_), .ZN(G1336gat));
  OAI21_X1  g590(.A(new_n560_), .B1(new_n784_), .B2(new_n508_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(KEYINPUT118), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n508_), .A2(new_n560_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n788_), .B2(new_n794_), .ZN(G1337gat));
  OR3_X1    g594(.A1(new_n784_), .A2(new_n502_), .A3(new_n553_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n788_), .A2(new_n501_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n797_), .B2(new_n568_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g598(.A1(new_n785_), .A2(new_n569_), .A3(new_n463_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n720_), .B1(new_n718_), .B2(KEYINPUT109), .ZN(new_n802_));
  AOI211_X1 g601(.A(new_n712_), .B(new_n716_), .C1(new_n512_), .C2(new_n645_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n463_), .B(new_n787_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT119), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n721_), .A2(KEYINPUT119), .A3(new_n463_), .A4(new_n787_), .ZN(new_n807_));
  AND4_X1   g606(.A1(new_n801_), .A2(new_n806_), .A3(G106gat), .A4(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n569_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n801_), .B1(new_n809_), .B2(new_n807_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n800_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT53), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n813_), .B(new_n800_), .C1(new_n808_), .C2(new_n810_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(G1339gat));
  NAND2_X1  g614(.A1(new_n501_), .A2(new_n397_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n816_), .A2(new_n509_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n606_), .A2(new_n551_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n606_), .A2(new_n551_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT55), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n606_), .A2(new_n822_), .A3(new_n551_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n819_), .B1(new_n821_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT56), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n824_), .A2(new_n825_), .A3(new_n612_), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n606_), .A2(new_n822_), .A3(new_n551_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n822_), .B1(new_n606_), .B2(new_n551_), .ZN(new_n828_));
  OAI22_X1  g627(.A1(new_n827_), .A2(new_n828_), .B1(new_n551_), .B2(new_n606_), .ZN(new_n829_));
  AOI21_X1  g628(.A(KEYINPUT56), .B1(new_n829_), .B2(new_n611_), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n548_), .B(new_n614_), .C1(new_n826_), .C2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n544_), .A2(new_n547_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n534_), .A2(new_n535_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n542_), .A2(new_n535_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n547_), .B1(new_n540_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n832_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n615_), .A2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n671_), .B1(new_n831_), .B2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n837_), .B1(new_n607_), .B2(new_n612_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n841_), .B(KEYINPUT58), .C1(new_n826_), .C2(new_n830_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n645_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n825_), .B1(new_n824_), .B2(new_n612_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n829_), .A2(KEYINPUT56), .A3(new_n611_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT58), .B1(new_n846_), .B2(new_n841_), .ZN(new_n847_));
  OAI22_X1  g646(.A1(new_n840_), .A2(KEYINPUT57), .B1(new_n843_), .B2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n548_), .A2(new_n614_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n849_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n837_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n851_));
  OAI211_X1 g650(.A(KEYINPUT57), .B(new_n670_), .C1(new_n850_), .C2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(KEYINPUT120), .B1(new_n848_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n847_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n855_), .A2(new_n645_), .A3(new_n842_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n670_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n856_), .A2(new_n859_), .A3(new_n860_), .A4(new_n852_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n854_), .A2(new_n657_), .A3(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n666_), .A2(new_n713_), .A3(new_n753_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(KEYINPUT54), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n818_), .B1(new_n862_), .B2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n865_), .A2(new_n348_), .A3(new_n548_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n863_), .B(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n856_), .A2(new_n859_), .A3(new_n852_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n669_), .B1(new_n869_), .B2(KEYINPUT120), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n868_), .B1(new_n870_), .B2(new_n861_), .ZN(new_n871_));
  OAI21_X1  g670(.A(KEYINPUT59), .B1(new_n871_), .B2(new_n818_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n817_), .A2(KEYINPUT121), .ZN(new_n873_));
  OR2_X1    g672(.A1(new_n817_), .A2(KEYINPUT121), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT59), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  AND2_X1   g675(.A1(new_n869_), .A2(new_n657_), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n873_), .B(new_n876_), .C1(new_n877_), .C2(new_n868_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n872_), .A2(new_n548_), .A3(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n866_), .B1(new_n880_), .B2(new_n348_), .ZN(G1340gat));
  OAI211_X1 g680(.A(new_n752_), .B(new_n878_), .C1(new_n865_), .C2(new_n875_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(KEYINPUT122), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n872_), .A2(new_n884_), .A3(new_n752_), .A4(new_n878_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n883_), .A2(new_n885_), .A3(G120gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n350_), .B1(new_n666_), .B2(KEYINPUT60), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n865_), .B(new_n887_), .C1(KEYINPUT60), .C2(new_n350_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n888_), .ZN(G1341gat));
  NAND3_X1  g688(.A1(new_n865_), .A2(new_n344_), .A3(new_n669_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n872_), .A2(new_n669_), .A3(new_n878_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n890_), .B1(new_n892_), .B2(new_n344_), .ZN(G1342gat));
  INV_X1    g692(.A(new_n674_), .ZN(new_n894_));
  AOI21_X1  g693(.A(G134gat), .B1(new_n865_), .B2(new_n894_), .ZN(new_n895_));
  OR2_X1    g694(.A1(new_n895_), .A2(KEYINPUT123), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(KEYINPUT123), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n872_), .A2(new_n878_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n713_), .A2(new_n346_), .ZN(new_n899_));
  AOI22_X1  g698(.A1(new_n896_), .A2(new_n897_), .B1(new_n898_), .B2(new_n899_), .ZN(G1343gat));
  NAND2_X1  g699(.A1(new_n862_), .A2(new_n864_), .ZN(new_n901_));
  NOR4_X1   g700(.A1(new_n680_), .A2(new_n501_), .A3(new_n475_), .A4(new_n464_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n903_), .A2(new_n664_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(new_n326_), .ZN(G1344gat));
  NOR2_X1   g704(.A1(new_n903_), .A2(new_n618_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(new_n327_), .ZN(G1345gat));
  NOR2_X1   g706(.A1(new_n903_), .A2(new_n657_), .ZN(new_n908_));
  XOR2_X1   g707(.A(KEYINPUT61), .B(G155gat), .Z(new_n909_));
  XNOR2_X1  g708(.A(new_n908_), .B(new_n909_), .ZN(G1346gat));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n911_));
  INV_X1    g710(.A(G162gat), .ZN(new_n912_));
  AND2_X1   g711(.A1(new_n901_), .A2(new_n902_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n645_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n894_), .A2(new_n912_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n903_), .A2(new_n915_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n911_), .B1(new_n914_), .B2(new_n916_), .ZN(new_n917_));
  OAI21_X1  g716(.A(G162gat), .B1(new_n903_), .B2(new_n713_), .ZN(new_n918_));
  OAI211_X1 g717(.A(new_n918_), .B(KEYINPUT124), .C1(new_n903_), .C2(new_n915_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n919_), .ZN(G1347gat));
  NOR2_X1   g719(.A1(new_n877_), .A2(new_n868_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n507_), .A2(new_n508_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(new_n701_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n921_), .A2(new_n923_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n225_), .B1(new_n924_), .B2(new_n548_), .ZN(new_n925_));
  OR2_X1    g724(.A1(new_n925_), .A2(KEYINPUT62), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n548_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n927_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n928_));
  NAND4_X1  g727(.A1(new_n924_), .A2(new_n231_), .A3(new_n233_), .A4(new_n548_), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n926_), .A2(new_n928_), .A3(new_n929_), .ZN(G1348gat));
  AOI21_X1  g729(.A(G176gat), .B1(new_n924_), .B2(new_n617_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n871_), .A2(new_n463_), .ZN(new_n932_));
  AND3_X1   g731(.A1(new_n752_), .A2(G176gat), .A3(new_n922_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n931_), .B1(new_n932_), .B2(new_n933_), .ZN(G1349gat));
  NAND3_X1  g733(.A1(new_n932_), .A2(new_n669_), .A3(new_n922_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n657_), .A2(new_n253_), .ZN(new_n936_));
  AOI22_X1  g735(.A1(new_n935_), .A2(new_n216_), .B1(new_n924_), .B2(new_n936_), .ZN(G1350gat));
  NAND2_X1  g736(.A1(new_n894_), .A2(new_n254_), .ZN(new_n938_));
  XOR2_X1   g737(.A(new_n938_), .B(KEYINPUT126), .Z(new_n939_));
  NAND2_X1  g738(.A1(new_n924_), .A2(new_n939_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n924_), .A2(new_n645_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n941_), .B1(new_n942_), .B2(G190gat), .ZN(new_n943_));
  AOI211_X1 g742(.A(KEYINPUT125), .B(new_n217_), .C1(new_n924_), .C2(new_n645_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n940_), .B1(new_n943_), .B2(new_n944_), .ZN(G1351gat));
  NAND3_X1  g744(.A1(new_n502_), .A2(new_n680_), .A3(new_n480_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n871_), .A2(new_n946_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(new_n548_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(G197gat), .ZN(G1352gat));
  NOR3_X1   g748(.A1(new_n871_), .A2(new_n618_), .A3(new_n946_), .ZN(new_n950_));
  OAI21_X1  g749(.A(new_n950_), .B1(KEYINPUT127), .B2(new_n265_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(KEYINPUT127), .B(G204gat), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n951_), .B1(new_n950_), .B2(new_n952_), .ZN(G1353gat));
  NOR3_X1   g752(.A1(new_n871_), .A2(new_n657_), .A3(new_n946_), .ZN(new_n954_));
  NOR3_X1   g753(.A1(new_n954_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n955_));
  XOR2_X1   g754(.A(KEYINPUT63), .B(G211gat), .Z(new_n956_));
  AOI21_X1  g755(.A(new_n955_), .B1(new_n954_), .B2(new_n956_), .ZN(G1354gat));
  NAND3_X1  g756(.A1(new_n947_), .A2(new_n275_), .A3(new_n894_), .ZN(new_n958_));
  NOR3_X1   g757(.A1(new_n871_), .A2(new_n713_), .A3(new_n946_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n958_), .B1(new_n959_), .B2(new_n275_), .ZN(G1355gat));
endmodule


