//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 0 1 0 1 0 0 1 0 1 1 1 0 1 1 1 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n877_, new_n878_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n915_, new_n916_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT1), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT1), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G155gat), .A3(G162gat), .ZN(new_n205_));
  OR2_X1    g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n203_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n207_), .A2(new_n208_), .A3(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT83), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT86), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT84), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n215_), .B1(new_n209_), .B2(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n218_));
  AND3_X1   g017(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n219_));
  NOR3_X1   g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT85), .B1(new_n209_), .B2(new_n216_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT85), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n222_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n223_));
  NOR3_X1   g022(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n224_));
  AOI22_X1  g023(.A1(new_n221_), .A2(new_n223_), .B1(new_n224_), .B2(new_n215_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n220_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n206_), .A2(new_n202_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n214_), .B1(new_n226_), .B2(new_n228_), .ZN(new_n229_));
  AOI211_X1 g028(.A(KEYINPUT86), .B(new_n227_), .C1(new_n220_), .C2(new_n225_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n213_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT28), .B1(new_n231_), .B2(KEYINPUT29), .ZN(new_n232_));
  INV_X1    g031(.A(G50gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n226_), .A2(new_n228_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT86), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n226_), .A2(new_n214_), .A3(new_n228_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT28), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT29), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .A4(new_n213_), .ZN(new_n240_));
  AND3_X1   g039(.A1(new_n232_), .A2(new_n233_), .A3(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n233_), .B1(new_n232_), .B2(new_n240_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G78gat), .B(G106gat), .ZN(new_n244_));
  INV_X1    g043(.A(G22gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n231_), .A2(KEYINPUT29), .ZN(new_n247_));
  XOR2_X1   g046(.A(G211gat), .B(G218gat), .Z(new_n248_));
  INV_X1    g047(.A(G197gat), .ZN(new_n249_));
  NOR2_X1   g048(.A1(KEYINPUT87), .A2(G204gat), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(KEYINPUT87), .A2(G204gat), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n249_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n249_), .A2(G204gat), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  OAI211_X1 g054(.A(KEYINPUT21), .B(new_n248_), .C1(new_n253_), .C2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT88), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G197gat), .A2(G204gat), .ZN(new_n259_));
  INV_X1    g058(.A(new_n252_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n260_), .A2(new_n250_), .ZN(new_n261_));
  OAI211_X1 g060(.A(KEYINPUT21), .B(new_n259_), .C1(new_n261_), .C2(G197gat), .ZN(new_n262_));
  OAI21_X1  g061(.A(G197gat), .B1(new_n260_), .B2(new_n250_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT21), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(new_n264_), .A3(new_n254_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n248_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n262_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n264_), .B1(new_n263_), .B2(new_n254_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n268_), .A2(KEYINPUT88), .A3(new_n248_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n258_), .A2(new_n267_), .A3(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT89), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n258_), .A2(new_n267_), .A3(new_n269_), .A4(KEYINPUT89), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(G228gat), .ZN(new_n275_));
  INV_X1    g074(.A(G233gat), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  AND3_X1   g077(.A1(new_n247_), .A2(new_n274_), .A3(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n278_), .B1(new_n247_), .B2(new_n270_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n246_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n247_), .A2(new_n270_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(new_n277_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n247_), .A2(new_n274_), .A3(new_n278_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n246_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n243_), .A2(new_n281_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n242_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n232_), .A2(new_n240_), .A3(new_n233_), .ZN(new_n289_));
  AOI22_X1  g088(.A1(new_n281_), .A2(new_n286_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n287_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT23), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n293_), .B1(G183gat), .B2(G190gat), .ZN(new_n294_));
  INV_X1    g093(.A(G169gat), .ZN(new_n295_));
  INV_X1    g094(.A(G176gat), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT22), .B(G169gat), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n299_), .A2(KEYINPUT79), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT79), .B1(new_n295_), .B2(KEYINPUT22), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n296_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n294_), .B(new_n298_), .C1(new_n300_), .C2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(G169gat), .A2(G176gat), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT24), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n293_), .A2(new_n306_), .ZN(new_n307_));
  NOR3_X1   g106(.A1(new_n297_), .A2(new_n305_), .A3(new_n304_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  OR2_X1    g108(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT26), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT78), .B1(new_n313_), .B2(G190gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT26), .B(G190gat), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n312_), .B(new_n314_), .C1(new_n315_), .C2(KEYINPUT78), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n307_), .A2(new_n309_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n303_), .A2(new_n317_), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n318_), .A2(G227gat), .A3(G233gat), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n318_), .B1(G227gat), .B2(G233gat), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G127gat), .B(G134gat), .ZN(new_n322_));
  INV_X1    g121(.A(G113gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(G120gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n321_), .A2(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n319_), .A2(new_n320_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n326_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G15gat), .B(G43gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT82), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(G71gat), .B(G99gat), .Z(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT81), .B(KEYINPUT30), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n334_), .B(new_n337_), .ZN(new_n338_));
  AND3_X1   g137(.A1(new_n327_), .A2(new_n330_), .A3(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n338_), .B1(new_n327_), .B2(new_n330_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n291_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n231_), .A2(new_n329_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n326_), .B(new_n213_), .C1(new_n229_), .C2(new_n230_), .ZN(new_n344_));
  AND3_X1   g143(.A1(new_n343_), .A2(KEYINPUT4), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT4), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n231_), .A2(new_n329_), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G225gat), .A2(G233gat), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n347_), .A2(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT92), .B1(new_n345_), .B2(new_n350_), .ZN(new_n351_));
  XOR2_X1   g150(.A(G57gat), .B(G85gat), .Z(new_n352_));
  XNOR2_X1  g151(.A(G1gat), .B(G29gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n355_));
  XOR2_X1   g154(.A(new_n354_), .B(new_n355_), .Z(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n343_), .A2(new_n344_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(new_n348_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n343_), .A2(KEYINPUT4), .A3(new_n344_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT92), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n360_), .A2(new_n361_), .A3(new_n349_), .A4(new_n347_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n351_), .A2(new_n357_), .A3(new_n359_), .A4(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT33), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT94), .ZN(new_n366_));
  INV_X1    g165(.A(new_n363_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT33), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n312_), .A2(KEYINPUT90), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT90), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n310_), .A2(new_n370_), .A3(new_n311_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n315_), .ZN(new_n373_));
  OAI211_X1 g172(.A(KEYINPUT91), .B(new_n309_), .C1(new_n372_), .C2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT91), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n373_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n375_), .B1(new_n376_), .B2(new_n308_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n374_), .A2(new_n307_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n299_), .A2(new_n296_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n294_), .A2(new_n298_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  OR2_X1    g180(.A1(new_n381_), .A2(new_n270_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT20), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n383_), .B1(new_n274_), .B2(new_n318_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G226gat), .A2(G233gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT19), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n385_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G8gat), .B(G36gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT18), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(G64gat), .ZN(new_n392_));
  INV_X1    g191(.A(G92gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n381_), .A2(new_n270_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n272_), .A2(new_n303_), .A3(new_n317_), .A4(new_n273_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n396_), .A2(new_n397_), .A3(KEYINPUT20), .A4(new_n387_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n389_), .A2(new_n395_), .A3(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n387_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n398_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n394_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n358_), .A2(new_n349_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n360_), .A2(new_n348_), .A3(new_n347_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(new_n404_), .A3(new_n356_), .ZN(new_n405_));
  AND3_X1   g204(.A1(new_n399_), .A2(new_n402_), .A3(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT94), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n363_), .A2(new_n407_), .A3(new_n364_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n366_), .A2(new_n368_), .A3(new_n406_), .A4(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n394_), .A2(KEYINPUT32), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n411_), .B1(new_n389_), .B2(new_n398_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n351_), .A2(new_n359_), .A3(new_n362_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n356_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n412_), .B1(new_n414_), .B2(new_n363_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n388_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n416_));
  AND4_X1   g215(.A1(KEYINPUT20), .A2(new_n396_), .A3(new_n388_), .A4(new_n397_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n411_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n415_), .A2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n342_), .B1(new_n409_), .B2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n341_), .B1(new_n287_), .B2(new_n290_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n327_), .A2(new_n330_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n338_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n327_), .A2(new_n330_), .A3(new_n338_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NOR3_X1   g225(.A1(new_n279_), .A2(new_n280_), .A3(new_n246_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n285_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n428_));
  OAI22_X1  g227(.A1(new_n427_), .A2(new_n428_), .B1(new_n242_), .B2(new_n241_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n243_), .A2(new_n281_), .A3(new_n286_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n426_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n421_), .A2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n395_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n402_), .A2(new_n433_), .A3(KEYINPUT27), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT95), .B(KEYINPUT27), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n435_), .B1(new_n399_), .B2(new_n402_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n414_), .A2(new_n363_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n432_), .A2(new_n437_), .A3(new_n439_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n420_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT13), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT68), .ZN(new_n443_));
  INV_X1    g242(.A(G78gat), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT66), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n445_), .A2(G71gat), .ZN(new_n446_));
  INV_X1    g245(.A(G71gat), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n447_), .A2(KEYINPUT66), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n444_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(G57gat), .ZN(new_n450_));
  INV_X1    g249(.A(G64gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT11), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G57gat), .A2(G64gat), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n447_), .A2(KEYINPUT66), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n445_), .A2(G71gat), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(new_n457_), .A3(G78gat), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n449_), .A2(new_n455_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT67), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT67), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n449_), .A2(new_n461_), .A3(new_n455_), .A4(new_n458_), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n452_), .A2(new_n454_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n463_), .A2(new_n453_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n460_), .A2(new_n462_), .A3(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n464_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n443_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n464_), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n456_), .A2(new_n457_), .A3(G78gat), .ZN(new_n469_));
  AOI21_X1  g268(.A(G78gat), .B1(new_n456_), .B2(new_n457_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n461_), .B1(new_n471_), .B2(new_n455_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n462_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n468_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n460_), .A2(new_n462_), .A3(new_n464_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(KEYINPUT68), .A3(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G99gat), .A2(G106gat), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT6), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  XOR2_X1   g279(.A(KEYINPUT10), .B(G99gat), .Z(new_n481_));
  INV_X1    g280(.A(G106gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(G85gat), .ZN(new_n484_));
  OR3_X1    g283(.A1(new_n484_), .A2(new_n393_), .A3(KEYINPUT9), .ZN(new_n485_));
  AND3_X1   g284(.A1(new_n480_), .A2(new_n483_), .A3(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(G85gat), .B(G92gat), .Z(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT9), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(G99gat), .A2(G106gat), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT7), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n487_), .B1(new_n492_), .B2(new_n479_), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n493_), .A2(KEYINPUT8), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n493_), .A2(KEYINPUT8), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n489_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n467_), .A2(new_n476_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT12), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n474_), .A2(KEYINPUT70), .A3(new_n475_), .ZN(new_n500_));
  AOI21_X1  g299(.A(KEYINPUT70), .B1(new_n474_), .B2(new_n475_), .ZN(new_n501_));
  OAI211_X1 g300(.A(KEYINPUT12), .B(new_n496_), .C1(new_n500_), .C2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n467_), .A2(new_n476_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n496_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G230gat), .A2(G233gat), .ZN(new_n506_));
  XOR2_X1   g305(.A(new_n506_), .B(KEYINPUT64), .Z(new_n507_));
  XOR2_X1   g306(.A(new_n507_), .B(KEYINPUT65), .Z(new_n508_));
  NAND4_X1  g307(.A1(new_n499_), .A2(new_n502_), .A3(new_n505_), .A4(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G120gat), .B(G148gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G176gat), .B(G204gat), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n512_), .B(new_n513_), .Z(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n497_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT69), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n505_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n503_), .A2(KEYINPUT69), .A3(new_n504_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n516_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  OAI211_X1 g319(.A(new_n509_), .B(new_n515_), .C1(new_n520_), .C2(new_n508_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n508_), .ZN(new_n523_));
  AOI21_X1  g322(.A(KEYINPUT69), .B1(new_n503_), .B2(new_n504_), .ZN(new_n524_));
  AOI211_X1 g323(.A(new_n517_), .B(new_n496_), .C1(new_n467_), .C2(new_n476_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n523_), .B1(new_n526_), .B2(new_n516_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n515_), .B1(new_n527_), .B2(new_n509_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n442_), .B1(new_n522_), .B2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G29gat), .B(G36gat), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n530_), .A2(G43gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(G43gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(new_n233_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n531_), .A2(G50gat), .A3(new_n532_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G15gat), .B(G22gat), .ZN(new_n537_));
  INV_X1    g336(.A(G1gat), .ZN(new_n538_));
  INV_X1    g337(.A(G8gat), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT14), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G1gat), .B(G8gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n536_), .B(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n544_), .A2(G229gat), .A3(G233gat), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT15), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n531_), .A2(G50gat), .A3(new_n532_), .ZN(new_n547_));
  AOI21_X1  g346(.A(G50gat), .B1(new_n531_), .B2(new_n532_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n546_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n534_), .A2(KEYINPUT15), .A3(new_n535_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(new_n543_), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n536_), .A2(new_n543_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G229gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT77), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n552_), .A2(new_n553_), .A3(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n545_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G113gat), .B(G141gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(new_n295_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(new_n249_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n557_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n560_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n545_), .A2(new_n556_), .A3(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n509_), .B1(new_n520_), .B2(new_n508_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(new_n514_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n566_), .A2(KEYINPUT13), .A3(new_n521_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n529_), .A2(new_n564_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n441_), .A2(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(G231gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n543_), .B(new_n571_), .ZN(new_n572_));
  OR3_X1    g371(.A1(new_n500_), .A2(new_n501_), .A3(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G127gat), .B(G155gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G183gat), .B(G211gat), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n576_), .B(new_n577_), .Z(new_n578_));
  INV_X1    g377(.A(KEYINPUT17), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n572_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n573_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT76), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n583_), .ZN(new_n585_));
  AND2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n503_), .A2(new_n572_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n587_), .A2(new_n580_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n578_), .A2(new_n579_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n503_), .A2(new_n572_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n588_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n586_), .A2(new_n591_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n496_), .A2(new_n536_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G232gat), .A2(G233gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT34), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n595_), .A2(KEYINPUT35), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n551_), .A2(new_n496_), .A3(KEYINPUT73), .ZN(new_n597_));
  AOI21_X1  g396(.A(KEYINPUT73), .B1(new_n551_), .B2(new_n496_), .ZN(new_n598_));
  OAI211_X1 g397(.A(new_n593_), .B(new_n596_), .C1(new_n597_), .C2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n595_), .A2(KEYINPUT35), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n600_), .B(KEYINPUT72), .Z(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n551_), .A2(new_n496_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT73), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n551_), .A2(new_n496_), .A3(KEYINPUT73), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n601_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n607_), .A2(new_n608_), .A3(new_n593_), .A4(new_n596_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G190gat), .B(G218gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(G134gat), .ZN(new_n611_));
  INV_X1    g410(.A(G162gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT36), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n602_), .A2(new_n609_), .A3(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n613_), .B(new_n614_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n617_), .B1(new_n602_), .B2(new_n609_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n592_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n570_), .A2(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(G1gat), .B1(new_n621_), .B2(new_n439_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT74), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT37), .B1(new_n619_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT37), .ZN(new_n625_));
  NOR4_X1   g424(.A1(new_n616_), .A2(new_n618_), .A3(KEYINPUT74), .A4(new_n625_), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n627_), .A2(new_n592_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n570_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n438_), .B(KEYINPUT96), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n630_), .A2(new_n538_), .A3(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT97), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT97), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n630_), .A2(new_n635_), .A3(new_n538_), .A4(new_n631_), .ZN(new_n636_));
  AND3_X1   g435(.A1(new_n633_), .A2(new_n634_), .A3(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n634_), .B1(new_n633_), .B2(new_n636_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n622_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT98), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  OAI211_X1 g440(.A(KEYINPUT98), .B(new_n622_), .C1(new_n637_), .C2(new_n638_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1324gat));
  INV_X1    g442(.A(new_n437_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n570_), .A2(new_n644_), .A3(new_n620_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(G8gat), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT39), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n646_), .A2(KEYINPUT99), .A3(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n630_), .A2(new_n539_), .A3(new_n644_), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n647_), .A2(KEYINPUT99), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n647_), .A2(KEYINPUT99), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n645_), .A2(G8gat), .A3(new_n650_), .A4(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n648_), .A2(new_n649_), .A3(new_n652_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g453(.A(G15gat), .B1(new_n621_), .B2(new_n341_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT41), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n629_), .A2(G15gat), .A3(new_n341_), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1326gat));
  OAI21_X1  g457(.A(G22gat), .B1(new_n621_), .B2(new_n291_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT42), .ZN(new_n660_));
  INV_X1    g459(.A(new_n291_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n630_), .A2(new_n245_), .A3(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT100), .ZN(G1327gat));
  INV_X1    g463(.A(new_n592_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n619_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  OAI211_X1 g466(.A(new_n568_), .B(new_n667_), .C1(new_n420_), .C2(new_n440_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT102), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n432_), .A2(new_n437_), .A3(new_n439_), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n363_), .A2(new_n407_), .A3(new_n364_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n407_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n399_), .A2(new_n402_), .A3(new_n405_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n675_), .B1(KEYINPUT33), .B2(new_n367_), .ZN(new_n676_));
  AOI22_X1  g475(.A1(new_n674_), .A2(new_n676_), .B1(new_n415_), .B2(new_n418_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n671_), .B1(new_n677_), .B2(new_n342_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n678_), .A2(KEYINPUT102), .A3(new_n568_), .A4(new_n667_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n670_), .A2(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(G29gat), .B1(new_n680_), .B2(new_n438_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n627_), .B1(new_n420_), .B2(new_n440_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n682_), .A2(KEYINPUT101), .A3(KEYINPUT43), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT43), .B1(new_n682_), .B2(KEYINPUT101), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n568_), .B(new_n592_), .C1(new_n683_), .C2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n682_), .A2(KEYINPUT101), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n682_), .A2(KEYINPUT101), .A3(KEYINPUT43), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n692_), .A2(KEYINPUT44), .A3(new_n568_), .A4(new_n592_), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n687_), .A2(new_n693_), .A3(G29gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n681_), .B1(new_n694_), .B2(new_n631_), .ZN(G1328gat));
  NAND3_X1  g494(.A1(new_n687_), .A2(new_n693_), .A3(new_n644_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(G36gat), .ZN(new_n697_));
  INV_X1    g496(.A(G36gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n680_), .A2(new_n698_), .A3(new_n644_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(KEYINPUT103), .B(KEYINPUT104), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT45), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n699_), .B(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n697_), .A2(new_n702_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n697_), .A2(new_n702_), .A3(new_n704_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1329gat));
  INV_X1    g507(.A(KEYINPUT47), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n426_), .A2(G43gat), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n687_), .A2(new_n693_), .A3(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n670_), .A2(new_n679_), .A3(new_n426_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(KEYINPUT106), .A2(G43gat), .ZN(new_n713_));
  OR2_X1    g512(.A1(KEYINPUT106), .A2(G43gat), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n712_), .A2(new_n713_), .A3(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT107), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n712_), .A2(new_n717_), .A3(new_n713_), .A4(new_n714_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT108), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n711_), .A2(new_n719_), .A3(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n711_), .B2(new_n719_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n709_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n711_), .A2(new_n719_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT108), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n711_), .A2(new_n719_), .A3(new_n720_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n725_), .A2(KEYINPUT47), .A3(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n723_), .A2(new_n727_), .ZN(G1330gat));
  AOI21_X1  g527(.A(G50gat), .B1(new_n680_), .B2(new_n661_), .ZN(new_n729_));
  AOI211_X1 g528(.A(new_n233_), .B(new_n291_), .C1(new_n685_), .C2(new_n686_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n730_), .B2(new_n693_), .ZN(G1331gat));
  AND2_X1   g530(.A1(new_n529_), .A2(new_n567_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n441_), .A2(new_n564_), .A3(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(new_n620_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n734_), .A2(new_n450_), .A3(new_n439_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n628_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT109), .Z(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n631_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n735_), .B1(new_n738_), .B2(new_n450_), .ZN(G1332gat));
  INV_X1    g538(.A(new_n736_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n740_), .A2(new_n451_), .A3(new_n644_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G64gat), .B1(new_n734_), .B2(new_n437_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT110), .Z(new_n743_));
  AND2_X1   g542(.A1(new_n743_), .A2(KEYINPUT48), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(KEYINPUT48), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n741_), .B1(new_n744_), .B2(new_n745_), .ZN(G1333gat));
  OAI21_X1  g545(.A(G71gat), .B1(new_n734_), .B2(new_n341_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT49), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n740_), .A2(new_n447_), .A3(new_n426_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1334gat));
  OAI21_X1  g549(.A(G78gat), .B1(new_n734_), .B2(new_n291_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT50), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n740_), .A2(new_n444_), .A3(new_n661_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(G1335gat));
  NAND2_X1  g553(.A1(new_n733_), .A2(new_n667_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(G85gat), .B1(new_n756_), .B2(new_n631_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n732_), .A2(new_n564_), .A3(new_n665_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n692_), .A2(new_n758_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n439_), .A2(new_n484_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n757_), .B1(new_n759_), .B2(new_n760_), .ZN(G1336gat));
  NOR3_X1   g560(.A1(new_n755_), .A2(G92gat), .A3(new_n437_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n759_), .A2(new_n644_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(G92gat), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT111), .ZN(G1337gat));
  AND3_X1   g564(.A1(new_n756_), .A2(new_n481_), .A3(new_n426_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n759_), .A2(new_n426_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n767_), .B2(G99gat), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT51), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n769_), .A2(KEYINPUT112), .ZN(new_n770_));
  XOR2_X1   g569(.A(new_n768_), .B(new_n770_), .Z(G1338gat));
  OAI211_X1 g570(.A(new_n661_), .B(new_n758_), .C1(new_n683_), .C2(new_n684_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(G106gat), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT113), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n772_), .A2(new_n775_), .A3(G106gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n774_), .A2(KEYINPUT52), .A3(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n756_), .A2(new_n482_), .A3(new_n661_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n773_), .A2(KEYINPUT113), .A3(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n777_), .A2(new_n778_), .A3(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT53), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n777_), .A2(new_n783_), .A3(new_n778_), .A4(new_n780_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(G1339gat));
  INV_X1    g584(.A(new_n631_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n786_), .A2(new_n644_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n431_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n566_), .A2(new_n521_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n544_), .A2(new_n555_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n552_), .A2(new_n553_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n791_), .B(new_n560_), .C1(new_n792_), .C2(new_n555_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n793_), .A2(new_n563_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n790_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n499_), .A2(new_n502_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n523_), .B1(new_n526_), .B2(new_n796_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n499_), .A2(new_n502_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n798_), .A2(KEYINPUT55), .A3(new_n505_), .A4(new_n508_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n509_), .A2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n797_), .A2(new_n799_), .A3(new_n801_), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n802_), .A2(KEYINPUT56), .A3(new_n514_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT56), .B1(new_n802_), .B2(new_n514_), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n803_), .A2(new_n804_), .A3(KEYINPUT115), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n802_), .A2(KEYINPUT115), .A3(KEYINPUT56), .A4(new_n514_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n521_), .A2(new_n564_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n795_), .B1(new_n805_), .B2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n809_), .A2(KEYINPUT57), .A3(new_n666_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT57), .ZN(new_n811_));
  INV_X1    g610(.A(new_n795_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n802_), .A2(new_n514_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT56), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n802_), .A2(KEYINPUT56), .A3(new_n514_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n815_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n806_), .A2(new_n807_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n812_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n811_), .B1(new_n820_), .B2(new_n619_), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n521_), .A2(KEYINPUT116), .A3(new_n794_), .ZN(new_n822_));
  AOI21_X1  g621(.A(KEYINPUT116), .B1(new_n521_), .B2(new_n794_), .ZN(new_n823_));
  OAI22_X1  g622(.A1(new_n803_), .A2(new_n804_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT58), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  OAI221_X1 g625(.A(KEYINPUT58), .B1(new_n822_), .B2(new_n823_), .C1(new_n803_), .C2(new_n804_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n827_), .A3(new_n627_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n810_), .A2(new_n821_), .A3(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n810_), .A2(new_n821_), .A3(KEYINPUT117), .A4(new_n828_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n592_), .A3(new_n832_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n624_), .A2(new_n626_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n564_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n835_), .A2(new_n584_), .A3(new_n591_), .A4(new_n585_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n836_), .B(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n732_), .A2(new_n834_), .A3(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n839_), .B(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n789_), .B1(new_n833_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n323_), .B1(new_n844_), .B2(new_n835_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n829_), .A2(new_n592_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n842_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT59), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n847_), .A2(new_n848_), .A3(new_n788_), .A4(new_n787_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n835_), .A2(new_n323_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n849_), .B(new_n850_), .C1(new_n843_), .C2(new_n848_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n845_), .A2(new_n851_), .ZN(G1340gat));
  XNOR2_X1  g651(.A(KEYINPUT118), .B(G120gat), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(new_n732_), .B2(KEYINPUT60), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n843_), .B(new_n855_), .C1(KEYINPUT60), .C2(new_n854_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n732_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n857_), .B(new_n849_), .C1(new_n843_), .C2(new_n848_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n856_), .B1(new_n859_), .B2(new_n854_), .ZN(G1341gat));
  INV_X1    g659(.A(G127gat), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n861_), .B1(new_n844_), .B2(new_n592_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n592_), .A2(new_n861_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n849_), .B(new_n863_), .C1(new_n843_), .C2(new_n848_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n862_), .A2(new_n864_), .ZN(G1342gat));
  INV_X1    g664(.A(G134gat), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n866_), .B1(new_n844_), .B2(new_n666_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n834_), .A2(new_n866_), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n849_), .B(new_n868_), .C1(new_n843_), .C2(new_n848_), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n867_), .A2(new_n869_), .ZN(G1343gat));
  NAND2_X1  g669(.A1(new_n833_), .A2(new_n842_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n786_), .A2(new_n644_), .A3(new_n421_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  OR3_X1    g672(.A1(new_n873_), .A2(G141gat), .A3(new_n835_), .ZN(new_n874_));
  OAI21_X1  g673(.A(G141gat), .B1(new_n873_), .B2(new_n835_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(G1344gat));
  OR3_X1    g675(.A1(new_n873_), .A2(G148gat), .A3(new_n732_), .ZN(new_n877_));
  OAI21_X1  g676(.A(G148gat), .B1(new_n873_), .B2(new_n732_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(G1345gat));
  NAND3_X1  g678(.A1(new_n871_), .A2(new_n665_), .A3(new_n872_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(KEYINPUT61), .B(G155gat), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(KEYINPUT119), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n880_), .B(new_n882_), .ZN(G1346gat));
  NOR3_X1   g682(.A1(new_n873_), .A2(new_n612_), .A3(new_n834_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n873_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n619_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n884_), .B1(new_n612_), .B2(new_n886_), .ZN(G1347gat));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n841_), .B1(new_n829_), .B2(new_n592_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n786_), .A2(new_n644_), .A3(new_n788_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n889_), .A2(new_n835_), .A3(new_n890_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n888_), .B1(new_n891_), .B2(new_n295_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n890_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n847_), .A2(new_n564_), .A3(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n894_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n891_), .A2(new_n299_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n892_), .A2(new_n895_), .A3(new_n896_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n892_), .A2(new_n895_), .A3(KEYINPUT120), .A4(new_n896_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(G1348gat));
  NOR2_X1   g700(.A1(new_n889_), .A2(new_n890_), .ZN(new_n902_));
  AOI21_X1  g701(.A(G176gat), .B1(new_n902_), .B2(new_n857_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n890_), .A2(new_n732_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n871_), .A2(G176gat), .A3(new_n904_), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n905_), .A2(KEYINPUT121), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(KEYINPUT121), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n903_), .B1(new_n906_), .B2(new_n907_), .ZN(G1349gat));
  NOR3_X1   g707(.A1(new_n889_), .A2(new_n592_), .A3(new_n890_), .ZN(new_n909_));
  AND3_X1   g708(.A1(new_n909_), .A2(KEYINPUT122), .A3(new_n372_), .ZN(new_n910_));
  AOI21_X1  g709(.A(KEYINPUT122), .B1(new_n909_), .B2(new_n372_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n909_), .A2(G183gat), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n910_), .A2(new_n911_), .A3(new_n912_), .ZN(G1350gat));
  NAND3_X1  g712(.A1(new_n902_), .A2(new_n315_), .A3(new_n619_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n889_), .A2(new_n834_), .A3(new_n890_), .ZN(new_n915_));
  INV_X1    g714(.A(G190gat), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n914_), .B1(new_n915_), .B2(new_n916_), .ZN(G1351gat));
  NOR2_X1   g716(.A1(new_n421_), .A2(new_n438_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  OR2_X1    g718(.A1(new_n919_), .A2(KEYINPUT123), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(KEYINPUT123), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n920_), .A2(new_n644_), .A3(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n922_), .B1(new_n833_), .B2(new_n842_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n564_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(KEYINPUT124), .B(G197gat), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n924_), .B(new_n925_), .ZN(G1352gat));
  NAND2_X1  g725(.A1(new_n923_), .A2(new_n857_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(G204gat), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n928_), .B1(new_n261_), .B2(new_n927_), .ZN(G1353gat));
  AOI211_X1 g728(.A(KEYINPUT63), .B(G211gat), .C1(new_n923_), .C2(new_n665_), .ZN(new_n930_));
  AND2_X1   g729(.A1(new_n923_), .A2(new_n665_), .ZN(new_n931_));
  XOR2_X1   g730(.A(KEYINPUT63), .B(G211gat), .Z(new_n932_));
  AOI21_X1  g731(.A(new_n930_), .B1(new_n931_), .B2(new_n932_), .ZN(G1354gat));
  XNOR2_X1  g732(.A(KEYINPUT125), .B(G218gat), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n934_), .B1(new_n923_), .B2(new_n619_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n922_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n627_), .A2(new_n934_), .ZN(new_n937_));
  XOR2_X1   g736(.A(new_n937_), .B(KEYINPUT126), .Z(new_n938_));
  AND3_X1   g737(.A1(new_n871_), .A2(new_n936_), .A3(new_n938_), .ZN(new_n939_));
  OAI21_X1  g738(.A(KEYINPUT127), .B1(new_n935_), .B2(new_n939_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n923_), .A2(new_n938_), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT127), .ZN(new_n942_));
  AOI211_X1 g741(.A(new_n666_), .B(new_n922_), .C1(new_n833_), .C2(new_n842_), .ZN(new_n943_));
  OAI211_X1 g742(.A(new_n941_), .B(new_n942_), .C1(new_n943_), .C2(new_n934_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n940_), .A2(new_n944_), .ZN(G1355gat));
endmodule


