//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 1 1 0 1 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n642_,
    new_n643_, new_n644_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n866_, new_n868_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n902_, new_n903_, new_n905_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  OR2_X1    g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n208_));
  INV_X1    g007(.A(G141gat), .ZN(new_n209_));
  INV_X1    g008(.A(G148gat), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .A4(KEYINPUT83), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT83), .ZN(new_n212_));
  OAI22_X1  g011(.A1(new_n212_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT84), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n215_), .A2(KEYINPUT2), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n211_), .B(new_n213_), .C1(new_n214_), .C2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n214_), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n215_), .A2(KEYINPUT2), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n215_), .A2(KEYINPUT2), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n218_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n206_), .B(new_n207_), .C1(new_n217_), .C2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n209_), .A2(new_n210_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n207_), .A2(KEYINPUT1), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(new_n206_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n207_), .A2(KEYINPUT1), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n214_), .B(new_n223_), .C1(new_n225_), .C2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n222_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT92), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n205_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n222_), .A2(KEYINPUT92), .A3(new_n227_), .A4(new_n204_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n230_), .A2(KEYINPUT4), .A3(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G225gat), .A2(G233gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT93), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT4), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n228_), .A2(new_n235_), .A3(new_n205_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n232_), .A2(new_n234_), .A3(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n234_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n230_), .A2(new_n238_), .A3(new_n231_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G1gat), .B(G29gat), .ZN(new_n241_));
  INV_X1    g040(.A(G85gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT0), .B(G57gat), .ZN(new_n244_));
  XOR2_X1   g043(.A(new_n243_), .B(new_n244_), .Z(new_n245_));
  NAND2_X1  g044(.A1(new_n240_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n245_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n237_), .A2(new_n239_), .A3(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n204_), .B(KEYINPUT31), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT22), .B(G169gat), .ZN(new_n253_));
  INV_X1    g052(.A(G176gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT81), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(G169gat), .A2(G176gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G183gat), .A2(G190gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT23), .ZN(new_n260_));
  OR2_X1    g059(.A1(G183gat), .A2(G190gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n257_), .A2(new_n258_), .A3(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(G169gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(new_n254_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(KEYINPUT24), .A3(new_n258_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT80), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n265_), .A2(KEYINPUT24), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n260_), .A2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT26), .B(G190gat), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(KEYINPUT79), .A2(G183gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT25), .ZN(new_n274_));
  OAI211_X1 g073(.A(new_n268_), .B(new_n270_), .C1(new_n272_), .C2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n263_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G227gat), .A2(G233gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G71gat), .B(G99gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(G43gat), .ZN(new_n280_));
  XOR2_X1   g079(.A(KEYINPUT30), .B(G15gat), .Z(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n278_), .B(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT82), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n282_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n278_), .B(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT82), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n252_), .B1(new_n285_), .B2(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n251_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n250_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n266_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT25), .B(G183gat), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n293_), .B1(new_n271_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(new_n270_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n255_), .A2(new_n258_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n298_), .A2(KEYINPUT89), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT89), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n300_), .B1(new_n255_), .B2(new_n258_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n260_), .A2(KEYINPUT90), .A3(new_n261_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(KEYINPUT90), .B1(new_n260_), .B2(new_n261_), .ZN(new_n304_));
  OAI22_X1  g103(.A1(new_n299_), .A2(new_n301_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT91), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n298_), .B(KEYINPUT89), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT91), .ZN(new_n308_));
  INV_X1    g107(.A(new_n304_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(new_n302_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n307_), .A2(new_n308_), .A3(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n297_), .B1(new_n306_), .B2(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G197gat), .B(G204gat), .Z(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT21), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G211gat), .B(G218gat), .ZN(new_n315_));
  OR2_X1    g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n313_), .A2(KEYINPUT21), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n314_), .A2(new_n315_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n316_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n312_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT20), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G226gat), .A2(G233gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  AOI211_X1 g124(.A(new_n322_), .B(new_n325_), .C1(new_n276_), .C2(new_n319_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n321_), .A2(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT20), .B1(new_n276_), .B2(new_n319_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n305_), .A2(KEYINPUT91), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n308_), .B1(new_n307_), .B2(new_n310_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n296_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n328_), .B1(new_n331_), .B2(new_n319_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n325_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n327_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G8gat), .B(G36gat), .ZN(new_n335_));
  INV_X1    g134(.A(G92gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT18), .B(G64gat), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n337_), .B(new_n338_), .Z(new_n339_));
  NAND2_X1  g138(.A1(new_n334_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n339_), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n327_), .B(new_n341_), .C1(new_n332_), .C2(new_n333_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT95), .B(KEYINPUT27), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT27), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n263_), .A2(new_n275_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n322_), .B1(new_n346_), .B2(new_n320_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n347_), .B1(new_n312_), .B2(new_n320_), .ZN(new_n348_));
  AOI22_X1  g147(.A1(new_n348_), .A2(new_n325_), .B1(new_n321_), .B2(new_n326_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n345_), .B1(new_n349_), .B2(new_n341_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n320_), .A2(new_n296_), .A3(new_n305_), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n351_), .B(KEYINPUT20), .C1(new_n346_), .C2(new_n320_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(new_n325_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n353_), .B1(new_n348_), .B2(new_n325_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n339_), .ZN(new_n355_));
  AOI22_X1  g154(.A1(new_n343_), .A2(new_n344_), .B1(new_n350_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT86), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n228_), .A2(KEYINPUT29), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n358_), .A2(KEYINPUT85), .A3(new_n319_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n359_), .A2(G228gat), .A3(G233gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G228gat), .A2(G233gat), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n358_), .A2(KEYINPUT85), .A3(new_n319_), .A4(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G78gat), .B(G106gat), .Z(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n357_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G22gat), .B(G50gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n228_), .A2(KEYINPUT29), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT28), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n369_), .A2(new_n370_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n368_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n373_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n375_), .A2(new_n371_), .A3(new_n367_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n360_), .A2(KEYINPUT86), .A3(new_n362_), .A4(new_n364_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n363_), .A2(new_n365_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n366_), .A2(new_n377_), .A3(new_n378_), .A4(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n363_), .B1(KEYINPUT87), .B2(new_n364_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n364_), .A2(KEYINPUT87), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n360_), .A2(new_n362_), .A3(new_n382_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n381_), .A2(new_n383_), .A3(new_n376_), .A4(new_n374_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n380_), .A2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT96), .B1(new_n356_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n342_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n348_), .A2(new_n325_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n341_), .B1(new_n388_), .B2(new_n327_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n344_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n350_), .A2(new_n355_), .ZN(new_n391_));
  AND4_X1   g190(.A1(KEYINPUT96), .A2(new_n390_), .A3(new_n391_), .A4(new_n385_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n292_), .B1(new_n386_), .B2(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n289_), .A2(new_n290_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n385_), .ZN(new_n395_));
  AND4_X1   g194(.A1(new_n250_), .A2(new_n390_), .A3(new_n395_), .A4(new_n391_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n248_), .B(KEYINPUT33), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n230_), .A2(KEYINPUT94), .A3(new_n231_), .ZN(new_n398_));
  AOI21_X1  g197(.A(KEYINPUT94), .B1(new_n230_), .B2(new_n231_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n234_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n232_), .A2(new_n238_), .A3(new_n236_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n400_), .A2(new_n245_), .A3(new_n401_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n397_), .A2(new_n340_), .A3(new_n402_), .A4(new_n342_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n354_), .A2(KEYINPUT32), .A3(new_n341_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n341_), .A2(KEYINPUT32), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n349_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n404_), .A2(new_n406_), .A3(new_n249_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n395_), .B1(new_n403_), .B2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n394_), .B1(new_n396_), .B2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n393_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G230gat), .A2(G233gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(KEYINPUT64), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT65), .B(KEYINPUT9), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  OR2_X1    g214(.A1(KEYINPUT9), .A2(G92gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n336_), .A2(G85gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n242_), .A2(G92gat), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n416_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n415_), .A2(new_n419_), .ZN(new_n420_));
  XOR2_X1   g219(.A(KEYINPUT10), .B(G99gat), .Z(new_n421_));
  INV_X1    g220(.A(G106gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n414_), .A2(new_n417_), .A3(new_n418_), .A4(new_n416_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G99gat), .A2(G106gat), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT6), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n420_), .A2(new_n423_), .A3(new_n424_), .A4(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT7), .ZN(new_n431_));
  INV_X1    g230(.A(G99gat), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(new_n432_), .A3(new_n422_), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n433_), .A2(new_n427_), .A3(new_n428_), .A4(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT8), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n417_), .A2(new_n418_), .A3(KEYINPUT66), .ZN(new_n437_));
  AOI21_X1  g236(.A(KEYINPUT66), .B1(new_n417_), .B2(new_n418_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n435_), .B(new_n436_), .C1(new_n437_), .C2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT66), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n242_), .A2(G92gat), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n336_), .A2(G85gat), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n441_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n417_), .A2(new_n418_), .A3(KEYINPUT66), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n436_), .B1(new_n446_), .B2(new_n435_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n430_), .B1(new_n440_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT11), .ZN(new_n449_));
  INV_X1    g248(.A(G78gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(G71gat), .ZN(new_n451_));
  INV_X1    g250(.A(G71gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(G78gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G57gat), .A2(G64gat), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(G57gat), .A2(G64gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT67), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(G57gat), .ZN(new_n459_));
  INV_X1    g258(.A(G64gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT67), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(new_n462_), .A3(new_n455_), .ZN(new_n463_));
  AOI211_X1 g262(.A(new_n449_), .B(new_n454_), .C1(new_n458_), .C2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n458_), .A2(new_n463_), .A3(new_n449_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n454_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n458_), .A2(new_n463_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n466_), .B1(new_n467_), .B2(KEYINPUT11), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n464_), .B1(new_n465_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n448_), .A2(new_n469_), .ZN(new_n470_));
  NOR3_X1   g269(.A1(new_n456_), .A2(new_n457_), .A3(KEYINPUT67), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n462_), .B1(new_n461_), .B2(new_n455_), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT11), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(new_n454_), .A3(new_n465_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n467_), .A2(KEYINPUT11), .A3(new_n466_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n435_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT8), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n439_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n476_), .A2(new_n479_), .A3(new_n430_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n413_), .B1(new_n470_), .B2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n470_), .A2(KEYINPUT12), .A3(new_n480_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT12), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n448_), .A2(new_n483_), .A3(new_n469_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n482_), .A2(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n481_), .B1(new_n485_), .B2(new_n413_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT68), .ZN(new_n487_));
  XOR2_X1   g286(.A(G176gat), .B(G204gat), .Z(new_n488_));
  XNOR2_X1  g287(.A(G120gat), .B(G148gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT68), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n412_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n493_), .B1(new_n494_), .B2(new_n481_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n487_), .A2(new_n492_), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT70), .ZN(new_n497_));
  INV_X1    g296(.A(new_n492_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n497_), .B1(new_n486_), .B2(new_n498_), .ZN(new_n499_));
  NOR4_X1   g298(.A1(new_n494_), .A2(KEYINPUT70), .A3(new_n481_), .A4(new_n492_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n496_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n501_), .A2(KEYINPUT13), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(KEYINPUT13), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G113gat), .B(G141gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G169gat), .B(G197gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G29gat), .B(G36gat), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G43gat), .B(G50gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(G43gat), .B(G50gat), .Z(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(new_n509_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT71), .B(KEYINPUT15), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G1gat), .A2(G8gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT14), .ZN(new_n519_));
  XOR2_X1   g318(.A(KEYINPUT73), .B(G15gat), .Z(new_n520_));
  INV_X1    g319(.A(G22gat), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n519_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT73), .B(G15gat), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n523_), .A2(G22gat), .ZN(new_n524_));
  OAI21_X1  g323(.A(KEYINPUT74), .B1(new_n522_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n518_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(G1gat), .A2(G8gat), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n523_), .A2(G22gat), .B1(KEYINPUT14), .B2(new_n518_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n520_), .A2(new_n521_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT74), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n529_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n525_), .A2(new_n528_), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n528_), .B1(new_n525_), .B2(new_n532_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n517_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n525_), .A2(new_n532_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n528_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n515_), .B(KEYINPUT78), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n539_), .A2(new_n540_), .A3(new_n533_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(G229gat), .A2(G233gat), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n536_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT78), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n515_), .B(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n546_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n542_), .B1(new_n547_), .B2(new_n541_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n508_), .B1(new_n544_), .B2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n542_), .ZN(new_n550_));
  NOR3_X1   g349(.A1(new_n534_), .A2(new_n546_), .A3(new_n535_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n540_), .B1(new_n539_), .B2(new_n533_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n550_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n508_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n553_), .A2(new_n543_), .A3(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n549_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n505_), .A2(new_n557_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n410_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G190gat), .B(G218gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G134gat), .B(G162gat), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n560_), .B(new_n561_), .Z(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT36), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n517_), .A2(new_n448_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(G232gat), .A2(G233gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT34), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n564_), .B1(KEYINPUT35), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n448_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n512_), .A2(new_n514_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n567_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n566_), .A2(KEYINPUT35), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n572_), .A2(new_n573_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n563_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n567_), .A2(new_n571_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n573_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT36), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n580_), .A2(new_n581_), .A3(new_n562_), .A4(new_n574_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n577_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n563_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n584_), .B1(new_n580_), .B2(new_n574_), .ZN(new_n585_));
  OAI21_X1  g384(.A(KEYINPUT37), .B1(new_n585_), .B2(KEYINPUT72), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n583_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT72), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT37), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n577_), .B(new_n582_), .C1(new_n588_), .C2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n587_), .A2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n476_), .B(KEYINPUT75), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G231gat), .A2(G233gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n534_), .A2(new_n535_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G127gat), .B(G155gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(G211gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(KEYINPUT16), .B(G183gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT17), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n597_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n596_), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n595_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n595_), .A2(new_n604_), .ZN(new_n606_));
  XOR2_X1   g405(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n607_));
  AND2_X1   g406(.A1(new_n601_), .A2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n605_), .A2(new_n606_), .A3(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(KEYINPUT77), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT77), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n597_), .A2(new_n611_), .A3(new_n608_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n603_), .B1(new_n610_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n592_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n559_), .A2(new_n615_), .ZN(new_n616_));
  NOR3_X1   g415(.A1(new_n616_), .A2(G1gat), .A3(new_n250_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT97), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n614_), .A2(new_n583_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n559_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(new_n249_), .ZN(new_n623_));
  AOI22_X1  g422(.A1(new_n619_), .A2(KEYINPUT38), .B1(G1gat), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT98), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT38), .ZN(new_n626_));
  AND3_X1   g425(.A1(new_n618_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n625_), .B1(new_n618_), .B2(new_n626_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n624_), .B1(new_n627_), .B2(new_n628_), .ZN(G1324gat));
  OAI21_X1  g428(.A(G8gat), .B1(new_n621_), .B2(new_n356_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT39), .ZN(new_n631_));
  OR3_X1    g430(.A1(new_n616_), .A2(G8gat), .A3(new_n356_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT40), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(G1325gat));
  OAI21_X1  g434(.A(G15gat), .B1(new_n621_), .B2(new_n394_), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n636_), .A2(KEYINPUT41), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(KEYINPUT41), .ZN(new_n638_));
  OR3_X1    g437(.A1(new_n616_), .A2(G15gat), .A3(new_n394_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n637_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT99), .ZN(G1326gat));
  OAI21_X1  g440(.A(G22gat), .B1(new_n621_), .B2(new_n385_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT42), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n395_), .A2(new_n521_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n643_), .B1(new_n616_), .B2(new_n644_), .ZN(G1327gat));
  INV_X1    g444(.A(new_n583_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n613_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n559_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(G29gat), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n649_), .A2(new_n650_), .A3(new_n249_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n558_), .A2(new_n614_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n390_), .A2(new_n391_), .A3(new_n385_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT96), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n356_), .A2(KEYINPUT96), .A3(new_n385_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n291_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n289_), .A2(new_n290_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n403_), .A2(new_n407_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(new_n385_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n390_), .A2(new_n395_), .A3(new_n391_), .A4(new_n250_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n659_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n592_), .B1(new_n658_), .B2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT43), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT43), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n410_), .A2(new_n666_), .A3(new_n592_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n653_), .B1(new_n665_), .B2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n250_), .B1(new_n668_), .B2(KEYINPUT44), .ZN(new_n669_));
  INV_X1    g468(.A(new_n653_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n666_), .B1(new_n410_), .B2(new_n592_), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n587_), .A2(new_n591_), .ZN(new_n672_));
  AOI211_X1 g471(.A(KEYINPUT43), .B(new_n672_), .C1(new_n393_), .C2(new_n409_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n670_), .B1(new_n671_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n669_), .A2(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n652_), .B1(new_n677_), .B2(G29gat), .ZN(new_n678_));
  AOI211_X1 g477(.A(KEYINPUT100), .B(new_n650_), .C1(new_n669_), .C2(new_n676_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n651_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT101), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  OAI211_X1 g481(.A(KEYINPUT101), .B(new_n651_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1328gat));
  NOR3_X1   g483(.A1(new_n648_), .A2(G36gat), .A3(new_n356_), .ZN(new_n685_));
  XOR2_X1   g484(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT103), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n685_), .B(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT104), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n689_), .A2(KEYINPUT46), .ZN(new_n690_));
  INV_X1    g489(.A(G36gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n356_), .B1(new_n668_), .B2(KEYINPUT44), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n691_), .B1(new_n692_), .B2(new_n676_), .ZN(new_n693_));
  OR3_X1    g492(.A1(new_n688_), .A2(new_n690_), .A3(new_n693_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n690_), .B1(new_n688_), .B2(new_n693_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1329gat));
  NAND2_X1  g495(.A1(new_n668_), .A2(KEYINPUT44), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n697_), .A2(G43gat), .A3(new_n659_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n676_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n648_), .A2(new_n394_), .ZN(new_n700_));
  OAI22_X1  g499(.A1(new_n698_), .A2(new_n699_), .B1(G43gat), .B2(new_n700_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g501(.A(G50gat), .B1(new_n649_), .B2(new_n395_), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n697_), .A2(G50gat), .A3(new_n395_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n704_), .B2(new_n676_), .ZN(G1331gat));
  NAND2_X1  g504(.A1(new_n615_), .A2(new_n505_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n556_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n708_), .B(new_n410_), .C1(new_n707_), .C2(new_n706_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n709_), .B(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n711_), .A2(new_n459_), .A3(new_n249_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n504_), .A2(new_n556_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n410_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n620_), .ZN(new_n715_));
  OAI21_X1  g514(.A(G57gat), .B1(new_n715_), .B2(new_n250_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n712_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT107), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT107), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n712_), .A2(new_n719_), .A3(new_n716_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n720_), .ZN(G1332gat));
  INV_X1    g520(.A(new_n356_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(new_n460_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT109), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n711_), .A2(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(G64gat), .B1(new_n715_), .B2(new_n356_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(KEYINPUT108), .B(KEYINPUT48), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n726_), .B(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n725_), .A2(new_n728_), .ZN(G1333gat));
  NAND3_X1  g528(.A1(new_n711_), .A2(new_n452_), .A3(new_n659_), .ZN(new_n730_));
  OAI21_X1  g529(.A(G71gat), .B1(new_n715_), .B2(new_n394_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT49), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(G1334gat));
  NAND3_X1  g532(.A1(new_n711_), .A2(new_n450_), .A3(new_n395_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G78gat), .B1(new_n715_), .B2(new_n385_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT50), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(G1335gat));
  NAND2_X1  g536(.A1(new_n714_), .A2(new_n647_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(G85gat), .B1(new_n739_), .B2(new_n249_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n713_), .A2(new_n614_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT110), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT110), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n713_), .A2(new_n743_), .A3(new_n614_), .ZN(new_n744_));
  AOI22_X1  g543(.A1(new_n665_), .A2(new_n667_), .B1(new_n742_), .B2(new_n744_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n250_), .A2(new_n242_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n740_), .B1(new_n745_), .B2(new_n746_), .ZN(G1336gat));
  AOI21_X1  g546(.A(G92gat), .B1(new_n739_), .B2(new_n722_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n356_), .A2(new_n336_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n745_), .B2(new_n749_), .ZN(G1337gat));
  INV_X1    g549(.A(new_n745_), .ZN(new_n751_));
  OAI21_X1  g550(.A(G99gat), .B1(new_n751_), .B2(new_n394_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n659_), .A2(new_n421_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n752_), .B1(new_n738_), .B2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g554(.A1(new_n739_), .A2(new_n422_), .A3(new_n395_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n745_), .A2(new_n395_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT52), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n757_), .A2(KEYINPUT111), .A3(new_n758_), .A4(G106gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n422_), .B1(new_n745_), .B2(new_n395_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n759_), .B1(new_n758_), .B2(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(KEYINPUT111), .B1(new_n760_), .B2(new_n758_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n756_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n756_), .B(new_n764_), .C1(new_n761_), .C2(new_n762_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(G1339gat));
  INV_X1    g567(.A(KEYINPUT54), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n613_), .B(new_n557_), .C1(new_n587_), .C2(new_n591_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n769_), .B1(new_n771_), .B2(new_n504_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n505_), .A2(new_n770_), .A3(KEYINPUT54), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n556_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT113), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n556_), .B(new_n777_), .C1(new_n499_), .C2(new_n500_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n482_), .A2(new_n412_), .A3(new_n484_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n780_), .B1(new_n485_), .B2(new_n413_), .ZN(new_n781_));
  AOI211_X1 g580(.A(KEYINPUT55), .B(new_n412_), .C1(new_n482_), .C2(new_n484_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n779_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT56), .B1(new_n783_), .B2(new_n492_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n783_), .A2(KEYINPUT56), .A3(new_n492_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n776_), .B(new_n778_), .C1(new_n784_), .C2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n542_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n536_), .A2(new_n541_), .A3(new_n550_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(new_n508_), .A3(new_n789_), .ZN(new_n790_));
  AND2_X1   g589(.A1(new_n555_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n501_), .A2(KEYINPUT114), .A3(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n495_), .A2(new_n492_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n485_), .A2(new_n413_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n481_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n796_), .A3(new_n498_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT70), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n486_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n799_));
  AOI22_X1  g598(.A1(new_n794_), .A2(new_n487_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n791_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n793_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n787_), .A2(new_n792_), .A3(new_n802_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n803_), .A2(new_n646_), .ZN(new_n804_));
  OAI21_X1  g603(.A(KEYINPUT115), .B1(new_n804_), .B2(KEYINPUT57), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n785_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n783_), .A2(new_n492_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT56), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n807_), .A2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n808_), .A2(new_n806_), .A3(new_n809_), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n791_), .B(KEYINPUT116), .C1(new_n499_), .C2(new_n500_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n791_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  AOI22_X1  g615(.A1(new_n811_), .A2(new_n812_), .B1(new_n813_), .B2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n592_), .B1(new_n817_), .B2(KEYINPUT58), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n813_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n784_), .B1(new_n806_), .B2(new_n785_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n812_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n819_), .B(KEYINPUT58), .C1(new_n820_), .C2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  OR2_X1    g622(.A1(new_n818_), .A2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n803_), .A2(KEYINPUT57), .A3(new_n646_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT57), .B1(new_n803_), .B2(new_n646_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n805_), .A2(new_n824_), .A3(new_n825_), .A4(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n774_), .B1(new_n829_), .B2(new_n614_), .ZN(new_n830_));
  AOI211_X1 g629(.A(new_n250_), .B(new_n394_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n830_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(G113gat), .B1(new_n833_), .B2(new_n556_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n829_), .A2(new_n614_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n774_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n837_), .A2(new_n831_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n825_), .B1(new_n818_), .B2(new_n823_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n614_), .B1(new_n839_), .B2(new_n826_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n774_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  OAI211_X1 g641(.A(KEYINPUT118), .B(new_n614_), .C1(new_n839_), .C2(new_n826_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n832_), .A2(KEYINPUT59), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n838_), .A2(KEYINPUT59), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n556_), .A2(G113gat), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n834_), .B1(new_n846_), .B2(new_n847_), .ZN(G1340gat));
  NAND2_X1  g647(.A1(new_n846_), .A2(new_n505_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(G120gat), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n504_), .A2(KEYINPUT60), .ZN(new_n851_));
  MUX2_X1   g650(.A(new_n851_), .B(KEYINPUT60), .S(G120gat), .Z(new_n852_));
  NAND2_X1  g651(.A1(new_n833_), .A2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT119), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n853_), .B(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n850_), .A2(new_n855_), .ZN(G1341gat));
  AOI21_X1  g655(.A(G127gat), .B1(new_n833_), .B2(new_n613_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n613_), .A2(G127gat), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n857_), .B1(new_n846_), .B2(new_n858_), .ZN(G1342gat));
  AOI21_X1  g658(.A(G134gat), .B1(new_n833_), .B2(new_n583_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n592_), .A2(G134gat), .ZN(new_n861_));
  XOR2_X1   g660(.A(new_n861_), .B(KEYINPUT120), .Z(new_n862_));
  AOI21_X1  g661(.A(new_n860_), .B1(new_n846_), .B2(new_n862_), .ZN(G1343gat));
  NOR2_X1   g662(.A1(new_n830_), .A2(new_n659_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n722_), .A2(new_n250_), .A3(new_n385_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n864_), .A2(new_n556_), .A3(new_n865_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g666(.A1(new_n864_), .A2(new_n505_), .A3(new_n865_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g668(.A1(new_n864_), .A2(new_n613_), .A3(new_n865_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(KEYINPUT61), .B(G155gat), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n870_), .B(new_n871_), .ZN(G1346gat));
  NAND4_X1  g671(.A1(new_n864_), .A2(G162gat), .A3(new_n592_), .A4(new_n865_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n865_), .ZN(new_n874_));
  NOR4_X1   g673(.A1(new_n830_), .A2(new_n646_), .A3(new_n659_), .A4(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n873_), .B1(G162gat), .B2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT121), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n873_), .B(new_n878_), .C1(G162gat), .C2(new_n875_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n879_), .ZN(G1347gat));
  NOR3_X1   g679(.A1(new_n291_), .A2(new_n395_), .A3(new_n356_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  AOI211_X1 g681(.A(new_n557_), .B(new_n882_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n253_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n885_), .B(KEYINPUT62), .C1(new_n883_), .C2(new_n264_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n844_), .A2(new_n556_), .A3(new_n881_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n887_), .A2(new_n888_), .A3(G169gat), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n886_), .A2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n887_), .A2(G169gat), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n885_), .B1(new_n891_), .B2(KEYINPUT62), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n884_), .B1(new_n890_), .B2(new_n892_), .ZN(G1348gat));
  NAND2_X1  g692(.A1(new_n844_), .A2(new_n881_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n254_), .B1(new_n894_), .B2(new_n504_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(KEYINPUT123), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT123), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n897_), .B(new_n254_), .C1(new_n894_), .C2(new_n504_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n830_), .A2(new_n882_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n504_), .A2(new_n254_), .ZN(new_n900_));
  AOI22_X1  g699(.A1(new_n896_), .A2(new_n898_), .B1(new_n899_), .B2(new_n900_), .ZN(G1349gat));
  NOR3_X1   g700(.A1(new_n894_), .A2(new_n614_), .A3(new_n294_), .ZN(new_n902_));
  AOI21_X1  g701(.A(G183gat), .B1(new_n899_), .B2(new_n613_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1350gat));
  OAI21_X1  g703(.A(G190gat), .B1(new_n894_), .B2(new_n672_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n583_), .A2(new_n271_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(KEYINPUT124), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n905_), .B1(new_n894_), .B2(new_n907_), .ZN(G1351gat));
  NOR3_X1   g707(.A1(new_n356_), .A2(new_n249_), .A3(new_n385_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n864_), .A2(new_n556_), .A3(new_n909_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(G197gat), .ZN(G1352gat));
  AND2_X1   g710(.A1(new_n864_), .A2(new_n909_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n505_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(G204gat), .ZN(new_n914_));
  INV_X1    g713(.A(G204gat), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n912_), .A2(new_n915_), .A3(new_n505_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n916_), .ZN(G1353gat));
  NAND2_X1  g716(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n613_), .A2(new_n918_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(KEYINPUT125), .ZN(new_n920_));
  NAND4_X1  g719(.A1(new_n837_), .A2(new_n394_), .A3(new_n909_), .A4(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n922_), .ZN(new_n924_));
  NAND4_X1  g723(.A1(new_n864_), .A2(new_n909_), .A3(new_n924_), .A4(new_n920_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(KEYINPUT126), .B(KEYINPUT127), .ZN(new_n926_));
  AND3_X1   g725(.A1(new_n923_), .A2(new_n925_), .A3(new_n926_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n926_), .B1(new_n923_), .B2(new_n925_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n927_), .A2(new_n928_), .ZN(G1354gat));
  AOI21_X1  g728(.A(G218gat), .B1(new_n912_), .B2(new_n583_), .ZN(new_n930_));
  AND2_X1   g729(.A1(new_n592_), .A2(G218gat), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n912_), .B2(new_n931_), .ZN(G1355gat));
endmodule


