//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n777_, new_n778_, new_n779_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n793_, new_n794_, new_n795_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n933_, new_n935_, new_n936_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n965_,
    new_n966_, new_n967_, new_n969_, new_n970_, new_n971_, new_n972_,
    new_n973_, new_n975_, new_n976_, new_n977_, new_n979_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n986_, new_n987_, new_n988_;
  XOR2_X1   g000(.A(G113gat), .B(G141gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT78), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G169gat), .B(G197gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT75), .B(G15gat), .ZN(new_n207_));
  INV_X1    g006(.A(G22gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G1gat), .ZN(new_n210_));
  INV_X1    g009(.A(G8gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT14), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n209_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G1gat), .B(G8gat), .ZN(new_n214_));
  AND2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n213_), .A2(new_n214_), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G29gat), .B(G36gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(G43gat), .B(G50gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n218_), .B(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n220_), .B(KEYINPUT15), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n217_), .A2(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n215_), .A2(new_n216_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(new_n220_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G229gat), .A2(G233gat), .ZN(new_n225_));
  AND3_X1   g024(.A1(new_n222_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n220_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n217_), .A2(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n225_), .B1(new_n228_), .B2(new_n224_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n206_), .B1(new_n226_), .B2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n225_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n224_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n223_), .A2(new_n220_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n231_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n222_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(new_n235_), .A3(new_n205_), .ZN(new_n236_));
  AOI21_X1  g035(.A(KEYINPUT79), .B1(new_n230_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n230_), .A2(KEYINPUT79), .A3(new_n236_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(G127gat), .B(G134gat), .Z(new_n241_));
  XNOR2_X1  g040(.A(G113gat), .B(G120gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G71gat), .B(G99gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(G43gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G227gat), .A2(G233gat), .ZN(new_n247_));
  INV_X1    g046(.A(G15gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n246_), .B(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NOR3_X1   g051(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(KEYINPUT80), .A2(G190gat), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(KEYINPUT80), .A2(G190gat), .ZN(new_n257_));
  NOR3_X1   g056(.A1(new_n256_), .A2(new_n257_), .A3(G183gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G183gat), .A2(G190gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT23), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n254_), .B1(new_n258_), .B2(new_n263_), .ZN(new_n264_));
  XOR2_X1   g063(.A(KEYINPUT25), .B(G183gat), .Z(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT26), .B1(new_n256_), .B2(new_n257_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n265_), .B1(new_n266_), .B2(new_n268_), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n261_), .A2(new_n262_), .ZN(new_n270_));
  INV_X1    g069(.A(G169gat), .ZN(new_n271_));
  INV_X1    g070(.A(G176gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G169gat), .A2(G176gat), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(KEYINPUT24), .A3(new_n274_), .ZN(new_n275_));
  OR3_X1    g074(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n270_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n264_), .B1(new_n269_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT30), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  OAI211_X1 g079(.A(KEYINPUT30), .B(new_n264_), .C1(new_n269_), .C2(new_n277_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT81), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT81), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n281_), .A2(new_n284_), .A3(new_n280_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n250_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT31), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n283_), .A2(new_n250_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n287_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n289_), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT31), .B1(new_n291_), .B2(new_n286_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT82), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n290_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n293_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n244_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n296_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(new_n243_), .A3(new_n294_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  AND2_X1   g100(.A1(G228gat), .A2(G233gat), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n302_), .A2(KEYINPUT95), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT91), .B(KEYINPUT92), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(G22gat), .B(G50gat), .Z(new_n307_));
  INV_X1    g106(.A(KEYINPUT85), .ZN(new_n308_));
  NOR2_X1   g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT84), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT84), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(G155gat), .A3(G162gat), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT1), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n308_), .B(new_n310_), .C1(new_n315_), .C2(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n316_), .B1(new_n312_), .B2(new_n314_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT85), .B1(new_n318_), .B2(new_n309_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n315_), .A2(new_n316_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n317_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G141gat), .A2(G148gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT83), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT83), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n324_), .A2(G141gat), .A3(G148gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  OR2_X1    g125(.A1(G141gat), .A2(G148gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT89), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(KEYINPUT89), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n332_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT88), .B(KEYINPUT2), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n326_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n327_), .A2(KEYINPUT86), .ZN(new_n338_));
  NOR2_X1   g137(.A1(KEYINPUT87), .A2(KEYINPUT3), .ZN(new_n339_));
  AND2_X1   g138(.A1(KEYINPUT87), .A2(KEYINPUT3), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n338_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n327_), .A2(KEYINPUT86), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n335_), .B(new_n337_), .C1(new_n341_), .C2(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n315_), .A2(new_n309_), .ZN(new_n344_));
  AOI22_X1  g143(.A1(new_n321_), .A2(new_n329_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT29), .ZN(new_n346_));
  XOR2_X1   g145(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n345_), .A2(new_n346_), .A3(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n348_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n307_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n321_), .A2(new_n329_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n343_), .A2(new_n344_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n347_), .B1(new_n355_), .B2(KEYINPUT29), .ZN(new_n356_));
  INV_X1    g155(.A(new_n307_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n356_), .A2(new_n357_), .A3(new_n349_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n352_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(G106gat), .ZN(new_n360_));
  INV_X1    g159(.A(G78gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n355_), .A2(KEYINPUT29), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G197gat), .B(G204gat), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT21), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(G218gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(G211gat), .ZN(new_n367_));
  INV_X1    g166(.A(G211gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(G218gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(G197gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(G204gat), .ZN(new_n373_));
  INV_X1    g172(.A(G204gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(G197gat), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n373_), .A2(new_n375_), .A3(KEYINPUT93), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT93), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n377_), .A2(new_n372_), .A3(G204gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT21), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n365_), .B(new_n371_), .C1(new_n376_), .C2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n364_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT94), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n381_), .A2(new_n382_), .A3(new_n370_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n382_), .B1(new_n381_), .B2(new_n370_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n380_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n302_), .A2(KEYINPUT95), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n361_), .B1(new_n362_), .B2(new_n388_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n388_), .B(new_n361_), .C1(new_n345_), .C2(new_n346_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n360_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n345_), .A2(new_n346_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n388_), .ZN(new_n394_));
  OAI21_X1  g193(.A(G78gat), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n395_), .A2(G106gat), .A3(new_n390_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n359_), .A2(new_n392_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n359_), .B1(new_n396_), .B2(new_n392_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n306_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n392_), .A2(new_n396_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n401_), .A2(new_n352_), .A3(new_n358_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(new_n305_), .A3(new_n397_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n400_), .A2(new_n403_), .ZN(new_n404_));
  XOR2_X1   g203(.A(G8gat), .B(G36gat), .Z(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT18), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G64gat), .B(G92gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n406_), .B(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT32), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G226gat), .A2(G233gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT19), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT20), .B1(new_n386_), .B2(new_n278_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n381_), .A2(new_n370_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT94), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(new_n383_), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT96), .B1(new_n252_), .B2(new_n253_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT22), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n417_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT96), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n419_), .A3(new_n251_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(G183gat), .A2(G190gat), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n416_), .B(new_n420_), .C1(new_n263_), .C2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT25), .B(G183gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT26), .B(G190gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n425_), .A2(new_n270_), .A3(new_n275_), .A4(new_n276_), .ZN(new_n426_));
  AOI22_X1  g225(.A1(new_n415_), .A2(new_n380_), .B1(new_n422_), .B2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n411_), .B1(new_n412_), .B2(new_n427_), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n422_), .A2(new_n426_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n363_), .A2(KEYINPUT93), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(KEYINPUT21), .A3(new_n378_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n370_), .B1(new_n364_), .B2(new_n363_), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n414_), .A2(new_n383_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n411_), .B1(new_n429_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT20), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n435_), .B1(new_n386_), .B2(new_n278_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n428_), .A2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n409_), .B1(new_n438_), .B2(KEYINPUT97), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n422_), .A2(new_n426_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n386_), .A2(new_n440_), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n441_), .B(KEYINPUT20), .C1(new_n278_), .C2(new_n386_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n442_), .A2(new_n411_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n411_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT98), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n440_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n422_), .A2(KEYINPUT98), .A3(new_n426_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n446_), .A2(new_n433_), .A3(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n444_), .B1(new_n448_), .B2(new_n436_), .ZN(new_n449_));
  OR3_X1    g248(.A1(new_n443_), .A2(new_n449_), .A3(new_n409_), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n442_), .A2(new_n411_), .B1(new_n436_), .B2(new_n434_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n451_), .A2(KEYINPUT97), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n439_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G225gat), .A2(G233gat), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n244_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT4), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n454_), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n312_), .A2(new_n314_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n309_), .B1(new_n458_), .B2(KEYINPUT1), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n459_), .A2(new_n308_), .B1(new_n316_), .B2(new_n315_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n328_), .B1(new_n460_), .B2(new_n319_), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n343_), .A2(new_n344_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n243_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n353_), .A2(new_n244_), .A3(new_n354_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n463_), .A2(KEYINPUT4), .A3(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n457_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT99), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n463_), .A2(new_n464_), .A3(new_n454_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G1gat), .B(G29gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(G85gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT0), .B(G57gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .A4(new_n473_), .ZN(new_n474_));
  AOI221_X4 g273(.A(new_n243_), .B1(new_n343_), .B2(new_n344_), .C1(new_n321_), .C2(new_n329_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n475_), .A2(new_n455_), .ZN(new_n476_));
  AOI22_X1  g275(.A1(new_n465_), .A2(new_n457_), .B1(new_n476_), .B2(new_n454_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n474_), .B1(new_n477_), .B2(new_n473_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n467_), .B1(new_n477_), .B2(new_n473_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n453_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT100), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n477_), .A2(KEYINPUT33), .A3(new_n473_), .ZN(new_n482_));
  AOI21_X1  g281(.A(KEYINPUT33), .B1(new_n477_), .B2(new_n473_), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n428_), .A2(new_n408_), .A3(new_n437_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n408_), .B1(new_n428_), .B2(new_n437_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n463_), .A2(G225gat), .A3(new_n464_), .A4(G233gat), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n463_), .A2(KEYINPUT4), .A3(new_n464_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n454_), .B1(new_n463_), .B2(KEYINPUT4), .ZN(new_n489_));
  OAI211_X1 g288(.A(new_n472_), .B(new_n487_), .C1(new_n488_), .C2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n486_), .A2(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n483_), .A2(new_n491_), .ZN(new_n492_));
  AOI22_X1  g291(.A1(new_n480_), .A2(new_n481_), .B1(new_n482_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n466_), .A2(new_n468_), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT99), .B1(new_n494_), .B2(new_n472_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n472_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(new_n496_), .A3(new_n474_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n497_), .A2(KEYINPUT100), .A3(new_n453_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n404_), .B1(new_n493_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n408_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n438_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n428_), .A2(new_n437_), .A3(new_n408_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT27), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n504_), .B1(new_n451_), .B2(new_n408_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n500_), .B1(new_n443_), .B2(new_n449_), .ZN(new_n506_));
  AOI22_X1  g305(.A1(new_n503_), .A2(new_n504_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n507_), .A2(new_n495_), .A3(new_n496_), .A4(new_n474_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n508_), .B1(new_n400_), .B2(new_n403_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n301_), .B1(new_n499_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n404_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n497_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n300_), .A2(new_n511_), .A3(new_n512_), .A4(new_n507_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n240_), .B1(new_n510_), .B2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G71gat), .B(G78gat), .ZN(new_n515_));
  INV_X1    g314(.A(G57gat), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n516_), .A2(G64gat), .ZN(new_n517_));
  INV_X1    g316(.A(G64gat), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n518_), .A2(G57gat), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT70), .B1(new_n517_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(G57gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n516_), .A2(G64gat), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT70), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n521_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n520_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT11), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n515_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n521_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n523_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT11), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT72), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT71), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT72), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n525_), .A2(new_n535_), .A3(KEYINPUT11), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n533_), .A2(new_n534_), .A3(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n534_), .B1(new_n533_), .B2(new_n536_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n529_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n535_), .B1(new_n525_), .B2(KEYINPUT11), .ZN(new_n540_));
  AOI211_X1 g339(.A(KEYINPUT72), .B(new_n527_), .C1(new_n520_), .C2(new_n524_), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT71), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n533_), .A2(new_n536_), .A3(new_n534_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n542_), .A2(new_n528_), .A3(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT8), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n545_), .A2(KEYINPUT69), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT7), .ZN(new_n547_));
  INV_X1    g346(.A(G99gat), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n547_), .A2(new_n548_), .A3(new_n360_), .A4(KEYINPUT68), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT68), .ZN(new_n550_));
  OAI22_X1  g349(.A1(new_n550_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT6), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT67), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT67), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT6), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G99gat), .A2(G106gat), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  AND2_X1   g358(.A1(G99gat), .A2(G106gat), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n554_), .A2(new_n556_), .A3(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n552_), .B1(new_n559_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G85gat), .A2(G92gat), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(G85gat), .A2(G92gat), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n546_), .B1(new_n562_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n546_), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n554_), .A2(new_n556_), .A3(new_n560_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n560_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n569_), .B(new_n566_), .C1(new_n572_), .C2(new_n552_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n568_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n572_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT64), .ZN(new_n576_));
  XOR2_X1   g375(.A(KEYINPUT10), .B(G99gat), .Z(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n576_), .B1(new_n578_), .B2(G106gat), .ZN(new_n579_));
  NAND3_X1  g378(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n580_), .B1(new_n565_), .B2(KEYINPUT66), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT9), .ZN(new_n582_));
  AND3_X1   g381(.A1(new_n563_), .A2(KEYINPUT65), .A3(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(KEYINPUT65), .B1(new_n563_), .B2(new_n582_), .ZN(new_n584_));
  OAI221_X1 g383(.A(new_n581_), .B1(KEYINPUT66), .B2(new_n580_), .C1(new_n583_), .C2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n577_), .A2(KEYINPUT64), .A3(new_n360_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n575_), .A2(new_n579_), .A3(new_n585_), .A4(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n574_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n539_), .A2(new_n544_), .A3(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n588_), .B1(new_n539_), .B2(new_n544_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT12), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n589_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n542_), .A2(new_n528_), .A3(new_n543_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n528_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n593_), .A2(new_n594_), .A3(new_n591_), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n574_), .A2(KEYINPUT73), .A3(new_n587_), .ZN(new_n596_));
  AOI21_X1  g395(.A(KEYINPUT73), .B1(new_n574_), .B2(new_n587_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n595_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G230gat), .A2(G233gat), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n592_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n588_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n602_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(new_n589_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n604_), .A2(G230gat), .A3(G233gat), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n601_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G120gat), .B(G148gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT5), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G176gat), .B(G204gat), .ZN(new_n609_));
  XOR2_X1   g408(.A(new_n608_), .B(new_n609_), .Z(new_n610_));
  NAND2_X1  g409(.A1(new_n606_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n610_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n601_), .A2(new_n605_), .A3(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT13), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n611_), .A2(KEYINPUT13), .A3(new_n613_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  XOR2_X1   g418(.A(G127gat), .B(G155gat), .Z(new_n620_));
  XNOR2_X1  g419(.A(G183gat), .B(G211gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  AND2_X1   g423(.A1(G231gat), .A2(G233gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n223_), .B(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n593_), .A2(new_n594_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n626_), .A2(new_n627_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n624_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n629_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n626_), .A2(new_n627_), .ZN(new_n633_));
  OAI21_X1  g432(.A(KEYINPUT77), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  AOI22_X1  g433(.A1(new_n631_), .A2(KEYINPUT17), .B1(new_n634_), .B2(new_n624_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n634_), .A2(KEYINPUT17), .A3(new_n624_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n598_), .A2(new_n221_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(G232gat), .A2(G233gat), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT34), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(KEYINPUT74), .B(KEYINPUT35), .ZN(new_n644_));
  AOI22_X1  g443(.A1(new_n602_), .A2(new_n220_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n640_), .A2(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n643_), .A2(new_n644_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n640_), .B(new_n645_), .C1(new_n643_), .C2(new_n644_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(G190gat), .B(G218gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(G134gat), .B(G162gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT36), .Z(new_n654_));
  NAND2_X1  g453(.A1(new_n650_), .A2(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n653_), .A2(KEYINPUT36), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n648_), .A2(new_n656_), .A3(new_n649_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n658_), .A2(KEYINPUT37), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(KEYINPUT37), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  AND4_X1   g460(.A1(new_n514_), .A2(new_n619_), .A3(new_n639_), .A4(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n662_), .A2(new_n210_), .A3(new_n497_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT38), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n658_), .B(KEYINPUT101), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(new_n510_), .B2(new_n513_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n230_), .A2(new_n236_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n618_), .A2(new_n638_), .A3(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n667_), .A2(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n210_), .B1(new_n671_), .B2(new_n497_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n665_), .A2(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n673_), .B1(new_n664_), .B2(new_n663_), .ZN(G1324gat));
  INV_X1    g473(.A(new_n507_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n671_), .A2(new_n675_), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n676_), .A2(KEYINPUT102), .A3(G8gat), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT102), .B1(new_n676_), .B2(G8gat), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT39), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n677_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n678_), .A2(new_n679_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n662_), .A2(new_n211_), .A3(new_n675_), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n681_), .A2(KEYINPUT40), .A3(new_n682_), .A4(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT40), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n682_), .A2(new_n683_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n685_), .B1(new_n680_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n684_), .A2(new_n687_), .ZN(G1325gat));
  AOI21_X1  g487(.A(new_n248_), .B1(new_n671_), .B2(new_n300_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT41), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n662_), .A2(new_n248_), .A3(new_n300_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1326gat));
  AOI21_X1  g491(.A(new_n208_), .B1(new_n671_), .B2(new_n404_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT42), .Z(new_n694_));
  NAND3_X1  g493(.A1(new_n662_), .A2(new_n208_), .A3(new_n404_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1327gat));
  NAND2_X1  g495(.A1(new_n666_), .A2(new_n638_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n697_), .A2(new_n618_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n514_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(G29gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(new_n700_), .A3(new_n497_), .ZN(new_n701_));
  NOR3_X1   g500(.A1(new_n639_), .A2(new_n669_), .A3(new_n618_), .ZN(new_n702_));
  AOI211_X1 g501(.A(KEYINPUT43), .B(new_n661_), .C1(new_n510_), .C2(new_n513_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n480_), .A2(new_n481_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n492_), .A2(new_n482_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n705_), .A2(new_n498_), .A3(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n509_), .B1(new_n707_), .B2(new_n511_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n513_), .B1(new_n708_), .B2(new_n300_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n661_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n704_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n702_), .B1(new_n703_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(KEYINPUT44), .B1(new_n712_), .B2(KEYINPUT103), .ZN(new_n715_));
  INV_X1    g514(.A(new_n702_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n709_), .A2(new_n710_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT43), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n709_), .A2(new_n704_), .A3(new_n710_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n716_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT103), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n714_), .B1(new_n715_), .B2(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n723_), .A2(KEYINPUT104), .A3(new_n497_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(G29gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(KEYINPUT104), .B1(new_n723_), .B2(new_n497_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n701_), .B1(new_n725_), .B2(new_n726_), .ZN(G1328gat));
  INV_X1    g526(.A(KEYINPUT46), .ZN(new_n728_));
  INV_X1    g527(.A(G36gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n729_), .B1(new_n723_), .B2(new_n675_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n507_), .B(KEYINPUT105), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n699_), .A2(new_n729_), .A3(new_n732_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT45), .Z(new_n734_));
  OAI21_X1  g533(.A(new_n728_), .B1(new_n730_), .B2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n720_), .A2(KEYINPUT44), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n713_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n712_), .A2(KEYINPUT103), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n675_), .B(new_n736_), .C1(new_n737_), .C2(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(G36gat), .ZN(new_n740_));
  INV_X1    g539(.A(new_n734_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n740_), .A2(new_n741_), .A3(KEYINPUT46), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n735_), .A2(new_n742_), .ZN(G1329gat));
  AOI21_X1  g542(.A(G43gat), .B1(new_n699_), .B2(new_n300_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n300_), .A2(G43gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n723_), .B2(new_n745_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n747_), .ZN(new_n749_));
  AOI211_X1 g548(.A(new_n744_), .B(new_n749_), .C1(new_n723_), .C2(new_n745_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n748_), .A2(new_n750_), .ZN(G1330gat));
  AOI21_X1  g550(.A(G50gat), .B1(new_n699_), .B2(new_n404_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n404_), .A2(G50gat), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n723_), .B2(new_n753_), .ZN(G1331gat));
  OAI21_X1  g553(.A(new_n240_), .B1(new_n635_), .B2(new_n637_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n619_), .A2(new_n755_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n667_), .A2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(G57gat), .B1(new_n758_), .B2(new_n512_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n668_), .B1(new_n510_), .B2(new_n513_), .ZN(new_n760_));
  AND4_X1   g559(.A1(new_n618_), .A2(new_n760_), .A3(new_n639_), .A4(new_n661_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(new_n516_), .A3(new_n497_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n759_), .A2(new_n762_), .ZN(G1332gat));
  NAND3_X1  g562(.A1(new_n761_), .A2(new_n518_), .A3(new_n732_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n757_), .A2(new_n732_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(KEYINPUT107), .B(KEYINPUT48), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n765_), .A2(G64gat), .A3(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n765_), .B2(G64gat), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n764_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT108), .ZN(G1333gat));
  INV_X1    g569(.A(G71gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n771_), .B1(new_n757_), .B2(new_n300_), .ZN(new_n772_));
  XOR2_X1   g571(.A(KEYINPUT109), .B(KEYINPUT49), .Z(new_n773_));
  XNOR2_X1  g572(.A(new_n772_), .B(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n761_), .A2(new_n771_), .A3(new_n300_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1334gat));
  AOI21_X1  g575(.A(new_n361_), .B1(new_n757_), .B2(new_n404_), .ZN(new_n777_));
  XOR2_X1   g576(.A(new_n777_), .B(KEYINPUT50), .Z(new_n778_));
  NAND3_X1  g577(.A1(new_n761_), .A2(new_n361_), .A3(new_n404_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(G1335gat));
  INV_X1    g579(.A(G85gat), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n697_), .A2(new_n619_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n760_), .A2(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n781_), .B1(new_n783_), .B2(new_n512_), .ZN(new_n784_));
  OR2_X1    g583(.A1(new_n784_), .A2(KEYINPUT110), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(KEYINPUT110), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n718_), .A2(new_n719_), .ZN(new_n787_));
  NOR3_X1   g586(.A1(new_n619_), .A2(new_n639_), .A3(new_n668_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n497_), .A2(G85gat), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT111), .ZN(new_n791_));
  AOI22_X1  g590(.A1(new_n785_), .A2(new_n786_), .B1(new_n789_), .B2(new_n791_), .ZN(G1336gat));
  INV_X1    g591(.A(G92gat), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n793_), .B1(new_n789_), .B2(new_n732_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n783_), .A2(G92gat), .A3(new_n507_), .ZN(new_n795_));
  OR2_X1    g594(.A1(new_n794_), .A2(new_n795_), .ZN(G1337gat));
  INV_X1    g595(.A(KEYINPUT112), .ZN(new_n797_));
  OR2_X1    g596(.A1(new_n797_), .A2(KEYINPUT51), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n548_), .B1(new_n789_), .B2(new_n300_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n783_), .A2(new_n301_), .A3(new_n578_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n798_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n797_), .A2(KEYINPUT51), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n801_), .B(new_n802_), .ZN(G1338gat));
  XNOR2_X1  g602(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n404_), .B(new_n788_), .C1(new_n703_), .C2(new_n711_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n805_), .A2(new_n806_), .A3(G106gat), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n805_), .B2(G106gat), .ZN(new_n808_));
  OR2_X1    g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n760_), .A2(new_n360_), .A3(new_n404_), .A4(new_n782_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n804_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n810_), .B(new_n804_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n811_), .A2(new_n813_), .ZN(G1339gat));
  NOR3_X1   g613(.A1(new_n301_), .A2(new_n512_), .A3(new_n675_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n816_));
  INV_X1    g615(.A(new_n613_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n817_), .A2(new_n669_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n603_), .A2(KEYINPUT12), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n819_), .A2(new_n589_), .B1(new_n598_), .B2(new_n595_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n820_), .A2(new_n821_), .A3(KEYINPUT55), .A4(new_n600_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n592_), .A2(new_n599_), .A3(KEYINPUT55), .A4(new_n600_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT115), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n592_), .A2(new_n599_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(G230gat), .A3(G233gat), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT55), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n601_), .A2(new_n827_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n822_), .A2(new_n824_), .A3(new_n826_), .A4(new_n828_), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n829_), .A2(KEYINPUT56), .A3(new_n610_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT56), .B1(new_n829_), .B2(new_n610_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n818_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n225_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n225_), .B1(new_n223_), .B2(new_n220_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n205_), .B1(new_n222_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n833_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n226_), .A2(new_n229_), .A3(new_n206_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n836_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n837_), .A2(new_n838_), .A3(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n612_), .B1(new_n601_), .B2(new_n605_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n840_), .B(KEYINPUT117), .C1(new_n841_), .C2(new_n817_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(KEYINPUT117), .B1(new_n614_), .B2(new_n840_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  AOI211_X1 g644(.A(new_n816_), .B(new_n666_), .C1(new_n832_), .C2(new_n845_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(KEYINPUT119), .A2(KEYINPUT58), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  NOR3_X1   g647(.A1(new_n830_), .A2(new_n831_), .A3(KEYINPUT118), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n829_), .A2(new_n610_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT56), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n850_), .A2(KEYINPUT118), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n840_), .A2(new_n613_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n848_), .B1(new_n849_), .B2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n850_), .A2(new_n851_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n829_), .A2(KEYINPUT56), .A3(new_n610_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n857_), .A2(new_n858_), .A3(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n853_), .B1(new_n831_), .B2(KEYINPUT118), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n860_), .A2(new_n847_), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n856_), .A2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n846_), .B1(new_n863_), .B2(new_n710_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n666_), .ZN(new_n865_));
  OR2_X1    g664(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n866_));
  INV_X1    g665(.A(new_n818_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n867_), .B1(new_n857_), .B2(new_n859_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n844_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n842_), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n865_), .B(new_n866_), .C1(new_n868_), .C2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n816_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n639_), .B1(new_n864_), .B2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n755_), .A2(KEYINPUT114), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT17), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT77), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n876_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n624_), .ZN(new_n878_));
  OAI22_X1  g677(.A1(new_n875_), .A2(new_n630_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n636_), .A2(new_n879_), .B1(new_n239_), .B2(new_n238_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT114), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n874_), .A2(new_n882_), .A3(new_n661_), .ZN(new_n883_));
  OAI21_X1  g682(.A(KEYINPUT54), .B1(new_n883_), .B2(new_n618_), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n880_), .A2(new_n881_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n885_), .A2(new_n886_), .A3(new_n619_), .A4(new_n874_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n884_), .A2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n511_), .B(new_n815_), .C1(new_n873_), .C2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT121), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n860_), .A2(new_n847_), .A3(new_n861_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n847_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n710_), .B1(new_n893_), .B2(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n666_), .B1(new_n832_), .B2(new_n845_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n896_), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n895_), .A2(new_n872_), .A3(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n638_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n888_), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n900_), .A2(KEYINPUT121), .A3(new_n511_), .A4(new_n815_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n892_), .A2(new_n668_), .A3(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(G113gat), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT59), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n890_), .A2(new_n904_), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n900_), .A2(KEYINPUT59), .A3(new_n511_), .A4(new_n815_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(KEYINPUT122), .B(G113gat), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n240_), .A2(new_n908_), .ZN(new_n909_));
  AOI22_X1  g708(.A1(new_n902_), .A2(new_n903_), .B1(new_n907_), .B2(new_n909_), .ZN(G1340gat));
  INV_X1    g709(.A(KEYINPUT60), .ZN(new_n911_));
  AOI21_X1  g710(.A(G120gat), .B1(new_n618_), .B2(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n912_), .B1(new_n911_), .B2(G120gat), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n892_), .A2(new_n901_), .A3(new_n913_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n619_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n915_));
  INV_X1    g714(.A(G120gat), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n914_), .B1(new_n915_), .B2(new_n916_), .ZN(G1341gat));
  NAND3_X1  g716(.A1(new_n892_), .A2(new_n639_), .A3(new_n901_), .ZN(new_n918_));
  INV_X1    g717(.A(G127gat), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n919_), .B1(new_n639_), .B2(KEYINPUT123), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n920_), .B1(KEYINPUT123), .B2(new_n919_), .ZN(new_n921_));
  AOI22_X1  g720(.A1(new_n918_), .A2(new_n919_), .B1(new_n907_), .B2(new_n921_), .ZN(G1342gat));
  INV_X1    g721(.A(G134gat), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n892_), .A2(new_n923_), .A3(new_n666_), .A4(new_n901_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n661_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n925_), .B2(new_n923_), .ZN(G1343gat));
  AOI21_X1  g725(.A(new_n889_), .B1(new_n898_), .B2(new_n638_), .ZN(new_n927_));
  NOR4_X1   g726(.A1(new_n300_), .A2(new_n511_), .A3(new_n732_), .A4(new_n512_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n927_), .A2(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(new_n668_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g731(.A1(new_n930_), .A2(new_n618_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g733(.A1(new_n930_), .A2(new_n639_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(KEYINPUT61), .B(G155gat), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n935_), .B(new_n936_), .ZN(G1346gat));
  INV_X1    g736(.A(KEYINPUT124), .ZN(new_n938_));
  INV_X1    g737(.A(G162gat), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n939_), .B1(new_n930_), .B2(new_n710_), .ZN(new_n940_));
  NOR4_X1   g739(.A1(new_n927_), .A2(G162gat), .A3(new_n865_), .A4(new_n929_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n938_), .B1(new_n940_), .B2(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n900_), .A2(new_n928_), .ZN(new_n943_));
  OAI21_X1  g742(.A(G162gat), .B1(new_n943_), .B2(new_n661_), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n930_), .A2(new_n939_), .A3(new_n666_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n944_), .A2(KEYINPUT124), .A3(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n942_), .A2(new_n946_), .ZN(G1347gat));
  NOR3_X1   g746(.A1(new_n301_), .A2(new_n497_), .A3(new_n731_), .ZN(new_n948_));
  NAND4_X1  g747(.A1(new_n900_), .A2(new_n511_), .A3(new_n668_), .A4(new_n948_), .ZN(new_n949_));
  OAI211_X1 g748(.A(KEYINPUT62), .B(G169gat), .C1(new_n949_), .C2(KEYINPUT22), .ZN(new_n950_));
  INV_X1    g749(.A(KEYINPUT62), .ZN(new_n951_));
  INV_X1    g750(.A(new_n948_), .ZN(new_n952_));
  NOR4_X1   g751(.A1(new_n927_), .A2(new_n404_), .A3(new_n669_), .A4(new_n952_), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n951_), .B1(new_n953_), .B2(new_n417_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n271_), .B1(new_n953_), .B2(new_n951_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n950_), .B1(new_n954_), .B2(new_n955_), .ZN(G1348gat));
  NAND3_X1  g755(.A1(new_n900_), .A2(new_n511_), .A3(new_n948_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n272_), .B1(new_n957_), .B2(new_n619_), .ZN(new_n958_));
  NAND3_X1  g757(.A1(new_n900_), .A2(KEYINPUT125), .A3(new_n511_), .ZN(new_n959_));
  INV_X1    g758(.A(KEYINPUT125), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n960_), .B1(new_n927_), .B2(new_n404_), .ZN(new_n961_));
  NOR3_X1   g760(.A1(new_n952_), .A2(new_n272_), .A3(new_n619_), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n959_), .A2(new_n961_), .A3(new_n962_), .ZN(new_n963_));
  AND2_X1   g762(.A1(new_n958_), .A2(new_n963_), .ZN(G1349gat));
  NOR3_X1   g763(.A1(new_n957_), .A2(new_n423_), .A3(new_n638_), .ZN(new_n965_));
  NAND4_X1  g764(.A1(new_n959_), .A2(new_n961_), .A3(new_n639_), .A4(new_n948_), .ZN(new_n966_));
  INV_X1    g765(.A(G183gat), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n965_), .B1(new_n966_), .B2(new_n967_), .ZN(G1350gat));
  NAND4_X1  g767(.A1(new_n900_), .A2(new_n511_), .A3(new_n710_), .A4(new_n948_), .ZN(new_n969_));
  INV_X1    g768(.A(KEYINPUT126), .ZN(new_n970_));
  AND3_X1   g769(.A1(new_n969_), .A2(new_n970_), .A3(G190gat), .ZN(new_n971_));
  AOI21_X1  g770(.A(new_n970_), .B1(new_n969_), .B2(G190gat), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n666_), .A2(new_n424_), .ZN(new_n973_));
  OAI22_X1  g772(.A1(new_n971_), .A2(new_n972_), .B1(new_n957_), .B2(new_n973_), .ZN(G1351gat));
  NAND3_X1  g773(.A1(new_n301_), .A2(new_n732_), .A3(new_n512_), .ZN(new_n975_));
  NOR3_X1   g774(.A1(new_n927_), .A2(new_n511_), .A3(new_n975_), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n976_), .A2(new_n668_), .ZN(new_n977_));
  XNOR2_X1  g776(.A(new_n977_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g777(.A1(new_n976_), .A2(new_n618_), .ZN(new_n979_));
  XNOR2_X1  g778(.A(new_n979_), .B(G204gat), .ZN(G1353gat));
  OR2_X1    g779(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n981_));
  AOI21_X1  g780(.A(new_n981_), .B1(new_n976_), .B2(new_n639_), .ZN(new_n982_));
  AND2_X1   g781(.A1(new_n976_), .A2(new_n639_), .ZN(new_n983_));
  XOR2_X1   g782(.A(KEYINPUT63), .B(G211gat), .Z(new_n984_));
  AOI21_X1  g783(.A(new_n982_), .B1(new_n983_), .B2(new_n984_), .ZN(G1354gat));
  AOI21_X1  g784(.A(G218gat), .B1(new_n976_), .B2(new_n666_), .ZN(new_n986_));
  NAND2_X1  g785(.A1(new_n710_), .A2(G218gat), .ZN(new_n987_));
  XNOR2_X1  g786(.A(new_n987_), .B(KEYINPUT127), .ZN(new_n988_));
  AOI21_X1  g787(.A(new_n986_), .B1(new_n976_), .B2(new_n988_), .ZN(G1355gat));
endmodule


