//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 1 0 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 0 0 0 1 0 0 0 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n601_, new_n602_, new_n603_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n679_, new_n680_,
    new_n681_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n811_, new_n813_, new_n814_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n844_, new_n846_,
    new_n847_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_;
  INV_X1    g000(.A(KEYINPUT76), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT25), .B(G183gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT26), .B(G190gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT24), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n205_), .B1(G169gat), .B2(G176gat), .ZN(new_n206_));
  INV_X1    g005(.A(G169gat), .ZN(new_n207_));
  INV_X1    g006(.A(G176gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  AOI22_X1  g008(.A1(new_n203_), .A2(new_n204_), .B1(new_n206_), .B2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(G183gat), .A3(G190gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  AND3_X1   g012(.A1(new_n213_), .A2(KEYINPUT73), .A3(KEYINPUT23), .ZN(new_n214_));
  AOI21_X1  g013(.A(KEYINPUT73), .B1(new_n213_), .B2(KEYINPUT23), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n212_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n205_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n210_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n207_), .A2(new_n208_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT22), .B(G169gat), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n219_), .B1(new_n220_), .B2(new_n208_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n213_), .A2(KEYINPUT23), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(new_n212_), .ZN(new_n223_));
  OR2_X1    g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n221_), .A2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n218_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT30), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT30), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n218_), .A2(new_n226_), .A3(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT74), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT74), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n228_), .A2(new_n233_), .A3(new_n230_), .ZN(new_n234_));
  XOR2_X1   g033(.A(G71gat), .B(G99gat), .Z(new_n235_));
  NAND2_X1  g034(.A1(G227gat), .A2(G233gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G15gat), .B(G43gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n232_), .A2(new_n234_), .A3(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT75), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n233_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n239_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n241_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT31), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n240_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n245_), .B1(new_n240_), .B2(new_n244_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G127gat), .B(G134gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G113gat), .B(G120gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NOR3_X1   g051(.A1(new_n247_), .A2(new_n248_), .A3(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n240_), .A2(new_n244_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT31), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n251_), .B1(new_n255_), .B2(new_n246_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n202_), .B1(new_n253_), .B2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n252_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n255_), .A2(new_n251_), .A3(new_n246_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n258_), .A2(new_n259_), .A3(KEYINPUT76), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(G155gat), .A2(G162gat), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT78), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n263_), .A2(KEYINPUT79), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT79), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n265_), .A2(KEYINPUT78), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n262_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(KEYINPUT78), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n263_), .A2(KEYINPUT79), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n269_), .B(new_n270_), .C1(G155gat), .C2(G162gat), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n267_), .A2(new_n268_), .A3(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT82), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G141gat), .A2(G148gat), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT2), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT3), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n276_), .B1(KEYINPUT81), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT77), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n279_), .B1(G141gat), .B2(G148gat), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n274_), .A2(KEYINPUT77), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n275_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT81), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n283_), .B1(KEYINPUT80), .B2(KEYINPUT3), .ZN(new_n284_));
  NOR2_X1   g083(.A1(G141gat), .A2(G148gat), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n285_), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n278_), .A2(new_n282_), .A3(new_n286_), .A4(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT82), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n267_), .A2(new_n271_), .A3(new_n289_), .A4(new_n268_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n273_), .A2(new_n288_), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT83), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT83), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n273_), .A2(new_n288_), .A3(new_n293_), .A4(new_n290_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n280_), .A2(new_n281_), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n267_), .A2(new_n271_), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n268_), .B(KEYINPUT1), .Z(new_n298_));
  AOI211_X1 g097(.A(new_n296_), .B(new_n285_), .C1(new_n297_), .C2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n295_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n252_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n299_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n251_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n302_), .A2(KEYINPUT4), .A3(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G225gat), .A2(G233gat), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n306_), .B(KEYINPUT92), .Z(new_n307_));
  INV_X1    g106(.A(KEYINPUT94), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n251_), .B1(new_n295_), .B2(new_n300_), .ZN(new_n309_));
  XOR2_X1   g108(.A(KEYINPUT93), .B(KEYINPUT4), .Z(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n308_), .B1(new_n309_), .B2(new_n311_), .ZN(new_n312_));
  NOR4_X1   g111(.A1(new_n303_), .A2(KEYINPUT94), .A3(new_n251_), .A4(new_n310_), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n305_), .B(new_n307_), .C1(new_n312_), .C2(new_n313_), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n302_), .A2(new_n304_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n306_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G1gat), .B(G29gat), .ZN(new_n318_));
  INV_X1    g117(.A(G85gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT0), .B(G57gat), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n320_), .B(new_n321_), .Z(new_n322_));
  NAND2_X1  g121(.A1(new_n317_), .A2(new_n322_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n324_));
  AND2_X1   g123(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n325_));
  AND2_X1   g124(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n326_));
  NOR2_X1   g125(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n327_));
  OAI22_X1  g126(.A1(new_n324_), .A2(new_n325_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n206_), .A2(new_n209_), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n328_), .A2(new_n329_), .A3(new_n217_), .ZN(new_n330_));
  AOI22_X1  g129(.A1(new_n330_), .A2(new_n216_), .B1(new_n225_), .B2(new_n221_), .ZN(new_n331_));
  AND2_X1   g130(.A1(G211gat), .A2(G218gat), .ZN(new_n332_));
  NOR2_X1   g131(.A1(G211gat), .A2(G218gat), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT21), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G197gat), .B(G204gat), .ZN(new_n337_));
  NOR3_X1   g136(.A1(new_n335_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(G204gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(G197gat), .ZN(new_n341_));
  INV_X1    g140(.A(G197gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(G204gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(new_n343_), .A3(new_n336_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT85), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT85), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n337_), .A2(new_n346_), .A3(new_n336_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n342_), .A2(G204gat), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n336_), .B1(new_n349_), .B2(KEYINPUT84), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT84), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n341_), .A2(new_n343_), .A3(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n334_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n348_), .A2(KEYINPUT86), .A3(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(KEYINPUT86), .B1(new_n348_), .B2(new_n353_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n331_), .B(new_n339_), .C1(new_n354_), .C2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n348_), .A2(new_n353_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT86), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n348_), .A2(new_n353_), .A3(KEYINPUT86), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n338_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n216_), .A2(new_n224_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n223_), .A2(new_n217_), .ZN(new_n363_));
  AOI22_X1  g162(.A1(new_n362_), .A2(new_n221_), .B1(new_n210_), .B2(new_n363_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n356_), .B(KEYINPUT20), .C1(new_n361_), .C2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G226gat), .A2(G233gat), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n366_), .B(new_n367_), .Z(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT90), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n365_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT20), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n339_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n371_), .B1(new_n372_), .B2(new_n227_), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n364_), .B(new_n339_), .C1(new_n354_), .C2(new_n355_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(new_n368_), .A3(new_n374_), .ZN(new_n375_));
  XOR2_X1   g174(.A(G64gat), .B(G92gat), .Z(new_n376_));
  XNOR2_X1  g175(.A(G8gat), .B(G36gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n370_), .A2(new_n375_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT27), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n374_), .B(KEYINPUT20), .C1(new_n361_), .C2(new_n331_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n368_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n364_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n371_), .B1(new_n372_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n369_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(new_n356_), .A3(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n381_), .B1(new_n386_), .B2(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n383_), .A2(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n384_), .A2(new_n385_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n389_), .B1(new_n388_), .B2(new_n356_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n380_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(KEYINPUT27), .B1(new_n395_), .B2(new_n382_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n392_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n322_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n314_), .A2(new_n316_), .A3(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n323_), .A2(new_n397_), .A3(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G22gat), .B(G50gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT28), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n301_), .A2(KEYINPUT29), .A3(new_n403_), .ZN(new_n404_));
  XOR2_X1   g203(.A(G78gat), .B(G106gat), .Z(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n406_), .A2(KEYINPUT88), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT29), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n402_), .B1(new_n303_), .B2(new_n408_), .ZN(new_n409_));
  OR3_X1    g208(.A1(new_n404_), .A2(new_n407_), .A3(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n372_), .B1(new_n303_), .B2(new_n408_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G228gat), .A2(G233gat), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n412_), .B1(new_n372_), .B2(KEYINPUT87), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n411_), .B(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n406_), .B1(new_n404_), .B2(new_n409_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n410_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n414_), .B1(new_n410_), .B2(new_n415_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n261_), .B1(new_n400_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT33), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n399_), .A2(new_n421_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n314_), .A2(KEYINPUT33), .A3(new_n316_), .A4(new_n398_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n395_), .A2(new_n382_), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n305_), .B(new_n306_), .C1(new_n312_), .C2(new_n313_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n398_), .B1(new_n315_), .B2(new_n307_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n424_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n422_), .A2(new_n423_), .A3(new_n427_), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n386_), .A2(new_n390_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n370_), .A2(new_n375_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n381_), .A2(KEYINPUT32), .ZN(new_n431_));
  MUX2_X1   g230(.A(new_n429_), .B(new_n430_), .S(new_n431_), .Z(new_n432_));
  AND3_X1   g231(.A1(new_n314_), .A2(new_n316_), .A3(new_n398_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n398_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n432_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n410_), .A2(new_n415_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n414_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n416_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n428_), .A2(new_n435_), .A3(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n420_), .A2(new_n440_), .A3(KEYINPUT95), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n258_), .A2(new_n259_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n439_), .A2(new_n397_), .A3(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n433_), .A2(new_n434_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n441_), .A2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT95), .B1(new_n420_), .B2(new_n440_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G43gat), .B(G50gat), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT66), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n450_), .A2(new_n451_), .ZN(new_n453_));
  XOR2_X1   g252(.A(G29gat), .B(G36gat), .Z(new_n454_));
  OR3_X1    g253(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n454_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT71), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G15gat), .B(G22gat), .ZN(new_n460_));
  INV_X1    g259(.A(G1gat), .ZN(new_n461_));
  INV_X1    g260(.A(G8gat), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT14), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n460_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G1gat), .B(G8gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n459_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n457_), .B(KEYINPUT15), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(new_n466_), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G229gat), .A2(G233gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n459_), .B(new_n467_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n472_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n473_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G113gat), .B(G141gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G169gat), .B(G197gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(KEYINPUT72), .ZN(new_n481_));
  XOR2_X1   g280(.A(new_n477_), .B(new_n481_), .Z(new_n482_));
  NAND2_X1  g281(.A1(G99gat), .A2(G106gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT6), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n485_));
  OR3_X1    g284(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n484_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  XOR2_X1   g286(.A(G85gat), .B(G92gat), .Z(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT8), .ZN(new_n490_));
  XOR2_X1   g289(.A(KEYINPUT10), .B(G99gat), .Z(new_n491_));
  INV_X1    g290(.A(G106gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n488_), .A2(KEYINPUT9), .ZN(new_n494_));
  INV_X1    g293(.A(G92gat), .ZN(new_n495_));
  OR3_X1    g294(.A1(new_n319_), .A2(new_n495_), .A3(KEYINPUT9), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n493_), .A2(new_n494_), .A3(new_n496_), .A4(new_n484_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n490_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G71gat), .B(G78gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G57gat), .B(G64gat), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n499_), .B1(KEYINPUT11), .B2(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n501_), .B1(KEYINPUT11), .B2(new_n500_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n500_), .A2(new_n499_), .A3(KEYINPUT11), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n498_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n490_), .A2(new_n497_), .A3(new_n504_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(KEYINPUT12), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT12), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n498_), .A2(new_n509_), .A3(new_n505_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G230gat), .A2(G233gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n506_), .A2(new_n507_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n513_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G176gat), .B(G204gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G120gat), .B(G148gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT64), .B(KEYINPUT5), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n515_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT65), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n515_), .A2(new_n520_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n521_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n515_), .A2(KEYINPUT65), .A3(new_n520_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT13), .ZN(new_n527_));
  NOR3_X1   g326(.A1(new_n449_), .A2(new_n482_), .A3(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G231gat), .A2(G233gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n466_), .B(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(new_n504_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G127gat), .B(G155gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(G211gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT16), .B(G183gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(new_n534_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n535_), .A2(KEYINPUT17), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n535_), .A2(KEYINPUT17), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n531_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n538_), .B1(new_n536_), .B2(new_n531_), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n539_), .B(KEYINPUT69), .Z(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT70), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT37), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G134gat), .B(G162gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT68), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G190gat), .B(G218gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT36), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n546_), .A2(new_n547_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G232gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT34), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n552_), .A2(KEYINPUT35), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n469_), .A2(new_n498_), .ZN(new_n554_));
  AND2_X1   g353(.A1(new_n554_), .A2(KEYINPUT67), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n490_), .A2(new_n497_), .A3(new_n457_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n556_), .B1(new_n554_), .B2(KEYINPUT67), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n553_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n552_), .A2(KEYINPUT35), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n553_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n554_), .A2(new_n556_), .A3(new_n560_), .ZN(new_n561_));
  AOI211_X1 g360(.A(new_n549_), .B(new_n550_), .C1(new_n558_), .C2(new_n561_), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n558_), .A2(new_n547_), .A3(new_n546_), .A4(new_n561_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n542_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n550_), .B1(new_n558_), .B2(new_n561_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(new_n548_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n567_), .A2(KEYINPUT37), .A3(new_n563_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n565_), .A2(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n541_), .A2(new_n569_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n528_), .A2(new_n461_), .A3(new_n570_), .A4(new_n445_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n572_), .A2(KEYINPUT38), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n573_), .B(KEYINPUT96), .Z(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(KEYINPUT38), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n567_), .A2(new_n563_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n577_), .A2(new_n540_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n528_), .A2(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(G1gat), .B1(new_n579_), .B2(new_n444_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n574_), .A2(new_n575_), .A3(new_n580_), .ZN(G1324gat));
  NAND2_X1  g380(.A1(new_n528_), .A2(new_n570_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n582_), .A2(G8gat), .A3(new_n397_), .ZN(new_n583_));
  OR3_X1    g382(.A1(new_n579_), .A2(KEYINPUT97), .A3(new_n397_), .ZN(new_n584_));
  OAI21_X1  g383(.A(KEYINPUT97), .B1(new_n579_), .B2(new_n397_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(G8gat), .A3(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT39), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT39), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n584_), .A2(new_n588_), .A3(G8gat), .A4(new_n585_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n583_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(KEYINPUT98), .B(KEYINPUT40), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n590_), .B(new_n592_), .ZN(G1325gat));
  INV_X1    g392(.A(new_n261_), .ZN(new_n594_));
  OAI21_X1  g393(.A(G15gat), .B1(new_n579_), .B2(new_n594_), .ZN(new_n595_));
  XOR2_X1   g394(.A(KEYINPUT99), .B(KEYINPUT41), .Z(new_n596_));
  OR2_X1    g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n596_), .ZN(new_n598_));
  OR3_X1    g397(.A1(new_n582_), .A2(G15gat), .A3(new_n594_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n597_), .A2(new_n598_), .A3(new_n599_), .ZN(G1326gat));
  OAI21_X1  g399(.A(G22gat), .B1(new_n579_), .B2(new_n439_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT42), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n439_), .A2(G22gat), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n602_), .B1(new_n582_), .B2(new_n603_), .ZN(G1327gat));
  INV_X1    g403(.A(new_n527_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n482_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n605_), .A2(new_n541_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n565_), .A2(KEYINPUT100), .A3(new_n568_), .ZN(new_n609_));
  AOI21_X1  g408(.A(KEYINPUT100), .B1(new_n565_), .B2(new_n568_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n611_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n612_), .A2(KEYINPUT101), .A3(KEYINPUT43), .ZN(new_n613_));
  INV_X1    g412(.A(new_n569_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n614_), .A2(KEYINPUT43), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n615_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n613_), .A2(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT101), .B1(new_n612_), .B2(KEYINPUT43), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n608_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT44), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  OAI211_X1 g420(.A(KEYINPUT44), .B(new_n608_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n621_), .A2(new_n445_), .A3(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(G29gat), .ZN(new_n624_));
  INV_X1    g423(.A(new_n541_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n625_), .A2(new_n576_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n528_), .A2(new_n626_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n444_), .A2(G29gat), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n624_), .B1(new_n627_), .B2(new_n628_), .ZN(G1328gat));
  NOR3_X1   g428(.A1(new_n627_), .A2(G36gat), .A3(new_n397_), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n630_), .B(KEYINPUT45), .Z(new_n631_));
  INV_X1    g430(.A(new_n397_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n621_), .A2(new_n632_), .A3(new_n622_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT102), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n633_), .A2(new_n634_), .A3(G36gat), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n634_), .B1(new_n633_), .B2(G36gat), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n631_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  OAI221_X1 g438(.A(new_n631_), .B1(KEYINPUT103), .B2(KEYINPUT46), .C1(new_n635_), .C2(new_n636_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1329gat));
  NOR3_X1   g440(.A1(new_n627_), .A2(G43gat), .A3(new_n594_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n621_), .A2(new_n442_), .A3(new_n622_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n642_), .B1(new_n643_), .B2(G43gat), .ZN(new_n644_));
  XNOR2_X1  g443(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(G1330gat));
  NAND3_X1  g445(.A1(new_n621_), .A2(new_n419_), .A3(new_n622_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(G50gat), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n439_), .A2(G50gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n648_), .B1(new_n627_), .B2(new_n649_), .ZN(G1331gat));
  NAND2_X1  g449(.A1(new_n527_), .A2(new_n570_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT105), .Z(new_n652_));
  NOR2_X1   g451(.A1(new_n449_), .A2(new_n606_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(G57gat), .B1(new_n655_), .B2(new_n445_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n653_), .A2(new_n527_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n658_), .A2(new_n576_), .A3(new_n625_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(G57gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n661_), .B1(new_n445_), .B2(KEYINPUT106), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n662_), .B1(KEYINPUT106), .B2(new_n661_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n656_), .B1(new_n660_), .B2(new_n663_), .ZN(G1332gat));
  OAI21_X1  g463(.A(G64gat), .B1(new_n659_), .B2(new_n397_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT48), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n397_), .A2(G64gat), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n666_), .B1(new_n654_), .B2(new_n667_), .ZN(G1333gat));
  NOR2_X1   g467(.A1(new_n594_), .A2(G71gat), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT107), .Z(new_n670_));
  NAND2_X1  g469(.A1(new_n655_), .A2(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(G71gat), .B1(new_n659_), .B2(new_n594_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n672_), .A2(KEYINPUT49), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT49), .ZN(new_n674_));
  OAI211_X1 g473(.A(new_n674_), .B(G71gat), .C1(new_n659_), .C2(new_n594_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n671_), .B1(new_n673_), .B2(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT108), .ZN(G1334gat));
  OAI21_X1  g477(.A(G78gat), .B1(new_n659_), .B2(new_n439_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT50), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n439_), .A2(G78gat), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n680_), .B1(new_n654_), .B2(new_n681_), .ZN(G1335gat));
  NAND2_X1  g481(.A1(new_n658_), .A2(new_n626_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n319_), .B1(new_n683_), .B2(new_n444_), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT109), .Z(new_n685_));
  OR2_X1    g484(.A1(new_n617_), .A2(new_n618_), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n605_), .A2(new_n625_), .A3(new_n606_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT110), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n686_), .A2(KEYINPUT110), .A3(new_n687_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n690_), .A2(G85gat), .A3(new_n445_), .A4(new_n691_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n685_), .A2(new_n692_), .ZN(G1336gat));
  NAND4_X1  g492(.A1(new_n690_), .A2(G92gat), .A3(new_n632_), .A4(new_n691_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n495_), .B1(new_n683_), .B2(new_n397_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1337gat));
  NAND3_X1  g495(.A1(new_n690_), .A2(new_n261_), .A3(new_n691_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(G99gat), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n658_), .A2(new_n491_), .A3(new_n442_), .A4(new_n626_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT51), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT51), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n698_), .A2(new_n702_), .A3(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(G1338gat));
  NAND4_X1  g503(.A1(new_n658_), .A2(new_n492_), .A3(new_n419_), .A4(new_n626_), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n419_), .B(new_n687_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT111), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT52), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n492_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n708_), .A2(new_n709_), .A3(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n709_), .B1(new_n708_), .B2(new_n710_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n705_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT53), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT53), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n715_), .B(new_n705_), .C1(new_n711_), .C2(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1339gat));
  INV_X1    g516(.A(KEYINPUT113), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n512_), .B1(new_n511_), .B2(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n719_), .B1(new_n718_), .B2(new_n511_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT55), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n513_), .A2(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(KEYINPUT114), .B1(new_n513_), .B2(new_n721_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT114), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n511_), .A2(new_n724_), .A3(KEYINPUT55), .A4(new_n512_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n720_), .A2(new_n722_), .A3(new_n723_), .A4(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT56), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n726_), .A2(new_n727_), .A3(new_n520_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n728_), .A2(new_n521_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n726_), .A2(new_n520_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT56), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n729_), .A2(new_n606_), .A3(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n480_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n471_), .A2(new_n475_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n474_), .A2(new_n472_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n733_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n480_), .B1(new_n473_), .B2(new_n476_), .ZN(new_n737_));
  OR3_X1    g536(.A1(new_n736_), .A2(new_n737_), .A3(KEYINPUT115), .ZN(new_n738_));
  OAI21_X1  g537(.A(KEYINPUT115), .B1(new_n736_), .B2(new_n737_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n526_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n577_), .B1(new_n732_), .B2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT58), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT118), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n738_), .A2(new_n739_), .A3(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n729_), .A2(new_n746_), .A3(new_n731_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT117), .ZN(new_n748_));
  AOI21_X1  g547(.A(KEYINPUT118), .B1(new_n748_), .B2(new_n744_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n614_), .B1(new_n747_), .B2(new_n750_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n729_), .A2(new_n746_), .A3(new_n731_), .A4(new_n749_), .ZN(new_n752_));
  AOI22_X1  g551(.A1(KEYINPUT57), .A2(new_n743_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n743_), .A2(KEYINPUT116), .A3(KEYINPUT57), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT116), .ZN(new_n755_));
  AND4_X1   g554(.A1(new_n606_), .A2(new_n731_), .A3(new_n521_), .A4(new_n728_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n576_), .B1(new_n756_), .B2(new_n741_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT57), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n755_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n753_), .B1(new_n754_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT119), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT119), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n753_), .B(new_n762_), .C1(new_n754_), .C2(new_n759_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n761_), .A2(new_n540_), .A3(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n570_), .A2(new_n482_), .ZN(new_n765_));
  OR4_X1    g564(.A1(KEYINPUT112), .A2(new_n765_), .A3(KEYINPUT54), .A4(new_n527_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n605_), .A2(new_n570_), .A3(new_n482_), .ZN(new_n767_));
  OAI21_X1  g566(.A(KEYINPUT112), .B1(new_n767_), .B2(KEYINPUT54), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(KEYINPUT54), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n766_), .A2(new_n768_), .A3(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n764_), .A2(new_n770_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n443_), .A2(new_n444_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT59), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n753_), .B1(KEYINPUT57), .B2(new_n743_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n541_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n770_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT59), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n777_), .A2(new_n778_), .A3(new_n772_), .ZN(new_n779_));
  INV_X1    g578(.A(G113gat), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n482_), .A2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n774_), .A2(new_n779_), .A3(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n780_), .B1(new_n773_), .B2(new_n482_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n782_), .A2(new_n783_), .ZN(G1340gat));
  INV_X1    g583(.A(new_n772_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n785_), .B1(new_n764_), .B2(new_n770_), .ZN(new_n786_));
  INV_X1    g585(.A(G120gat), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n787_), .B1(new_n605_), .B2(KEYINPUT60), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n786_), .B(new_n788_), .C1(KEYINPUT60), .C2(new_n787_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n527_), .B(new_n779_), .C1(new_n786_), .C2(new_n778_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n789_), .B1(new_n791_), .B2(new_n787_), .ZN(G1341gat));
  XNOR2_X1  g591(.A(KEYINPUT120), .B(G127gat), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n540_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n774_), .A2(new_n779_), .A3(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(G127gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n796_), .B1(new_n773_), .B2(new_n541_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n795_), .A2(new_n797_), .ZN(G1342gat));
  INV_X1    g597(.A(G134gat), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n614_), .A2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n774_), .A2(new_n779_), .A3(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n799_), .B1(new_n773_), .B2(new_n576_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n801_), .A2(new_n802_), .ZN(G1343gat));
  NOR2_X1   g602(.A1(new_n261_), .A2(new_n439_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n805_), .B1(new_n764_), .B2(new_n770_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n444_), .A2(new_n632_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n806_), .A2(new_n606_), .A3(new_n807_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(KEYINPUT121), .B(G141gat), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n808_), .B(new_n809_), .ZN(G1344gat));
  NAND3_X1  g609(.A1(new_n806_), .A2(new_n527_), .A3(new_n807_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g611(.A1(new_n806_), .A2(new_n625_), .A3(new_n807_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(KEYINPUT61), .B(G155gat), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n813_), .B(new_n814_), .ZN(G1346gat));
  AND2_X1   g614(.A1(new_n806_), .A2(new_n807_), .ZN(new_n816_));
  INV_X1    g615(.A(G162gat), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n609_), .A2(new_n610_), .A3(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n806_), .A2(new_n577_), .A3(new_n807_), .ZN(new_n819_));
  AOI22_X1  g618(.A1(new_n816_), .A2(new_n818_), .B1(new_n819_), .B2(new_n817_), .ZN(G1347gat));
  NOR2_X1   g619(.A1(new_n445_), .A2(new_n397_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n261_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(KEYINPUT122), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n439_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n824_), .B1(new_n776_), .B2(new_n770_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(new_n606_), .A3(new_n220_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n207_), .B1(new_n825_), .B2(new_n606_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT62), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n827_), .A2(KEYINPUT123), .A3(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n828_), .B2(new_n827_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT123), .B1(new_n827_), .B2(new_n828_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n826_), .B1(new_n830_), .B2(new_n831_), .ZN(G1348gat));
  INV_X1    g631(.A(new_n825_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n208_), .B1(new_n833_), .B2(new_n605_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n771_), .A2(new_n439_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n823_), .A2(G176gat), .A3(new_n527_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n834_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT124), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n834_), .B(KEYINPUT124), .C1(new_n835_), .C2(new_n836_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(G1349gat));
  NOR3_X1   g640(.A1(new_n833_), .A2(new_n540_), .A3(new_n203_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n771_), .A2(new_n625_), .A3(new_n439_), .A4(new_n823_), .ZN(new_n843_));
  INV_X1    g642(.A(G183gat), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n842_), .B1(new_n843_), .B2(new_n844_), .ZN(G1350gat));
  OAI21_X1  g644(.A(G190gat), .B1(new_n833_), .B2(new_n614_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n825_), .A2(new_n577_), .A3(new_n204_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(G1351gat));
  NAND3_X1  g647(.A1(new_n806_), .A2(new_n606_), .A3(new_n821_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g649(.A(new_n821_), .ZN(new_n851_));
  AOI211_X1 g650(.A(new_n805_), .B(new_n851_), .C1(new_n764_), .C2(new_n770_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n527_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n853_), .A2(KEYINPUT125), .A3(G204gat), .ZN(new_n854_));
  NAND2_X1  g653(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n852_), .A2(new_n527_), .A3(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n856_), .ZN(G1353gat));
  INV_X1    g656(.A(new_n540_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n771_), .A2(new_n858_), .A3(new_n804_), .A4(new_n821_), .ZN(new_n859_));
  XOR2_X1   g658(.A(KEYINPUT63), .B(G211gat), .Z(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(KEYINPUT126), .B1(new_n859_), .B2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT126), .ZN(new_n863_));
  NAND4_X1  g662(.A1(new_n852_), .A2(new_n863_), .A3(new_n858_), .A4(new_n860_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n859_), .A2(new_n865_), .ZN(new_n866_));
  AND3_X1   g665(.A1(new_n862_), .A2(new_n864_), .A3(new_n866_), .ZN(G1354gat));
  NAND2_X1  g666(.A1(new_n852_), .A2(new_n577_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(KEYINPUT127), .B(G218gat), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n614_), .A2(new_n869_), .ZN(new_n870_));
  AOI22_X1  g669(.A1(new_n868_), .A2(new_n869_), .B1(new_n852_), .B2(new_n870_), .ZN(G1355gat));
endmodule


