//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 0 1 1 0 1 0 1 0 1 1 1 0 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 1 1 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n619_, new_n620_, new_n621_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n810_, new_n811_, new_n812_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n819_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n856_, new_n857_,
    new_n859_, new_n860_, new_n861_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_,
    new_n881_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(G1gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n202_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT72), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G231gat), .A2(G233gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n209_), .B(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G57gat), .B(G64gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT11), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(KEYINPUT11), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT67), .B(G71gat), .ZN(new_n216_));
  INV_X1    g015(.A(G78gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n216_), .B(new_n217_), .ZN(new_n218_));
  MUX2_X1   g017(.A(new_n214_), .B(new_n215_), .S(new_n218_), .Z(new_n219_));
  XNOR2_X1  g018(.A(new_n212_), .B(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT73), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G127gat), .B(G155gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(KEYINPUT16), .ZN(new_n224_));
  XOR2_X1   g023(.A(G183gat), .B(G211gat), .Z(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT17), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n222_), .B(new_n228_), .ZN(new_n229_));
  OR3_X1    g028(.A1(new_n220_), .A2(KEYINPUT17), .A3(new_n227_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT37), .ZN(new_n232_));
  XOR2_X1   g031(.A(G85gat), .B(G92gat), .Z(new_n233_));
  NOR2_X1   g032(.A1(G99gat), .A2(G106gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT7), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G99gat), .A2(G106gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT6), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n233_), .B1(new_n236_), .B2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT8), .ZN(new_n241_));
  INV_X1    g040(.A(G85gat), .ZN(new_n242_));
  INV_X1    g041(.A(G92gat), .ZN(new_n243_));
  NOR3_X1   g042(.A1(new_n242_), .A2(new_n243_), .A3(KEYINPUT9), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n239_), .A2(new_n244_), .ZN(new_n245_));
  XOR2_X1   g044(.A(KEYINPUT10), .B(G99gat), .Z(new_n246_));
  XOR2_X1   g045(.A(KEYINPUT66), .B(G106gat), .Z(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n233_), .A2(KEYINPUT9), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n245_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n241_), .A2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G29gat), .B(G36gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G43gat), .B(G50gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G232gat), .A2(G233gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT34), .ZN(new_n257_));
  OAI22_X1  g056(.A1(new_n251_), .A2(new_n255_), .B1(KEYINPUT35), .B2(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n254_), .B(KEYINPUT15), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n251_), .A2(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n257_), .A2(KEYINPUT35), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  OAI211_X1 g062(.A(KEYINPUT35), .B(new_n257_), .C1(new_n258_), .C2(new_n260_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G190gat), .B(G218gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G134gat), .B(G162gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n267_), .A2(KEYINPUT36), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n263_), .A2(new_n264_), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n263_), .A2(new_n264_), .ZN(new_n270_));
  XOR2_X1   g069(.A(new_n267_), .B(KEYINPUT36), .Z(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n269_), .B1(new_n272_), .B2(KEYINPUT71), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n274_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n232_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n272_), .A2(KEYINPUT37), .A3(new_n269_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n231_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n251_), .A2(new_n219_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n251_), .A2(new_n219_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n281_), .B1(new_n282_), .B2(KEYINPUT12), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G230gat), .A2(G233gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n251_), .A2(new_n219_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT68), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT12), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n287_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n288_), .B1(new_n287_), .B2(new_n289_), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n283_), .B(new_n286_), .C1(new_n291_), .C2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT69), .ZN(new_n294_));
  OAI21_X1  g093(.A(KEYINPUT68), .B1(new_n282_), .B2(KEYINPUT12), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(new_n290_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT69), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n296_), .A2(new_n297_), .A3(new_n286_), .A4(new_n283_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n286_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n299_), .B1(new_n282_), .B2(new_n281_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n294_), .A2(new_n298_), .A3(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G120gat), .B(G148gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT5), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G176gat), .B(G204gat), .ZN(new_n304_));
  XOR2_X1   g103(.A(new_n303_), .B(new_n304_), .Z(new_n305_));
  NAND2_X1  g104(.A1(new_n301_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n305_), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n294_), .A2(new_n298_), .A3(new_n300_), .A4(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT70), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n309_), .B1(new_n310_), .B2(KEYINPUT13), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n312_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT85), .B(G43gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT31), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G227gat), .A2(G233gat), .ZN(new_n318_));
  INV_X1    g117(.A(G15gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(G71gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(G99gat), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT24), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n324_), .B1(G169gat), .B2(G176gat), .ZN(new_n325_));
  NOR2_X1   g124(.A1(G169gat), .A2(G176gat), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT81), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n325_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT80), .ZN(new_n331_));
  INV_X1    g130(.A(G190gat), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT26), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT25), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT78), .B1(new_n334_), .B2(G183gat), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT78), .ZN(new_n336_));
  INV_X1    g135(.A(G183gat), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n336_), .A2(new_n337_), .A3(KEYINPUT25), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT26), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n339_), .A2(KEYINPUT80), .A3(G190gat), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n333_), .A2(new_n335_), .A3(new_n338_), .A4(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT79), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n342_), .B1(new_n334_), .B2(G183gat), .ZN(new_n343_));
  NOR3_X1   g142(.A1(new_n337_), .A2(KEYINPUT79), .A3(KEYINPUT25), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n330_), .B1(new_n341_), .B2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT82), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT82), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n348_), .B(new_n330_), .C1(new_n341_), .C2(new_n345_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n328_), .A2(new_n329_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n324_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G183gat), .A2(G190gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT23), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT23), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n354_), .A2(G183gat), .A3(G190gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n347_), .A2(new_n349_), .A3(new_n351_), .A4(new_n356_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(G183gat), .A2(G190gat), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n358_), .B1(new_n354_), .B2(new_n352_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n360_));
  AOI22_X1  g159(.A1(new_n359_), .A2(new_n360_), .B1(G169gat), .B2(G176gat), .ZN(new_n361_));
  XOR2_X1   g160(.A(KEYINPUT84), .B(G176gat), .Z(new_n362_));
  INV_X1    g161(.A(G169gat), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT83), .B1(new_n363_), .B2(KEYINPUT22), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT22), .B(G169gat), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n366_), .A2(KEYINPUT83), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n361_), .B1(new_n365_), .B2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n357_), .A2(KEYINPUT30), .A3(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(KEYINPUT30), .B1(new_n357_), .B2(new_n368_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n323_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n357_), .A2(new_n368_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT30), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n375_), .A2(new_n369_), .A3(new_n322_), .ZN(new_n376_));
  XOR2_X1   g175(.A(G127gat), .B(G134gat), .Z(new_n377_));
  XOR2_X1   g176(.A(G113gat), .B(G120gat), .Z(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n372_), .A2(new_n376_), .A3(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n379_), .B1(new_n372_), .B2(new_n376_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n317_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n372_), .A2(new_n376_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n379_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n372_), .A2(new_n376_), .A3(new_n379_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(new_n316_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n382_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G1gat), .B(G29gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(G85gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT0), .B(G57gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n390_), .B(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G141gat), .A2(G148gat), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT86), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(G141gat), .ZN(new_n397_));
  INV_X1    g196(.A(G148gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(KEYINPUT86), .A2(G141gat), .A3(G148gat), .ZN(new_n400_));
  NAND3_X1  g199(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n396_), .A2(new_n399_), .A3(new_n400_), .A4(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G155gat), .A2(G162gat), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT1), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(G155gat), .A2(G162gat), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT87), .B1(new_n402_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n400_), .ZN(new_n409_));
  AOI21_X1  g208(.A(KEYINPUT86), .B1(G141gat), .B2(G148gat), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  AND2_X1   g210(.A1(G155gat), .A2(G162gat), .ZN(new_n412_));
  AOI22_X1  g211(.A1(new_n412_), .A2(KEYINPUT1), .B1(new_n397_), .B2(new_n398_), .ZN(new_n413_));
  OR2_X1    g212(.A1(G155gat), .A2(G162gat), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n414_), .A2(new_n404_), .A3(new_n403_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT87), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n411_), .A2(new_n413_), .A3(new_n415_), .A4(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n408_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT2), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n396_), .A2(new_n419_), .A3(new_n400_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n421_));
  NAND3_X1  g220(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  OR3_X1    g222(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n420_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n412_), .A2(new_n406_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n418_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n428_), .A2(KEYINPUT100), .A3(new_n384_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT100), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n408_), .A2(new_n417_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n430_), .B1(new_n431_), .B2(new_n379_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n429_), .A2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT101), .B1(new_n428_), .B2(new_n384_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT101), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n431_), .A2(new_n435_), .A3(new_n379_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n433_), .A2(KEYINPUT4), .A3(new_n434_), .A4(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G225gat), .A2(G233gat), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n431_), .A2(new_n379_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT4), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n438_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n437_), .A2(new_n441_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n433_), .A2(new_n438_), .A3(new_n434_), .A4(new_n436_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n393_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n442_), .A2(new_n443_), .A3(new_n393_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n388_), .A2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(G228gat), .B1(KEYINPUT89), .B2(G233gat), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n449_), .B1(KEYINPUT89), .B2(G233gat), .ZN(new_n450_));
  INV_X1    g249(.A(G197gat), .ZN(new_n451_));
  INV_X1    g250(.A(G204gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G197gat), .A2(G204gat), .ZN(new_n454_));
  AOI21_X1  g253(.A(KEYINPUT21), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  OR2_X1    g254(.A1(new_n455_), .A2(KEYINPUT90), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT91), .ZN(new_n457_));
  INV_X1    g256(.A(G218gat), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n458_), .A2(G211gat), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n458_), .A2(G211gat), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n457_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G211gat), .B(G218gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT91), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n453_), .A2(new_n454_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT21), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n455_), .A2(KEYINPUT90), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n456_), .A2(new_n464_), .A3(new_n468_), .A4(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n467_), .A2(new_n463_), .A3(new_n461_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT88), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n450_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT29), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n472_), .B1(new_n475_), .B2(new_n431_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  OAI221_X1 g276(.A(new_n472_), .B1(new_n473_), .B2(new_n450_), .C1(new_n475_), .C2(new_n431_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G78gat), .B(G106gat), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G22gat), .B(G50gat), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n431_), .A2(new_n475_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT28), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n483_), .A2(KEYINPUT28), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n482_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n486_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(new_n484_), .A3(new_n481_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n480_), .A2(new_n487_), .A3(new_n489_), .ZN(new_n490_));
  AOI211_X1 g289(.A(KEYINPUT93), .B(new_n479_), .C1(new_n477_), .C2(new_n478_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n479_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT93), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n487_), .A2(new_n489_), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n477_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n496_), .B1(new_n497_), .B2(new_n493_), .ZN(new_n498_));
  AOI22_X1  g297(.A1(new_n492_), .A2(new_n495_), .B1(new_n498_), .B2(KEYINPUT92), .ZN(new_n499_));
  OR2_X1    g298(.A1(new_n498_), .A2(KEYINPUT92), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G226gat), .A2(G233gat), .ZN(new_n503_));
  XOR2_X1   g302(.A(new_n502_), .B(new_n503_), .Z(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  AOI22_X1  g304(.A1(new_n357_), .A2(new_n368_), .B1(new_n471_), .B2(new_n470_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT95), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n366_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n366_), .A2(new_n507_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(new_n509_), .A3(new_n362_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(new_n361_), .ZN(new_n511_));
  AOI22_X1  g310(.A1(new_n353_), .A2(new_n355_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n512_));
  XOR2_X1   g311(.A(KEYINPUT25), .B(G183gat), .Z(new_n513_));
  XOR2_X1   g312(.A(KEYINPUT26), .B(G190gat), .Z(new_n514_));
  OAI211_X1 g313(.A(new_n330_), .B(new_n512_), .C1(new_n513_), .C2(new_n514_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n511_), .A2(new_n470_), .A3(new_n471_), .A4(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT20), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n505_), .B1(new_n506_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT20), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n511_), .A2(new_n515_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n519_), .B1(new_n520_), .B2(new_n472_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n521_), .B(new_n504_), .C1(new_n373_), .C2(new_n472_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n518_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT104), .ZN(new_n524_));
  XOR2_X1   g323(.A(G64gat), .B(G92gat), .Z(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT98), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT99), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n526_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G8gat), .B(G36gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n523_), .A2(new_n524_), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n506_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n516_), .A2(KEYINPUT20), .A3(new_n504_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT96), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n534_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n521_), .B1(new_n373_), .B2(new_n472_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(new_n505_), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT96), .B1(new_n506_), .B2(new_n535_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n538_), .A2(new_n540_), .A3(new_n531_), .A4(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n533_), .A2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n524_), .B1(new_n523_), .B2(new_n532_), .ZN(new_n544_));
  OAI21_X1  g343(.A(KEYINPUT27), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n538_), .A2(new_n540_), .A3(new_n541_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n532_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT27), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n547_), .A2(new_n548_), .A3(new_n542_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n545_), .A2(new_n549_), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n448_), .A2(new_n501_), .A3(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n523_), .A2(KEYINPUT32), .A3(new_n531_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n531_), .A2(KEYINPUT32), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n553_), .A2(new_n541_), .A3(new_n538_), .A4(new_n540_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n446_), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n552_), .B(new_n554_), .C1(new_n555_), .C2(new_n444_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT102), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT33), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n392_), .A2(new_n558_), .ZN(new_n559_));
  AND4_X1   g358(.A1(new_n557_), .A2(new_n442_), .A3(new_n443_), .A4(new_n559_), .ZN(new_n560_));
  AND2_X1   g359(.A1(new_n443_), .A2(new_n559_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n557_), .B1(new_n561_), .B2(new_n442_), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n542_), .B(new_n547_), .C1(new_n560_), .C2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n446_), .A2(new_n558_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n438_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n565_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n437_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT103), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n433_), .A2(new_n565_), .A3(new_n434_), .A4(new_n436_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(new_n392_), .A3(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n567_), .A2(KEYINPUT103), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n564_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n556_), .B1(new_n563_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(new_n501_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n447_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(new_n550_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n551_), .B1(new_n577_), .B2(new_n388_), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n208_), .A2(new_n255_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT74), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n208_), .A2(new_n255_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n582_), .A2(G229gat), .A3(G233gat), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n259_), .A2(new_n208_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT75), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G229gat), .A2(G233gat), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n587_), .B(KEYINPUT76), .Z(new_n588_));
  NAND3_X1  g387(.A1(new_n586_), .A2(new_n579_), .A3(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n583_), .A2(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(G113gat), .B(G141gat), .Z(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT77), .ZN(new_n592_));
  XOR2_X1   g391(.A(G169gat), .B(G197gat), .Z(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n590_), .B(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NOR4_X1   g395(.A1(new_n280_), .A2(new_n314_), .A3(new_n578_), .A4(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n597_), .A2(new_n203_), .A3(new_n447_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT105), .Z(new_n599_));
  AND2_X1   g398(.A1(new_n599_), .A2(KEYINPUT38), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n448_), .A2(new_n501_), .A3(new_n550_), .ZN(new_n601_));
  AOI22_X1  g400(.A1(new_n573_), .A2(new_n501_), .B1(new_n575_), .B2(new_n550_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n388_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n601_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n273_), .A2(new_n275_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  NOR4_X1   g406(.A1(new_n607_), .A2(new_n314_), .A3(new_n596_), .A4(new_n231_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n203_), .B1(new_n608_), .B2(new_n447_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n600_), .A2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n610_), .B1(KEYINPUT38), .B2(new_n599_), .ZN(G1324gat));
  INV_X1    g410(.A(new_n550_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n204_), .B1(new_n608_), .B2(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT39), .Z(new_n614_));
  NAND3_X1  g413(.A1(new_n597_), .A2(new_n204_), .A3(new_n612_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(G1325gat));
  AOI21_X1  g417(.A(new_n319_), .B1(new_n608_), .B2(new_n603_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT41), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n597_), .A2(new_n319_), .A3(new_n603_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(G1326gat));
  INV_X1    g421(.A(G22gat), .ZN(new_n623_));
  INV_X1    g422(.A(new_n501_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n623_), .B1(new_n608_), .B2(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT42), .Z(new_n626_));
  NAND3_X1  g425(.A1(new_n597_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(G1327gat));
  NAND2_X1  g427(.A1(new_n231_), .A2(new_n605_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT109), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n311_), .A2(new_n313_), .ZN(new_n631_));
  AND4_X1   g430(.A1(new_n604_), .A2(new_n630_), .A3(new_n595_), .A4(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(G29gat), .B1(new_n632_), .B2(new_n447_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT43), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n603_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n634_), .B(new_n278_), .C1(new_n635_), .C2(new_n551_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT107), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n604_), .A2(KEYINPUT107), .A3(new_n634_), .A4(new_n278_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n278_), .ZN(new_n640_));
  OAI21_X1  g439(.A(KEYINPUT43), .B1(new_n578_), .B2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n638_), .A2(new_n639_), .A3(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n631_), .A2(new_n595_), .A3(new_n231_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT108), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT44), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT108), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n642_), .A2(new_n648_), .A3(new_n644_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n646_), .A2(new_n647_), .A3(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n642_), .A2(KEYINPUT44), .A3(new_n644_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n447_), .A2(G29gat), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n633_), .B1(new_n653_), .B2(new_n654_), .ZN(G1328gat));
  INV_X1    g454(.A(G36gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n632_), .A2(new_n656_), .A3(new_n612_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT45), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n651_), .A2(new_n612_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n650_), .A2(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT110), .B1(new_n661_), .B2(G36gat), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT110), .ZN(new_n663_));
  AOI211_X1 g462(.A(new_n663_), .B(new_n656_), .C1(new_n650_), .C2(new_n660_), .ZN(new_n664_));
  OAI211_X1 g463(.A(KEYINPUT46), .B(new_n658_), .C1(new_n662_), .C2(new_n664_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n657_), .B(KEYINPUT45), .Z(new_n666_));
  NAND3_X1  g465(.A1(new_n661_), .A2(KEYINPUT110), .A3(G36gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(KEYINPUT44), .B1(new_n645_), .B2(KEYINPUT108), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n659_), .B1(new_n668_), .B2(new_n649_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n663_), .B1(new_n669_), .B2(new_n656_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n666_), .B1(new_n667_), .B2(new_n670_), .ZN(new_n671_));
  XOR2_X1   g470(.A(KEYINPUT111), .B(KEYINPUT46), .Z(new_n672_));
  OAI21_X1  g471(.A(new_n665_), .B1(new_n671_), .B2(new_n672_), .ZN(G1329gat));
  INV_X1    g472(.A(KEYINPUT112), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n632_), .A2(new_n603_), .ZN(new_n675_));
  INV_X1    g474(.A(G43gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n674_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n388_), .A2(new_n676_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n677_), .B1(new_n652_), .B2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT47), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n650_), .A2(new_n674_), .A3(new_n651_), .A4(new_n678_), .ZN(new_n682_));
  AND3_X1   g481(.A1(new_n680_), .A2(new_n681_), .A3(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n681_), .B1(new_n680_), .B2(new_n682_), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1330gat));
  NOR2_X1   g484(.A1(new_n501_), .A2(G50gat), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT114), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n632_), .A2(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n653_), .A2(KEYINPUT113), .A3(new_n624_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(G50gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT113), .B1(new_n653_), .B2(new_n624_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n688_), .B1(new_n690_), .B2(new_n691_), .ZN(G1331gat));
  NAND2_X1  g491(.A1(new_n314_), .A2(new_n596_), .ZN(new_n693_));
  OR3_X1    g492(.A1(new_n693_), .A2(new_n607_), .A3(new_n231_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n447_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G57gat), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  NOR4_X1   g495(.A1(new_n631_), .A2(new_n280_), .A3(new_n578_), .A4(new_n595_), .ZN(new_n697_));
  INV_X1    g496(.A(G57gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n697_), .A2(new_n698_), .A3(new_n447_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n696_), .A2(new_n699_), .ZN(G1332gat));
  OAI21_X1  g499(.A(G64gat), .B1(new_n694_), .B2(new_n550_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT48), .ZN(new_n702_));
  INV_X1    g501(.A(G64gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n697_), .A2(new_n703_), .A3(new_n612_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(G1333gat));
  OAI21_X1  g504(.A(G71gat), .B1(new_n694_), .B2(new_n388_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT49), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n388_), .A2(G71gat), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT115), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n697_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n707_), .A2(new_n710_), .ZN(G1334gat));
  OAI21_X1  g510(.A(G78gat), .B1(new_n694_), .B2(new_n501_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT50), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n697_), .A2(new_n217_), .A3(new_n624_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1335gat));
  INV_X1    g514(.A(new_n231_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n693_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n642_), .A2(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(G85gat), .B1(new_n718_), .B2(new_n695_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n630_), .A2(new_n314_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n578_), .A2(new_n595_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n447_), .A2(new_n242_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n719_), .B1(new_n722_), .B2(new_n723_), .ZN(G1336gat));
  INV_X1    g523(.A(new_n722_), .ZN(new_n725_));
  AOI21_X1  g524(.A(G92gat), .B1(new_n725_), .B2(new_n612_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n718_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n612_), .A2(G92gat), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT116), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n726_), .B1(new_n727_), .B2(new_n729_), .ZN(G1337gat));
  OAI21_X1  g529(.A(G99gat), .B1(new_n718_), .B2(new_n388_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n603_), .A2(new_n246_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(new_n722_), .B2(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g533(.A1(new_n725_), .A2(new_n624_), .A3(new_n247_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n727_), .A2(new_n624_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT52), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n736_), .A2(new_n737_), .A3(G106gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n736_), .B2(G106gat), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g540(.A(KEYINPUT57), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT55), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n294_), .A2(new_n298_), .A3(new_n743_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n296_), .A2(KEYINPUT55), .A3(new_n286_), .A4(new_n283_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n283_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(new_n299_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n305_), .B1(new_n744_), .B2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT56), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n745_), .A2(new_n747_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n294_), .A2(new_n298_), .A3(new_n743_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(KEYINPUT56), .A3(new_n305_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n751_), .A2(new_n755_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n595_), .A2(new_n308_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n588_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n586_), .A2(new_n579_), .A3(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n594_), .B1(new_n582_), .B2(new_n588_), .ZN(new_n760_));
  AOI22_X1  g559(.A1(new_n590_), .A2(new_n594_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  AOI22_X1  g560(.A1(new_n756_), .A2(new_n757_), .B1(new_n309_), .B2(new_n761_), .ZN(new_n762_));
  OAI211_X1 g561(.A(KEYINPUT118), .B(new_n742_), .C1(new_n762_), .C2(new_n605_), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT56), .B1(new_n754_), .B2(new_n305_), .ZN(new_n764_));
  AOI211_X1 g563(.A(new_n750_), .B(new_n307_), .C1(new_n752_), .C2(new_n753_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n757_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n309_), .A2(new_n761_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n605_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT118), .ZN(new_n769_));
  OAI21_X1  g568(.A(KEYINPUT57), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n308_), .A2(new_n761_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n771_), .B1(new_n751_), .B2(new_n755_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT119), .ZN(new_n773_));
  OAI21_X1  g572(.A(KEYINPUT58), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT58), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n764_), .A2(new_n765_), .ZN(new_n776_));
  OAI211_X1 g575(.A(KEYINPUT119), .B(new_n775_), .C1(new_n776_), .C2(new_n771_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n774_), .A2(new_n777_), .A3(new_n278_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n763_), .A2(new_n770_), .A3(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n231_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n279_), .B(new_n596_), .C1(new_n313_), .C2(new_n311_), .ZN(new_n781_));
  XOR2_X1   g580(.A(KEYINPUT117), .B(KEYINPUT54), .Z(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(KEYINPUT117), .A2(KEYINPUT54), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n783_), .B1(new_n781_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n780_), .A2(new_n786_), .ZN(new_n787_));
  NOR4_X1   g586(.A1(new_n624_), .A2(new_n612_), .A3(new_n695_), .A4(new_n388_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(G113gat), .B1(new_n790_), .B2(new_n595_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(KEYINPUT59), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT59), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n789_), .A2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n595_), .A2(G113gat), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT120), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n791_), .B1(new_n795_), .B2(new_n797_), .ZN(G1340gat));
  INV_X1    g597(.A(G120gat), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n799_), .B1(new_n631_), .B2(KEYINPUT60), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n790_), .B(new_n800_), .C1(KEYINPUT60), .C2(new_n799_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n631_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(new_n799_), .ZN(G1341gat));
  INV_X1    g602(.A(G127gat), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n804_), .B1(new_n789_), .B2(new_n231_), .ZN(new_n805_));
  OR2_X1    g604(.A1(new_n805_), .A2(KEYINPUT121), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(KEYINPUT121), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n231_), .A2(new_n804_), .ZN(new_n808_));
  AOI22_X1  g607(.A1(new_n806_), .A2(new_n807_), .B1(new_n795_), .B2(new_n808_), .ZN(G1342gat));
  INV_X1    g608(.A(G134gat), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n790_), .A2(new_n810_), .A3(new_n605_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n640_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n812_), .B2(new_n810_), .ZN(G1343gat));
  NOR4_X1   g612(.A1(new_n612_), .A2(new_n501_), .A3(new_n695_), .A4(new_n603_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(KEYINPUT122), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n787_), .A2(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n816_), .A2(new_n596_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(new_n397_), .ZN(G1344gat));
  NOR2_X1   g617(.A1(new_n816_), .A2(new_n631_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(new_n398_), .ZN(G1345gat));
  INV_X1    g619(.A(KEYINPUT123), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n821_), .B1(new_n816_), .B2(new_n231_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n787_), .A2(KEYINPUT123), .A3(new_n716_), .A4(new_n815_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(KEYINPUT61), .B(G155gat), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n822_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n824_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(G1346gat));
  OAI21_X1  g626(.A(G162gat), .B1(new_n816_), .B2(new_n640_), .ZN(new_n828_));
  OR2_X1    g627(.A1(new_n606_), .A2(G162gat), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n816_), .B2(new_n829_), .ZN(G1347gat));
  INV_X1    g629(.A(KEYINPUT62), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n785_), .B1(new_n779_), .B2(new_n231_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n612_), .A2(new_n448_), .ZN(new_n833_));
  NOR4_X1   g632(.A1(new_n832_), .A2(new_n624_), .A3(new_n596_), .A4(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(G169gat), .B1(new_n834_), .B2(KEYINPUT124), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n832_), .A2(new_n624_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n833_), .ZN(new_n837_));
  AND4_X1   g636(.A1(KEYINPUT124), .A2(new_n836_), .A3(new_n595_), .A4(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n831_), .B1(new_n835_), .B2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n836_), .A2(new_n595_), .A3(new_n837_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT124), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n834_), .A2(KEYINPUT124), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n842_), .A2(KEYINPUT62), .A3(new_n843_), .A4(G169gat), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n834_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n839_), .A2(new_n844_), .A3(new_n845_), .ZN(G1348gat));
  INV_X1    g645(.A(new_n836_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT125), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT125), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n836_), .A2(new_n849_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n848_), .A2(new_n850_), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n314_), .A2(G176gat), .A3(new_n837_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n847_), .A2(new_n833_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n314_), .ZN(new_n854_));
  AOI22_X1  g653(.A1(new_n851_), .A2(new_n852_), .B1(new_n854_), .B2(new_n362_), .ZN(G1349gat));
  NAND4_X1  g654(.A1(new_n848_), .A2(new_n850_), .A3(new_n716_), .A4(new_n837_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n716_), .A2(new_n513_), .ZN(new_n857_));
  AOI22_X1  g656(.A1(new_n856_), .A2(new_n337_), .B1(new_n853_), .B2(new_n857_), .ZN(G1350gat));
  INV_X1    g657(.A(new_n514_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n853_), .A2(new_n859_), .A3(new_n605_), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n847_), .A2(new_n640_), .A3(new_n833_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n861_), .B2(new_n332_), .ZN(G1351gat));
  AND3_X1   g661(.A1(new_n612_), .A2(new_n575_), .A3(new_n388_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n787_), .A2(new_n863_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n864_), .A2(new_n596_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(new_n451_), .ZN(G1352gat));
  INV_X1    g665(.A(new_n864_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n314_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT126), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(G204gat), .ZN(new_n870_));
  XNOR2_X1  g669(.A(KEYINPUT126), .B(G204gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n868_), .B2(new_n871_), .ZN(G1353gat));
  NOR2_X1   g671(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n873_));
  AND2_X1   g672(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n874_));
  NOR4_X1   g673(.A1(new_n864_), .A2(new_n231_), .A3(new_n873_), .A4(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n867_), .A2(new_n716_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n876_), .B2(new_n873_), .ZN(G1354gat));
  NOR3_X1   g676(.A1(new_n864_), .A2(new_n458_), .A3(new_n640_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n864_), .A2(new_n606_), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n879_), .A2(KEYINPUT127), .ZN(new_n880_));
  AOI21_X1  g679(.A(G218gat), .B1(new_n879_), .B2(KEYINPUT127), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n878_), .B1(new_n880_), .B2(new_n881_), .ZN(G1355gat));
endmodule


