//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 0 0 1 0 0 1 0 1 0 1 1 1 1 0 0 1 0 1 0 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n631_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n863_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_;
  NOR2_X1   g000(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G169gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G183gat), .A3(G190gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  AOI21_X1  g005(.A(new_n204_), .B1(G183gat), .B2(G190gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n203_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G169gat), .ZN(new_n211_));
  INV_X1    g010(.A(G176gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT24), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  MUX2_X1   g013(.A(new_n213_), .B(KEYINPUT24), .S(new_n214_), .Z(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT25), .B(G183gat), .ZN(new_n216_));
  INV_X1    g015(.A(G190gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(KEYINPUT81), .A3(KEYINPUT26), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT81), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT26), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n219_), .B1(new_n220_), .B2(G190gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n216_), .A2(new_n218_), .A3(new_n221_), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n220_), .A2(KEYINPUT82), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n220_), .A2(KEYINPUT82), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n217_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n215_), .B1(new_n222_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT83), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n205_), .B(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n228_), .A2(new_n207_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n210_), .B1(new_n226_), .B2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT30), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G227gat), .A2(G233gat), .ZN(new_n232_));
  INV_X1    g031(.A(G15gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(G71gat), .ZN(new_n235_));
  INV_X1    g034(.A(G99gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n231_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT86), .B(KEYINPUT31), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT87), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n238_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G127gat), .B(G134gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G113gat), .B(G120gat), .ZN(new_n244_));
  AOI21_X1  g043(.A(KEYINPUT85), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  XOR2_X1   g044(.A(G127gat), .B(G134gat), .Z(new_n246_));
  XOR2_X1   g045(.A(G113gat), .B(G120gat), .Z(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n245_), .B(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(KEYINPUT84), .B(G43gat), .Z(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n242_), .B(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G22gat), .B(G50gat), .ZN(new_n253_));
  XOR2_X1   g052(.A(KEYINPUT89), .B(G197gat), .Z(new_n254_));
  NOR2_X1   g053(.A1(new_n254_), .A2(G204gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT90), .B(G204gat), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n256_), .A2(G197gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT21), .B1(new_n255_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n254_), .A2(G204gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT21), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n256_), .A2(G197gat), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n259_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G211gat), .B(G218gat), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n258_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n259_), .A2(new_n261_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n263_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(KEYINPUT21), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G141gat), .A2(G148gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT2), .ZN(new_n269_));
  NOR2_X1   g068(.A1(G141gat), .A2(G148gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT88), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT3), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n270_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n271_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT3), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n269_), .A2(new_n273_), .A3(new_n275_), .ZN(new_n276_));
  AND2_X1   g075(.A1(G155gat), .A2(G162gat), .ZN(new_n277_));
  NOR2_X1   g076(.A1(G155gat), .A2(G162gat), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n276_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT1), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n277_), .A2(KEYINPUT1), .ZN(new_n283_));
  INV_X1    g082(.A(new_n270_), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n282_), .A2(new_n283_), .A3(new_n268_), .A4(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n280_), .A2(new_n285_), .ZN(new_n286_));
  AOI22_X1  g085(.A1(new_n264_), .A2(new_n267_), .B1(new_n286_), .B2(KEYINPUT29), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G228gat), .A2(G233gat), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT91), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  NOR3_X1   g090(.A1(new_n287_), .A2(G78gat), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(G78gat), .B1(new_n287_), .B2(new_n291_), .ZN(new_n294_));
  AOI21_X1  g093(.A(G106gat), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(G78gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n264_), .A2(new_n267_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n286_), .A2(KEYINPUT29), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n296_), .B1(new_n299_), .B2(new_n290_), .ZN(new_n300_));
  INV_X1    g099(.A(G106gat), .ZN(new_n301_));
  NOR3_X1   g100(.A1(new_n300_), .A2(new_n292_), .A3(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n253_), .B1(new_n295_), .B2(new_n302_), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n286_), .A2(KEYINPUT29), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT28), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n288_), .A2(new_n289_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n305_), .B(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n293_), .A2(G106gat), .A3(new_n294_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n301_), .B1(new_n300_), .B2(new_n292_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n253_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  AND3_X1   g111(.A1(new_n303_), .A2(new_n308_), .A3(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n308_), .B1(new_n303_), .B2(new_n312_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(G8gat), .B(G36gat), .Z(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT93), .ZN(new_n317_));
  XOR2_X1   g116(.A(G64gat), .B(G92gat), .Z(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT94), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n317_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G226gat), .A2(G233gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT19), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n203_), .B1(new_n229_), .B2(new_n209_), .ZN(new_n325_));
  XOR2_X1   g124(.A(KEYINPUT26), .B(G190gat), .Z(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n208_), .B1(new_n216_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(new_n215_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n325_), .A2(new_n264_), .A3(new_n267_), .A4(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT20), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT101), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n297_), .A2(new_n230_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n331_), .A2(new_n332_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n324_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT20), .B1(new_n297_), .B2(new_n230_), .ZN(new_n338_));
  AOI22_X1  g137(.A1(new_n325_), .A2(new_n329_), .B1(new_n264_), .B2(new_n267_), .ZN(new_n339_));
  OR3_X1    g138(.A1(new_n338_), .A2(new_n339_), .A3(new_n324_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n322_), .B1(new_n337_), .B2(new_n340_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n324_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n324_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n334_), .A2(KEYINPUT20), .A3(new_n330_), .A4(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n342_), .A2(new_n322_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT103), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND4_X1  g146(.A1(new_n342_), .A2(new_n322_), .A3(KEYINPUT103), .A4(new_n344_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT27), .B1(new_n341_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT95), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n345_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n342_), .A2(new_n344_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n322_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT27), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n342_), .A2(new_n322_), .A3(KEYINPUT95), .A4(new_n344_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n352_), .A2(new_n355_), .A3(new_n356_), .A4(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n350_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G225gat), .A2(G233gat), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT4), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n249_), .A2(new_n286_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n246_), .B(new_n244_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n363_), .B(KEYINPUT96), .C1(new_n286_), .C2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT96), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n249_), .A2(new_n366_), .A3(new_n286_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n362_), .B1(new_n365_), .B2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n363_), .A2(KEYINPUT4), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n361_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n365_), .A2(new_n360_), .A3(new_n367_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G1gat), .B(G29gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(G85gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT0), .B(G57gat), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n374_), .B(new_n375_), .Z(new_n376_));
  NAND2_X1  g175(.A1(new_n372_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n376_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n370_), .A2(new_n378_), .A3(new_n371_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n377_), .A2(KEYINPUT102), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT102), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n372_), .A2(new_n381_), .A3(new_n376_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n315_), .A2(new_n359_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT104), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT104), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n315_), .A2(new_n359_), .A3(new_n386_), .A4(new_n383_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n352_), .A2(new_n357_), .A3(new_n355_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n365_), .A2(new_n367_), .ZN(new_n390_));
  OR2_X1    g189(.A1(new_n390_), .A2(KEYINPUT99), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n360_), .B1(new_n390_), .B2(KEYINPUT99), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n376_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n369_), .B1(new_n390_), .B2(KEYINPUT4), .ZN(new_n394_));
  AOI21_X1  g193(.A(KEYINPUT100), .B1(new_n394_), .B2(new_n360_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT100), .ZN(new_n396_));
  NOR4_X1   g195(.A1(new_n368_), .A2(new_n396_), .A3(new_n361_), .A4(new_n369_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n393_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n389_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT97), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n378_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n400_), .B1(new_n401_), .B2(KEYINPUT33), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n399_), .A2(new_n402_), .ZN(new_n403_));
  OR3_X1    g202(.A1(new_n401_), .A2(KEYINPUT98), .A3(KEYINPUT33), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT98), .B1(new_n401_), .B2(KEYINPUT33), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n401_), .A2(new_n400_), .A3(KEYINPUT33), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n403_), .A2(new_n406_), .A3(new_n408_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n322_), .A2(KEYINPUT32), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n410_), .A2(new_n353_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n337_), .A2(new_n340_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n411_), .B1(new_n412_), .B2(new_n410_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n380_), .A2(new_n382_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n315_), .B1(new_n409_), .B2(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n252_), .B1(new_n388_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n359_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n383_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n252_), .A2(new_n315_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n417_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT70), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G57gat), .B(G64gat), .ZN(new_n425_));
  OR2_X1    g224(.A1(new_n425_), .A2(KEYINPUT11), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(KEYINPUT11), .ZN(new_n427_));
  XOR2_X1   g226(.A(G71gat), .B(G78gat), .Z(new_n428_));
  NAND3_X1  g227(.A1(new_n426_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n427_), .A2(new_n428_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(KEYINPUT10), .B(G99gat), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n432_), .A2(G106gat), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n433_), .A2(KEYINPUT64), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(KEYINPUT64), .ZN(new_n435_));
  INV_X1    g234(.A(G85gat), .ZN(new_n436_));
  INV_X1    g235(.A(G92gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G85gat), .A2(G92gat), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(KEYINPUT9), .A3(new_n439_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n439_), .A2(KEYINPUT9), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT6), .B1(new_n236_), .B2(new_n301_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT6), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n443_), .A2(G99gat), .A3(G106gat), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n441_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n434_), .A2(new_n435_), .A3(new_n440_), .A4(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT8), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT65), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT7), .ZN(new_n449_));
  OAI211_X1 g248(.A(new_n448_), .B(new_n449_), .C1(G99gat), .C2(G106gat), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n236_), .B(new_n301_), .C1(KEYINPUT65), .C2(KEYINPUT7), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT67), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n450_), .A2(new_n451_), .A3(KEYINPUT67), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n442_), .A2(new_n444_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n454_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n438_), .A2(new_n439_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT66), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n438_), .A2(KEYINPUT66), .A3(new_n439_), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n447_), .B1(new_n457_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n460_), .A2(new_n461_), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n450_), .A2(new_n451_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n465_));
  NOR3_X1   g264(.A1(new_n464_), .A2(new_n465_), .A3(KEYINPUT8), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n431_), .B(new_n446_), .C1(new_n463_), .C2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G230gat), .A2(G233gat), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n467_), .A2(KEYINPUT69), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(KEYINPUT69), .B1(new_n467_), .B2(new_n468_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n431_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT68), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n473_), .A2(KEYINPUT12), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n457_), .A2(new_n462_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n466_), .B1(new_n476_), .B2(KEYINPUT8), .ZN(new_n477_));
  INV_X1    g276(.A(new_n446_), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n472_), .B(new_n475_), .C1(new_n477_), .C2(new_n478_), .ZN(new_n479_));
  AOI22_X1  g278(.A1(new_n452_), .A2(new_n453_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n464_), .B1(new_n480_), .B2(new_n455_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n462_), .A2(new_n447_), .ZN(new_n482_));
  OAI22_X1  g281(.A1(new_n481_), .A2(new_n447_), .B1(new_n482_), .B2(new_n465_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n431_), .B1(new_n483_), .B2(new_n446_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT68), .B(KEYINPUT12), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n479_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n424_), .B1(new_n471_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n468_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n467_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n488_), .B1(new_n484_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n467_), .A2(new_n468_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT69), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n467_), .A2(KEYINPUT69), .A3(new_n468_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n446_), .B1(new_n463_), .B2(new_n466_), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n496_), .A2(new_n472_), .A3(new_n475_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n485_), .B1(new_n496_), .B2(new_n472_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n495_), .A2(new_n499_), .A3(KEYINPUT70), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n487_), .A2(new_n490_), .A3(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(KEYINPUT71), .B(KEYINPUT5), .Z(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT72), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G120gat), .B(G148gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G176gat), .B(G204gat), .ZN(new_n506_));
  XOR2_X1   g305(.A(new_n505_), .B(new_n506_), .Z(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n501_), .A2(new_n508_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n487_), .A2(new_n500_), .A3(new_n490_), .A4(new_n507_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT13), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n509_), .A2(KEYINPUT13), .A3(new_n510_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(G29gat), .B(G36gat), .Z(new_n516_));
  XOR2_X1   g315(.A(G43gat), .B(G50gat), .Z(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G29gat), .B(G36gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G43gat), .B(G50gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n518_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT80), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G15gat), .B(G22gat), .ZN(new_n524_));
  INV_X1    g323(.A(G1gat), .ZN(new_n525_));
  INV_X1    g324(.A(G8gat), .ZN(new_n526_));
  OAI21_X1  g325(.A(KEYINPUT14), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT77), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n524_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n527_), .A2(new_n528_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G1gat), .B(G8gat), .ZN(new_n531_));
  OR3_X1    g330(.A1(new_n529_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n531_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n523_), .B(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G229gat), .A2(G233gat), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n535_), .A2(new_n537_), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n523_), .A2(new_n534_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n522_), .B(KEYINPUT15), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n534_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n539_), .A2(new_n536_), .A3(new_n541_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n538_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G113gat), .B(G141gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G169gat), .B(G197gat), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n544_), .B(new_n545_), .Z(new_n546_));
  XNOR2_X1  g345(.A(new_n543_), .B(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n515_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n423_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT79), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G231gat), .A2(G233gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n534_), .B(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(new_n472_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n554_), .A2(KEYINPUT78), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(G127gat), .B(G155gat), .Z(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT16), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G183gat), .B(G211gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n560_), .A2(KEYINPUT17), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n560_), .B1(new_n554_), .B2(KEYINPUT17), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n556_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n556_), .B1(new_n562_), .B2(new_n561_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n551_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n562_), .A2(new_n561_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(new_n555_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n568_), .A2(KEYINPUT79), .A3(new_n563_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n566_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n496_), .A2(new_n540_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n483_), .A2(new_n522_), .A3(new_n446_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(G232gat), .A2(G233gat), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n573_), .B(KEYINPUT34), .Z(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT73), .B(KEYINPUT35), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n574_), .A2(new_n575_), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n571_), .A2(new_n572_), .A3(new_n577_), .A4(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT74), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n571_), .A2(new_n572_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n580_), .B1(new_n581_), .B2(new_n576_), .ZN(new_n582_));
  AOI211_X1 g381(.A(KEYINPUT74), .B(new_n577_), .C1(new_n571_), .C2(new_n572_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n579_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G190gat), .B(G218gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT75), .ZN(new_n586_));
  XOR2_X1   g385(.A(G134gat), .B(G162gat), .Z(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n588_), .A2(KEYINPUT36), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(KEYINPUT36), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n584_), .A2(new_n590_), .A3(new_n591_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n589_), .B(new_n579_), .C1(new_n582_), .C2(new_n583_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT76), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n593_), .A2(new_n594_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n592_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT37), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  OAI211_X1 g398(.A(KEYINPUT37), .B(new_n592_), .C1(new_n595_), .C2(new_n596_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n570_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n550_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n602_), .A2(new_n525_), .A3(new_n419_), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n603_), .B(KEYINPUT38), .Z(new_n604_));
  INV_X1    g403(.A(new_n597_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n564_), .A2(new_n565_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n550_), .A2(new_n605_), .A3(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n525_), .B1(new_n608_), .B2(new_n419_), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n604_), .A2(new_n609_), .ZN(G1324gat));
  NAND3_X1  g409(.A1(new_n602_), .A2(new_n526_), .A3(new_n418_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT39), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n608_), .A2(new_n418_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n612_), .B1(new_n613_), .B2(G8gat), .ZN(new_n614_));
  AOI211_X1 g413(.A(KEYINPUT39), .B(new_n526_), .C1(new_n608_), .C2(new_n418_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n611_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT40), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  OAI211_X1 g417(.A(KEYINPUT40), .B(new_n611_), .C1(new_n614_), .C2(new_n615_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(G1325gat));
  INV_X1    g419(.A(new_n252_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n233_), .B1(new_n608_), .B2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT41), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n602_), .A2(new_n233_), .A3(new_n621_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(G1326gat));
  INV_X1    g424(.A(G22gat), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n602_), .A2(new_n626_), .A3(new_n315_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n608_), .A2(new_n315_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n628_), .A2(G22gat), .A3(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n628_), .B2(G22gat), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n627_), .B1(new_n630_), .B2(new_n631_), .ZN(G1327gat));
  INV_X1    g431(.A(new_n422_), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n399_), .A2(new_n407_), .A3(new_n402_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n414_), .B1(new_n634_), .B2(new_n406_), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n385_), .B(new_n387_), .C1(new_n635_), .C2(new_n315_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n633_), .B1(new_n636_), .B2(new_n252_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n549_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n570_), .A2(new_n597_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  OR3_X1    g440(.A1(new_n641_), .A2(G29gat), .A3(new_n383_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n599_), .A2(new_n600_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n423_), .A2(KEYINPUT107), .A3(KEYINPUT43), .A4(new_n643_), .ZN(new_n644_));
  OR2_X1    g443(.A1(KEYINPUT107), .A2(KEYINPUT43), .ZN(new_n645_));
  NAND2_X1  g444(.A1(KEYINPUT107), .A2(KEYINPUT43), .ZN(new_n646_));
  INV_X1    g445(.A(new_n643_), .ZN(new_n647_));
  OAI211_X1 g446(.A(new_n645_), .B(new_n646_), .C1(new_n637_), .C2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n570_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n549_), .A2(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT106), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n644_), .A2(new_n648_), .A3(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT44), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n644_), .A2(new_n648_), .A3(KEYINPUT44), .A4(new_n651_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n419_), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT108), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n656_), .A2(new_n657_), .A3(G29gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n656_), .B2(G29gat), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n642_), .B1(new_n658_), .B2(new_n659_), .ZN(G1328gat));
  NAND3_X1  g459(.A1(new_n654_), .A2(new_n418_), .A3(new_n655_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(G36gat), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n359_), .A2(G36gat), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n423_), .A2(new_n549_), .A3(new_n640_), .A4(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT109), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT109), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n639_), .A2(new_n666_), .A3(new_n640_), .A4(new_n663_), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n665_), .A2(new_n667_), .A3(KEYINPUT45), .ZN(new_n668_));
  AOI21_X1  g467(.A(KEYINPUT45), .B1(new_n665_), .B2(new_n667_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n662_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT46), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n662_), .A2(KEYINPUT46), .A3(new_n670_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1329gat));
  NAND4_X1  g474(.A1(new_n654_), .A2(G43gat), .A3(new_n621_), .A4(new_n655_), .ZN(new_n676_));
  INV_X1    g475(.A(G43gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n677_), .B1(new_n641_), .B2(new_n252_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g479(.A1(new_n654_), .A2(G50gat), .A3(new_n315_), .A4(new_n655_), .ZN(new_n681_));
  INV_X1    g480(.A(G50gat), .ZN(new_n682_));
  INV_X1    g481(.A(new_n315_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n682_), .B1(new_n641_), .B2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n681_), .A2(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT110), .ZN(G1331gat));
  INV_X1    g485(.A(new_n515_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n601_), .A2(new_n687_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT111), .Z(new_n689_));
  NOR3_X1   g488(.A1(new_n689_), .A2(new_n547_), .A3(new_n637_), .ZN(new_n690_));
  INV_X1    g489(.A(G57gat), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n690_), .A2(new_n691_), .A3(new_n419_), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n637_), .A2(new_n547_), .A3(new_n687_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n693_), .A2(new_n597_), .A3(new_n570_), .ZN(new_n694_));
  OAI21_X1  g493(.A(G57gat), .B1(new_n694_), .B2(new_n383_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n692_), .A2(new_n695_), .ZN(G1332gat));
  OAI21_X1  g495(.A(G64gat), .B1(new_n694_), .B2(new_n359_), .ZN(new_n697_));
  XOR2_X1   g496(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(G64gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n690_), .A2(new_n700_), .A3(new_n418_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(G1333gat));
  OAI21_X1  g501(.A(G71gat), .B1(new_n694_), .B2(new_n252_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT49), .ZN(new_n704_));
  INV_X1    g503(.A(G71gat), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n690_), .A2(new_n705_), .A3(new_n621_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(G1334gat));
  NAND2_X1  g506(.A1(new_n315_), .A2(new_n296_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT113), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n690_), .A2(new_n709_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n693_), .A2(new_n315_), .A3(new_n597_), .A4(new_n570_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT50), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n711_), .A2(new_n712_), .A3(G78gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n712_), .B1(new_n711_), .B2(G78gat), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n710_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT114), .ZN(G1335gat));
  NAND3_X1  g515(.A1(new_n649_), .A2(new_n548_), .A3(new_n515_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n644_), .A2(new_n648_), .A3(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT115), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n644_), .A2(new_n648_), .A3(KEYINPUT115), .A4(new_n718_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n383_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n693_), .A2(new_n640_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n419_), .A2(new_n436_), .ZN(new_n725_));
  OAI22_X1  g524(.A1(new_n723_), .A2(new_n436_), .B1(new_n724_), .B2(new_n725_), .ZN(G1336gat));
  OAI21_X1  g525(.A(new_n437_), .B1(new_n724_), .B2(new_n359_), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n727_), .B(KEYINPUT116), .Z(new_n728_));
  NAND2_X1  g527(.A1(new_n721_), .A2(new_n722_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n359_), .A2(new_n437_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n728_), .B1(new_n729_), .B2(new_n730_), .ZN(G1337gat));
  OR3_X1    g530(.A1(new_n724_), .A2(new_n432_), .A3(new_n252_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n252_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(new_n236_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(KEYINPUT51), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT51), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n736_), .B(new_n732_), .C1(new_n733_), .C2(new_n236_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1338gat));
  NAND4_X1  g537(.A1(new_n693_), .A2(new_n301_), .A3(new_n315_), .A4(new_n640_), .ZN(new_n739_));
  NAND4_X1  g538(.A1(new_n644_), .A2(new_n648_), .A3(new_n315_), .A4(new_n718_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT52), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n740_), .A2(new_n741_), .A3(G106gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n740_), .B2(G106gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n739_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT53), .ZN(G1339gat));
  XNOR2_X1  g544(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n515_), .A2(new_n547_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n747_), .B1(new_n749_), .B2(new_n601_), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n748_), .A2(new_n647_), .A3(new_n570_), .A4(new_n746_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n538_), .A2(new_n542_), .A3(new_n546_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT118), .ZN(new_n754_));
  AND3_X1   g553(.A1(new_n539_), .A2(new_n754_), .A3(new_n541_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n539_), .B2(new_n541_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n755_), .A2(new_n756_), .A3(new_n536_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n535_), .A2(new_n536_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n546_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n753_), .B1(new_n757_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n511_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT119), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT119), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n511_), .A2(new_n765_), .A3(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n547_), .A2(new_n510_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n487_), .A2(new_n769_), .A3(new_n500_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n486_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n479_), .B(new_n467_), .C1(new_n484_), .C2(new_n485_), .ZN(new_n772_));
  AOI22_X1  g571(.A1(new_n771_), .A2(KEYINPUT55), .B1(new_n488_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n770_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n508_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT56), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n774_), .A2(KEYINPUT56), .A3(new_n508_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n768_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n597_), .B1(new_n767_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT57), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n777_), .A2(new_n778_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n762_), .A2(new_n510_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT58), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT56), .B1(new_n774_), .B2(new_n508_), .ZN(new_n788_));
  AOI211_X1 g587(.A(new_n776_), .B(new_n507_), .C1(new_n770_), .C2(new_n773_), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n784_), .B(KEYINPUT58), .C1(new_n788_), .C2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n787_), .A2(new_n643_), .A3(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n768_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n792_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n793_), .A2(new_n764_), .A3(new_n766_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(KEYINPUT57), .A3(new_n597_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n782_), .A2(new_n791_), .A3(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n752_), .B1(new_n796_), .B2(new_n607_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n421_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n418_), .A2(new_n383_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n797_), .A2(new_n798_), .A3(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT59), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n752_), .B1(new_n796_), .B2(new_n649_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n800_), .A2(new_n798_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n802_), .ZN(new_n805_));
  OAI22_X1  g604(.A1(new_n801_), .A2(new_n802_), .B1(new_n803_), .B2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(G113gat), .B1(new_n806_), .B2(new_n548_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT120), .ZN(new_n808_));
  INV_X1    g607(.A(new_n752_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n765_), .B1(new_n511_), .B2(new_n762_), .ZN(new_n810_));
  AOI211_X1 g609(.A(KEYINPUT119), .B(new_n761_), .C1(new_n509_), .C2(new_n510_), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  AOI211_X1 g611(.A(new_n781_), .B(new_n605_), .C1(new_n812_), .C2(new_n793_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT57), .B1(new_n794_), .B2(new_n597_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT58), .B1(new_n783_), .B2(new_n784_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n790_), .A2(new_n643_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n813_), .A2(new_n814_), .A3(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n809_), .B1(new_n818_), .B2(new_n606_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n804_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n820_), .A2(G113gat), .A3(new_n548_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n807_), .A2(new_n808_), .A3(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(G113gat), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n803_), .A2(new_n805_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n825_), .B1(new_n820_), .B2(KEYINPUT59), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n824_), .B1(new_n826_), .B2(new_n547_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT120), .B1(new_n827_), .B2(new_n821_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n823_), .A2(new_n828_), .ZN(G1340gat));
  XOR2_X1   g628(.A(KEYINPUT121), .B(G120gat), .Z(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(new_n687_), .B2(KEYINPUT60), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n801_), .B(new_n831_), .C1(KEYINPUT60), .C2(new_n830_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n806_), .A2(new_n687_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n832_), .B1(new_n833_), .B2(new_n830_), .ZN(G1341gat));
  INV_X1    g633(.A(G127gat), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n806_), .A2(new_n835_), .A3(new_n607_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n820_), .B2(new_n649_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT122), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n837_), .A2(new_n838_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n836_), .A2(new_n839_), .A3(new_n840_), .ZN(G1342gat));
  OAI21_X1  g640(.A(G134gat), .B1(new_n806_), .B2(new_n647_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT123), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n820_), .A2(G134gat), .A3(new_n597_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n842_), .A2(new_n843_), .A3(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(G134gat), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n847_), .B1(new_n826_), .B2(new_n643_), .ZN(new_n848_));
  OAI21_X1  g647(.A(KEYINPUT123), .B1(new_n848_), .B2(new_n844_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n846_), .A2(new_n849_), .ZN(G1343gat));
  NOR2_X1   g649(.A1(new_n621_), .A2(new_n683_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n799_), .ZN(new_n852_));
  OAI21_X1  g651(.A(KEYINPUT124), .B1(new_n797_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT124), .ZN(new_n854_));
  INV_X1    g653(.A(new_n852_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n813_), .A2(new_n814_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n606_), .B1(new_n856_), .B2(new_n791_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n854_), .B(new_n855_), .C1(new_n857_), .C2(new_n752_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n853_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n547_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n860_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g660(.A1(new_n859_), .A2(new_n515_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT125), .B(G148gat), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(G1345gat));
  XNOR2_X1  g663(.A(KEYINPUT126), .B(KEYINPUT127), .ZN(new_n865_));
  INV_X1    g664(.A(new_n865_), .ZN(new_n866_));
  XOR2_X1   g665(.A(KEYINPUT61), .B(G155gat), .Z(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n868_), .B1(new_n859_), .B2(new_n570_), .ZN(new_n869_));
  AOI211_X1 g668(.A(new_n649_), .B(new_n867_), .C1(new_n853_), .C2(new_n858_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n866_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n854_), .B1(new_n819_), .B2(new_n855_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n797_), .A2(KEYINPUT124), .A3(new_n852_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n570_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n867_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n859_), .A2(new_n570_), .A3(new_n868_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n875_), .A2(new_n865_), .A3(new_n876_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n871_), .A2(new_n877_), .ZN(G1346gat));
  INV_X1    g677(.A(new_n859_), .ZN(new_n879_));
  OR3_X1    g678(.A1(new_n879_), .A2(G162gat), .A3(new_n597_), .ZN(new_n880_));
  OAI21_X1  g679(.A(G162gat), .B1(new_n879_), .B2(new_n647_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1347gat));
  INV_X1    g681(.A(KEYINPUT62), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n421_), .A2(new_n383_), .A3(new_n418_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n803_), .A2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n886_), .A2(new_n548_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT22), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n883_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(G169gat), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n211_), .B1(new_n887_), .B2(new_n883_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n889_), .B2(new_n891_), .ZN(G1348gat));
  OR2_X1    g691(.A1(new_n797_), .A2(new_n884_), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n893_), .A2(new_n212_), .A3(new_n687_), .ZN(new_n894_));
  AOI21_X1  g693(.A(G176gat), .B1(new_n885_), .B2(new_n515_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1349gat));
  OR2_X1    g695(.A1(new_n893_), .A2(new_n649_), .ZN(new_n897_));
  INV_X1    g696(.A(G183gat), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n607_), .A2(new_n216_), .ZN(new_n899_));
  AOI22_X1  g698(.A1(new_n897_), .A2(new_n898_), .B1(new_n885_), .B2(new_n899_), .ZN(G1350gat));
  OAI21_X1  g699(.A(G190gat), .B1(new_n886_), .B2(new_n647_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n885_), .A2(new_n327_), .A3(new_n605_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1351gat));
  NAND3_X1  g702(.A1(new_n851_), .A2(new_n383_), .A3(new_n418_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n797_), .A2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n547_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g706(.A1(new_n905_), .A2(new_n515_), .ZN(new_n908_));
  MUX2_X1   g707(.A(new_n256_), .B(G204gat), .S(new_n908_), .Z(G1353gat));
  NAND2_X1  g708(.A1(new_n905_), .A2(new_n606_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n911_));
  AND2_X1   g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n910_), .A2(new_n911_), .A3(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n913_), .B1(new_n910_), .B2(new_n911_), .ZN(G1354gat));
  INV_X1    g713(.A(G218gat), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n905_), .A2(new_n915_), .A3(new_n605_), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n797_), .A2(new_n647_), .A3(new_n904_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(new_n915_), .ZN(G1355gat));
endmodule


